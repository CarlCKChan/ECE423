��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�+����Rq�����������+�nS�U�F7&���S����"�M ��U���@�˴�5��.� -;P�~�oa|
)k���BЖ�@�o�v�4ߘ<��4�l��D�4Ak���-.b���mC*��D�i�M%��%�k�~&ʳ��0!����nY�qe��3��ck����o��z"��,f�ը��%$���|�;+#�0f�UhOǃ��2刑�Lc�����|��|����Q��Ol�pf��\�4Y�
A�Y�a@��qnNAz�pד��ݮiF�?��'~&{�X�v����H�	���Gʲ���dӤ�>v�� ���K�B�x��X�[#s��W�V��.��f$�n���:Qn��24"M��<48�}[�� �(�5��t�L�6����ئe3Xa�|=�X$nD�H"ď�Vl��⼞=��5��n�Q���6;#٬"I�L���P����/P=�}�㟂���C���?�ZI�r�	5��]%���ē�2FTC�Sh��Ds]鉬�@�0:�?"ܮAۙ�>���?��i+c��$�vf�:��P����LX�Z��+�'��Y�}�G��)��q��ʋ�X�]���ۅЅ�aڴG��i����(ް?	�P9���y�
�����E==6�iS��=م�gU����!��8�د�§���g��d���B�Rx%��E}��8�!-�U��@=�R ��s�/�ǥ�;,'�f��|�<�\W�21u�a���{-��������k�����@b��G�9SK{[O��Y��7�vb���yS�����	�63ǲ�Sr�,B�/�t�(��� bc";W���"-�����?�1\�ؤ'

`�x��4Q.�H����E�l���5��S���kd1��{+Hڔ�խ8�|$�������؄+����)���gn��+砯y���>3T��Xw5ӗ<,�C���   ̰�78ys
7�s�m�MO���_���t�3���d���*�۱�)!܃�9��-�J���.��qkT�*)�
0�Fx����t�g#@p��s���(��ܐ�q��U)ײ�Zƚś�!����qp� }�̚ޒ��	�v4����l�a�+|Eۺ�m�%��~�K~�u/+Em����	����������O�����閐��q�p�4��H@n�� N}���dv��m?�:�>!���GK���7r�H�0O��ߙ�	�N,���;�XG�Hw���2�d�lD��
�ϻY>�R���`������R�i�[~�~�<0�|�8t!��l*�,p49Ọ�2Vj������N~EG8��!S�K���͙�}IjV���l���1��Cz&3���\'(��]AG�0Z}?���=�bLϛ�A��3%�$�[G�j�fuA'�ٰ0�q�,����\�I���w�%�7pc�/ ���'t|�M�-�X3U �������fܨ�ZI	�:�:͙(:��}$@Fۢ��q|Le)Q�>C���ӆ[�1���E=A�	��j��WQ��;9�L�S�V����X�,�`������DY,�m�?��!!vC�yu��Ȣ%������S!G=3��i �t�2h,q�&�"���'+t����L�G��_�/QNvsN�UK�@+���[#��yfK�+�2)��/� =�v>3�(>r�'�(Abz!8{��>�G��Y��ϕ���5�
aiY��%ZӰ^#�KJ�7�_����r�90�"Hf�T�F ĳ#4�˟��?��ف�2@�F���Ƃ����M�]>�6Sy3!����=,C Zʺ�}p���݂�<�\��	kI�O�>�~�?=�jXF[XX�� �\)�h�\�v�GE�hOZ��y��6*I�(�ϱJgٕ6� {�� �l``;ʟ�`F�%{Tѱ� ?I�K�^�?�G��V�}t"��V��oń\���V׿� ��{9q_�� �\���F���LJ�����tn
ǏK�񍱖��}c88+¾R�Yd�]���R�2���W�+�Pw`ބ�������%[E�J"+�����q��0� �Ȏ��vML�צ��g֒��3��|��`��&9} ������\t�y9��w�*���k�[��x����f�!��캩�G;�ǻ
VA'�XS�B�g��ҼG������~����Np�*�G��F��|zH�3��t����d�'��Lk�p���1�~'QB��A�v�ah�[����7a�yJ��ӻ�t%-�0ۘ*�
��>(�޹-�=yG�?KK��:K�~�� 2���j��Xv���d��=��|�8Z��F���약_��䋨��8E�;���I��|�j�+�����h.aC�i"��j�T�y�F�>��_qS�,�j�*9eG2ʺ}��-f]g殺���-�hGk�ViR��q���~�l�_��WX^��"����{f��h������ԁhQ���×���uC1���������������6���<q��L��TZ�r��|�&�ҫ���|}FJ��T~KȪԅ�_��H�-u�x_8Fg�<�2���Y �CW�tnO�HZc������}XD���u����M��r�!
��pi��R�����{Q���
����ک5;G�d�Ƽ�'Z�%�����\��5B�P5��*J�{�r���N��J�vlF?�/>�V	��Rf��)�2�RX-���}&�Ө�AH�t3�����Q�/iӢw	wۛs1N���#*_�U�A��ڂ�ہH�a6H�^�Ѐ�}����Q
FQ�2%�c�T�������xD���#H��H�}C��K�ܿ<�a���-�0K�#�����@PȖ���B&�����A
�@g��~�^���XR�E��Z�'�=�8�v{���Y�^���"(���2 ('�a�7�ƬR���r��9���s:��<�."��ʌyP�mE�ۃt�^�g����y~�H�ヤH(3)�k�9E�J^�l~O��'z�?��v�I���LJ���<��>�?�k���U�m���pцpbV �#���~hB�t#$etU�m��r5l�l�5U�v�(_D{���q�����7��˟=��2T�d�s�K/٪7ԓ�^��� ˠ�?v�jץ��)Q����,�ͽ������8��9��q��v���H�͖҃0��L�-Õ$7���()?����n��P���7Nn[igx����ȡ48xm�ɴFju,/RVu�0���{k��̙���?��И�}Q��ے+9��_t&�O?e���K�)Fa"lx��&����P*��e�����"�U/1���Q*j��0�Ö��"_�ֹ��goE1
l�P	�ދ�걽69�щ��	3
4����ﭙ)�U���T��H�dҽcͺh�C_�t����,�,����4��)A�f�=�d���\���x9	tWU����h%�p -<��˷�7C@�f������k7`ڋy}�!󃩊p��窅���V�LO�6e0���V� �*�Y���0ltδt��74�ϏM��j
*"8Xkr�e�)�W{5�#�+������M���Q0�mSZ��8�{�[��kܨ��h��N�/�;����h}Y�)_�f{p�o(@��������c88bUej�`o���|�,�#�P�&��9���|�Oe�;���4	�O�}�ẎB ��Ԫ]-.�Y���A��_A������2}rO=���R��&��g68l�6\�!�n��YJ�О5�q�t"�tܣp;�t�ctд����i�����ԏ�
0v��%C��	��!}��)��ͫ'L��q�ɿs�����d�6#�4lr-�}�m�뮭������B�{��ON9v2������׀W��c�����.hi��g[��i"�Ш	�q�b�Ct�
��s�|�A}(Hs��(��p�R@��ړ9BӠ˔�]�`$�-�K�C���;ɹ I�;P����x\\Ȣ��*,A����j'�(���N3�3֑�ǣ�jF���]H�&�聪�:B�I�
9��L��U5�.�F�%xD���1�Y��A�۶�U.#�I/p����D�ף���B�JQ�C�
<�/�y�����ܤ����|��r�:�~z�G��_�MO�K�m��i:� 8θ.�FUo��V�'^�ꇩC����9�UM;���^{�������˺�E�Jmh�5�]��}�{#(U�1\N�+�`~�1���~�:�SМ�B�>��HاHB�_�uЉ%�1�>�5]�w��rHD�V�c�egeI;�/��6&98E��b�e]q���H*�$ѱ���{I���\�dhI4���O |�ś�t�uӕ���	���u�Ղe��.�?�ڛ;�.	j��!$f ��0I����R���[�#519W�/��]�<	 H�[fhE4�Prs9"J���F�B�/��|᭒����an��L��
4NV�(m�ݗ�:s�xU�}�쁆��W KK � ���ޯ��['>��9��:��_�VV��/�Z_�EYd�M0e��]A!/�m_C�����z�m�ҽB��Z���q��(,L�ˉbj���H
�������B;��0�Ă�Y��p�=e��9�
乞1:���X��lj=��L�IR����q�q����=�����Rah�2I�k� %�h� ~9�)�������aQTn�)�P5n�~&�d�F�y�j�>�D����v3��،�W��C%��p��Kn�K��\�a�pY_G^�	݁;☽�{:���Ig���[�;2���St�jA~��ld�G�Gd3--z��Ii8�*�
�t�
��.Dؙ\[�"?�Y�#&M{�-�I��V�܁Y#����G7qDc`��{�l���e3��(��9�?���A�x�YD��� [\�8�à�k�ӂ���\ZAH�G���җ�?��3��4�HI�sy�c�P���aӟ���9���dx�%	0︣z'��zm (W�s�.���Y�a�B,6�,�3?9���`�PˊQ�V5R�B�w��#zs�YK�l��}A����*�'�=�Ǔ~) ��AJ��8����q�:O
_v�bK���<,?^�.	3CK�jQ�<�41U@㥑���"n�$��9]�,Zy9D��e��>�H7��J���te>��e���R�T������ٓ��ܪ�P��ɾ���v+�h|�@���Ѧ}���2rΞ�>�ͨ�Tk�h/G��,.���p M��>����8�K�}c�H��i�JuO�p��s8�x�f;�E�&�dj!1S���j�q�p\�Wd��F6�mjsq�&��B��{�������X�ڞ�<|������.OY����xL聙B���w�T�0y��37��ƚ�60M�Ӛ,ݢө�
����Ϗ�G���|�����;QX���}B� �[�z�љ�.7_A�03�e�ؽA歚������Ƒ`SQ{Ԝ��y����e��W�ˡ>X|��[b@M�qg(���FC�i�ϟ���v���@T
X�����K�-��{3���{�I�$NT n�,�qV�����X�QO2��LH>���+�&���k��n���`��~{Z"<�y]7�2v�p��مx��EDG�P	��G��1���x��ʷj���Ȣ����Sg}G�8̃����̪�����|�i�-�"�D�]�F�S1�F�Ư:�5Q��Ζ˫��R���a�aB;�{�aO?mF|��P�u516럧��}y����ނ���uv�o�E�h9��6�yt�[�2>���\��ug'*3�{�b�@���G�76�e��<�t)y4}Gg�~��8��IͰ|7���V\%�W�qЙ��q��M�~�A�1bKu�SoM���M���TWp�緥��7ƿ:�nˡ�Cjq�(bͨ'Q���J����5`����Â^��y���$yA�l�S��jc�Q�8�u����21��wQ|Bt�k��8<�K��
Ouj���IH�7��]<E�sȷ�6��S��_�[}�^�E��:.��tL��QD�]H۸n&,-����g۱�:��J����r0�4ohQ�u�?jO��Ҏ�޲'��I!�jE՞�r��ZZfsgc��aF���Y���n��E�8�0L\7V���]�����:E}�]�&ܨ: ���ǌI�x��Yi>��r����[SsRW�z���L!�9.zܒ�Z%,hFk����9�s?d���`��.�rSl�����O�ŕ���*]߁���I��8���i<��Ͼ�0̱�V�[�9�̹I�-�e�SՁ���]>��+G`(����Q։as	�I��_�L�Y�h}VV|�T��@�B��5�f�|���b�l�0,{�.뭺߰�c����?:T���UJ��i�ȑ�gĔ������*���d-�Hw.�e"Y6ng���p��.���j �iz��zwr���o"�N:�K��ɔխ����1��&�a��n�r���ױ�:y����fU��pU��`-��';�-
���2�.{@�a�kp��"ϡ���8�e����xP��(M�,Y�mH9k=�K�����<Z�b}#���j���t}����k~q��.= $�˧3�
���z��I�Z@��R�c�E��t���	�I���H�џ��e	����)\b���^<�/�dk=�
���:n�|�����b������o��K^?2�aaq)�~�`=�[�0b�>|���M��5%ǈ�����s��H��Q�j����c����[�C翷7�G�6�SJ��.f�c5��?FN*�D_7 �f�D�Qt,a*��.Oºi5�/�T�n��6"�d�38��J���5��/2٠"��Q�1-���y�c[��d@��öF��9C7���@��=��_��ޏ����J�I�c/��i;���>�.L��yT�15��ܴ-�.t
�%�������L*�>]�d1�H��?����!�z�x�no���|�SPL�=���I�],���Y
���?����/�C��J��Џ�(�`�5Gjg�>ʁ.�np�Hݨt;�^�A�9gQ��Qv%�D��Iwt�h�=h�UP�r�����ޯ.>���r�\m�H)��<�����UY��-�S�?iA�� ���@8�sL:�$0[����Y��[�o
f"B�5�=Jg�eC��A39���Օꠖ�ݘ��Rο�ag���q�8�F���Bu�	��j�Z�؅h*ܡJ�;�y�w��@�s�r�5���k �c�?�uW�R�v�|lG�xy�*��?�7��j-5�59dT"s�X���:)k�m��
�T6��Եj�J��  ��@V�o4��;�M	uZ�Xe�^k��R�$(�M=*������[A��(.���t#�;¼XYݧ��O5����'#ht\�n������:�����Rs�->��4�s#���M�(�y ��H�L�d��?�7�϶�����22"c`ؙr�HAg���R��P���w8Yz��<xW|tD��$T�A���w'l9��3�k0dyy�3N�1�A9nP������Y��8�rqrX�����-�G!C�ϝ��6��6Iu�X��~/�(���Bq���=��+XD�0�%[��b�Il����\J���5t����g�����K��b�����-)��d��<;�C�8���y}���s7c���C��0�Y|H���!2��w4�9���I]�U�Q����"yK�ڟݪi�"��KH�t�8)"Q��|t9V�A�)@�_�j]��3>���kISձ3��}6x��E�@�=���|����<l����[��H�U��.u%�;q�C��S���2�����5yo�#�M��p���{cV����+N�P����y�?�J�Fn�H����tj��T��1�O!�����>��`5!�r,E��!��E�oC �/��H�*TL����0��� �ϝ`���_��ck8O�c��Q����/�Dsw|$ҡ�&�T�/>t���b�U�����Da�u��;
B)�ձc�6��m˻O�m��#%.�T�8����Ww�͂ն>�[��icx58"ij;�??�y����.���p5ɲ�2J��L�e��ژ.:�(/�
������
��ذgiJ�g�'��Uǲ+�3<�ރ1�hϗº�-����:�y\�y������A�w��-�8X)A=߬`;�ҢԀ6���L-M�����=E�>��ݬ���>��(V|���C��l�����`���IZ�!^y��H;.\���̚:d�%ȟ��}�}L.�ƯY�e�y*��V��3�_~32��7k�/�ʾ�Zݼ��g�1���������'�n�Km}4�1}���Ê!y���xf3���^���Cm��B�=h(���R��).p9��]0�H�>�,������"���w�惻�pt#���"x�9TC˧�ۍQ�f'?;F�`�N����<|!�5�h���� ~�{��Ԕ��[�1�|
^��zɓ<�q��@��]�e���x�M�A[�`���1�Jq'I��3 �c�C�q[�V�k�:sō�\�z�}W�]�G�0k�G�YDUǌ��t�0/}!�:�����r8��1ú��� �&��}�!���G�L���}C�y_Ԍ'����x��&�Q��`DOI�c��3�#J�,��[	%�_��(�O�_w��X(-�/�r���2�]�/grB��~U[�M�&D�IW�c?uw�թ%u����1�\�������&Fi4oW����ۘlSI��)א�<��]�&;�P��`r��5����5�K��Ω�ԫ^��Tn�K���q�|���gԣ �n��="���)�״c6�dk��^�~��z��m��cJ֗�nM��
:W��ݺ��&�
F3r"�ʆ�qÐ�Y�
���:-���p��ƍ��	,A��1����3�^�0�����TRl�����'Ca1����Bh�'&n�*�mP����/1�C���O��7A����0�m9\�`���%���|�S\	(X��ewn����������j=��B����`ddW�$��ө�(�}&#�S�D�w��\��챺����I�پ'B�4��z���ԠX�K���@$�'����q6-5�DF����-�X��_bw-�=M6��>���֩ԓ"A�_W{YO_�/�ύ�-5��j�?�`t/r�Ȏ��2M��� �7sנ+�gt��{���F]J�� lb�� �Se(�u�3�� |�.������&�T=M���+�A�����V���~��`��+�sX�QXQ�v@5�/ν�G�)�|�C������6nܿ&�$	���j��``U����
��5��P�C �t�S��L�Ԗ�RIB����d^�� ��~��ྖt�}_TX�2bϵ���������vw#ѮE��*�d��Q��m��?;y��q8Ë��eD_8O�I���b�JW�Mj��='����r�GI^^	D�v�ɬih_���b�1"b���&#V���?	�����3l5��j��k�~�7�_(q^r:q0z�x��$����:"��[�� �:�i��v�椷�nL�/d����y�	�l��$��ם��-���k=�0+����0U�[��\z�Ȃ�ʏ_v2�y�)wَ�OƦVs��J'5'�x������|����5vL
�ޝ���#�ד@�;�FO�]@�"�Fo[����bPmͣ@�9����m�E���[�[{�+��J}#,!� �<'Yv�ߛqqH���o�kH�$c%����ߓd��\�4Pb�@C��h�������ȑ'9ׯ�lhQq�zj�-/��ԥ�^ղf_ͱ�r�.���qƮy�jG��D��6XH���vN �wLN�XR�������͢�E�%�E]�����N}��G�+�DSz(�NF|!EHR�zK�X
S./��솄�@v��)ݹ�Z�陵7���K[�w�yF�_z:%8ךX=�i�8w���=���;}ɛ}h�)�A���U�^�0Sw���&�=0WJ�1����_ ��K c�
��k�z��{"M����E/D�?���m�h��;ξ��Ӯ	N:�fG�Á!8�N����%#���9}���`�g�3��7�q�"���q7����ǧF��tV��[<4�J�>Z�Ȗ',��.�}9��!��w3�Y
��
�mC�v� Xy�$t���{��,�j\zx\��p��1O��Ê,k�x�TY:+����G?��z�K�1�����r 1�[:0Q�r�>��Κ���RC�xn<�w�������1��S����(����, ���p>ǠD�Ќ�y��[����(>� 6ZHv��-D=�P��������ݓ{VϚ!�+ �����8hŤl-wrKh��CNHA~f�c��][Bp���>������0�r��b��S �:��w��u�r�{E��l�@ �<mZS}x�����wi�|��^��Ut�v�~s��'��;/Á1kC�eS4Y
u���"��_V!���]w�koO�@�]�$��eF�ß�K���<�?�D���O|��%D���D92}x� ��60QٚNi��mX��ǜ�d%�o��ȋe��Z�ÝW�rc�zz��l�1c�͏ҧse���ժ���J� ��1A��r�w`l_*}L�ei�ak���j�0B�@}Yϳhg_�$�uH�sc�U�=����פ3�l��D1�be9]6s�7ơ�`5���q������䊘~k�
7'��w��wo>�G��x�P0͞y;�/�^X!��RY2v�e$��i,�WR��cN�ya^:�a{��%�s�́R��+T��>dN>�9#�����~u%�h�ϟ��4�-�||�ð�4�	C|DM"�wb��1F�@<)M�3��u ���#8�t��MĖ�"�'H�r0"Ė�ꮞ������)W�u�~��4T�p@j�dӅ�t�5}T݁w�Ĺu�꛾���H.���v�݈/6���eTX��~w�&��&�~���Y�e�
޺�}ں�_4��>�f�tf_� ��c�-�*$��zG�3)S��IE0�q���W��_<w�
U*�L���-��w?L��t��y��-R�h%C"\��m�c<ᵜ��7f�>����x����]���v�]u�u��ų�B�E��Ė�w�~�mt�W˥����`4�G��*��ދjށZl'���0A�ě�\S�r�-�3�Hg��`&�`)a��������-N�Q� 0؇�ST(�%n_CCv�� �UP�A��#���]Zg��'*�!��a�?i�U$��K"D�}����2��g~Q�+���&��J����L������杄�L>e�o����z]1���{�����9�l�po�v  Jx˗��$Q׷k��;H3���D~ ;bϪy�]��t�F�6��oBfI��%;պ�BH�M���\� �J���՜���;��^�����[i (S%	ne���߬�Ƅ5�����e��<Q)�F7�l�Ƣ��La:��oʩ�.���F����L,����!1��s�r�Nl=�*<8� ���j.��G�q3M�Y7G�������ldg�a�G��ی�>�3h�Ȉ�'⤰����K��c��m=N/�g������dzy/�pf��L?�:~��wr�����լ�R�L�䮌k�,�P�zK��!�Z��/k1u�IV��!�<��Q�R�4��3���`:�p'�FJK>3�\��FC�>\i����w7#����6�F۽�x
3��[e�C�Y�a��j�!�:\����j��\լU[oBʛ�U�@�Pj�������H�o尫��;��L��E �6Gɮ�F�)�KsW�!ev���4��݇���Fe��{Zuv��M���2梉�)��UI%���6ۙÅ?�Uy+����P����Y��0�$v}���ZF��<&�F�#&	!�1(b��IV�(�e���0��G���Ϣ�� y�&+n�N���p6J_�n�A$$������[N�IB���[!�j�54@��lɄ$�ƁB��P m�S�]"۳��;)�{�h<j�t���A������b<��,8��Jxq���cH5t�1˙
�xDD�������Y��Sr�����}A|b�����U��sv�<ӽ�#t�E��KU�7_��^l���c13~�@Z�V�2I��G`�L`V"��~Ǐ�Z���?t晸����_wO�d��;���6C�$����ڃcy��~��ZQ���2���M-''�ejˎh�h���s����r�����l��3��� ���
��w�b�d��H��O��<l�|�,��ջ+��O��N�,p�����р�uGb�6I ڍ����i�r�/�����[�0�!%�e���?<F�f; Cg�xU��Kdj�����*4�Γ�!�\P_~"�Q6���yr�p�|3�W)���7��4��y|�#20z�t�}��-��ۯcq���X�yL�*�&ddz�.��,e��l�8��H7}�"�n�o�%uN��\t�Wh�����4����`�r�9�4u��wz�kV?��s7��m��C���1O��A�Zq�m�J�	L3��󩓎y��a5΍���K��Bz ���_E9�I���$�$�%�yɦ5�4��}�kP�X�����t�����<ӸA!��Ԭ'�{fO��T��E�	��mc�(��)��X����Ruy�9��qYsD�"�0�N��	,-n<Jag ��(��C�p��k�H�\�	�AL$0F�^�d���}Y�$t�ES,lD��D�W��K��0C[r�xoY\\�p+F��q�Ȃ�n����<��a]�I��/�&`�k�di� 6�T|<פO�@u���k�U�a�;E&�,�)C�A��OO�XFf���������an�r�#�FwP����&(D�������%^H�ek1`������0#�z�l��1QD!%	���t���u>(�R������j��*� ��y�(�,S�0i�@d(4L&�כ��f������~,�u,��h �V!���ѺaR&�l����@O���}�a�t/��F技�Z
�n��h�.O�u���j!������CMdd5kܟ��������5��S�ˢE� 1 ?R&��M��g>ek�/�:2Ga�ǧ�C�Q�v�%�<9<uܡ)�߰��r��|�2ޑ��Ϣ(��:ޥo,���0����s~�C���j��[C9�c^�~��U]=�xƽ�Y6SX�1�%��G�)�pUg{~I7����T�u��T��ہ��%RaΞ��oz��Z��}?�W�PѦ,��nB3h5���K͏ ����5R�|��i*�?BQH�D'c�����o�aN��8��v�Ᵽ��7��W�C�H|[j�2-�9N�9�,��n�<�9N�1�:`{��ah�[�f�:oY�5F�F�Y*��蛓��=).�ө 1=�O[�`�b���en�j>��y�$�PՍߐ"�g�r �*�![�օ�����yVp�m�P��	j~�ֈu��5£��������E�۩JZ�5�qe��1z��j�%ǡq찡G�OS�]�`��I�4��Ш:�'�ҍ�[�'�Fu���>.�ҏRAISyhJU�Q�_Ug9�D���ER�BĈ��T��:=���3����&:�\ZC�6�m���vB���		�h�/�=���kw�c����r�B��Xj3ȗ�E^\a���<�����
xߦ�$w,��"�H�R��?s�x��n�C!� �r��T��DܸU]0)?yǐ���!����G�fJC�6qm�$| ��+8���_p�*w�}X�r�K�AD�����ٚ�@��`Q���:�6[���|`?��w�H<ce���I�L��i��H�m����M���R���M���Ң��N�P2ت�!`���>�X�']�fθ�*�A��x�&ibȬ�ZlS��!���� ���������s���2�lє��9�V�&�ε�7��Y���ލ� R�0��!_�u
� ����Ο�Ų:�u��X�����Z>B~k���l(�����O��sv�Iջ�NJ�?o����f8 ��p/�6��,5ƭG��'!8!h�X�P�	��������9Vtvdt��Fr�Q��s��/iA���@5)'�<%򓣸���R��g�xu����e�HW�@��BF�(xm,���"ەn��R���Е��O8Ch :
9��o��8�����2�Z�"�1�g��AR��w�1�Hx��q�A�^�lG��+B�oh�6���ܹܘ���EH���9�w���V`�/�
h�^�w�Z��<�����'����p��������M�����xCEu��"S7]ډ���x�o?��w`4��7��m��N�R4k������~�����^_B� j ��l,f�RFE���9��޸&i���4跨^�dX[�ȍ�*fnqU��;'4�ZK���MB#�a��1�b�l3���.��U�}���^}غ�DF�B�ˋ(��K�v8/D��+�+9I;�̅*�ν�:�n �v*Z=�|x��ox���>��p�B�p���w�)|��sQ�J��ZlKY����/^�V���d܃J��Ƒ��<���G��<��VFA!E�?��
ռI�vp����� ���SM�x8��q�tx�;��+�rTm*�c�$�
Lwݽ�"hq�EHn`��|{}.�w#/�ˊ���B�[�+������ �3I��3Φ�B�>���z���T�#��_���5�A��V����ӥE��c�A:�HMy�����h��&����c�?NqԖ�dQy��������.h�!�/<�M�� �� ���q��FVy��U����S�)F�=����lD���a�(^�+M
��/Wi|�{�~��E�K��Zk=D�3-�Jn{�ue�Nנ�
�h����_CY�Q��j_]�>�3$N^ށ�}� ~��p���G�<*������8��mw���i�@X]֧?x�&M��p6�w���J�}�n�p{	�>��r߅]��̑��J&������<�H/�o>vf��Q��һ�ïR��o�j�3:1M�b�z��1��\! ��{Nvl7�mJ�	�b��CzP��۱����Ë���z?�
�n��Q�?�����m$W-�_;nc}2a�k�*����$�T��B��.@�ʫa������|��(2�F77�T5���o/� x���g�2��0r����cY�v�1�C��q���8�B*�u[/����RZ��@��>z�g���j�Ǝ���`'��R�g�2|m��g�E䦭�<��NU-���7���K�TH�E�ʱ3�?0#:BN�Ks1$,^��H�ps/���j�'Z�]��)kft)=�ٍ�ꜷ3*
�����*�\l�	L���U����ɎwA-� �\݊��Iٹ�m�1�,�ɷ��PP �u\a*Y�g�z.�w���v�V��U��p�>oN���'����" v�e{��]�!�*�O!_"쇭Z�/P�-k�w6+�ZHm9����3��
�%4��oG�᩽�l����<!�{,fN֨��:���V�D���f��I��`�+����d	*�k���5�kI�A�6"���a�[� ����oy�rt閹�Cl��m�׎^�3Yk��qnJЛ3��	u��w
rQ�6g:��c�n�,��9��}���&Ҝ�qW��R���![�4ު��P���eܸ+kyQ�e7���Mn��4X��H�fPBIـV���Y�������j�s����nT"&Pe�d�L�PZ���۸������e�|���4�U1��4fl�{��h����,�<��L�kU`A����]f��XN.hR�~����0Oǐ��x+.�%D�dDK�>�R8H�c����;�ߚ��Ex�&�J��־�����;X��΃�Q���=���oӌ���L��C4�{���TP�������8 }4�n?��P��o"b��ص���n�io@��)yǩC�m��X��CU�i-����sOw����ᾁ���}x�Z�Й3����z5�A�ˁZ�0��P�o\o�
��`Z�k� tc9�'���GD��8�{��o�?f�E��ɈI���i�k���X�풻�hR�ݺ񜋺3Ϟ2����2-n	�6������f��p���0�t���K#��t;�|-,5^tq��¹�s���:.υ���+�"���S�	(8�ȟ�ԇK&��,��"C�C41|��r���A�o;Ē�b*ҤO�?�n?s�.��~o� y�A��,>V�X�M\Y�I�4�WeT�Y\�~�5����w�ox�I�����⭃����MyK�v�'c ��N��ulM�weS~Al$"�Wc8�:��>�$�5u?+��J�1O���ç�؅�\q
��p���c>|H��ԝG#�A��!��ͷ޺W"���vۘƅ>����e���> ��:��@�h�bĜQ�����k'���d�~�G>z2&�k�m�⪝��<�9��W!݆w�a/��^C��\0�!5h'�J���o[e3�@�����3�,R�:L���ݑԸ!QL�db;��sy�S�@n�GJ�fS��o��&Dp��� 5��Zm%���������H�Ƌ���m6M��rTBY=]���*��}�sg!���Fl�_dH��׼4�Fi��S�v>���L.޶���<���9{ŕc�B��6�[,9�s�`J����O?�W��{���E�D�KבF�	�n]Cd�Qw+;�)
�}T�[Av�Z��=�c��xc�=�~��x>ćJ�]� 0� ����)ݚ����z�#E�R���·	Ukse�%
D�=8���4�Re6�u�T���(��`6/x��)lh����wÍ_�}��,wp#�DL\`���������v(��pUoP�MC.�L�c�=T����.&�(�.�:�v�~m9>!�<�c0߬��P�7���"��J�1W�'c�0÷�?%�����ʪPv�=bf�馎��O������д� ٻ��{����3���xw�gXPZKęo�=���dZ�%h�ĳ4�Q��g׃kb<ܪi���o�f@�G�b���'�"߸����`�pM���i
j�FPS�m�_?^��Աh�]���|��'�h�.���>�fx�)J���H�#Y�Ѥ>O2%R �R������������0�c�0@���E̓qkG���nB,��h�%�?_��s/�b�/(@@Z�̒ᰎ��$�S�il��NO���ϟߐ\���rf�[x�����!����(-v��nE��גr��;����V�GN;�e/>A�G%D1�ߤ�ĥ3�N��K���t��P��V�X�����dib+UD�i=�:��k����wˁ��%"���P$0
�8�Y�W��;���3��T�H݄j�g*�� ��k��޿w2�.,O��r�����o��j�!*#�x[�W�]xtDK���V�P��Ra/uŴ9�/�->�o<�4���r��M�X�*e�U�7�ݢ�E�}����>{{�'��ғ�M���R�vB�Ay�<�*1|p��<g��V��TC�E^K��D?�����.�Χu�����U`���Q���-#��D��4b%�����:�N�R���9"5�G��"��C9� �H��.�l�.��0��	�Whu�?�i;����6�9���3n�e,��&nuQ@�\�`T�ԅ�eY��7��0�&��)
���ԏ��4�`��#{�{�0 ?�85�y�=�����O��0�㴩�i���������\�7g,�zm��XRF̸�UP��6����w&�#��ƿK ��z��R:◍�A�K"R�UF��m]���~Jضh���$�|�za{N>1&p��@�w�0�ib���Dq�~߳��Աf��f"}��N��}��O�f59*ꔣQ��N�*)46����ߟ����7͑��V-1��18I;a��YA[UZ��QAI	Bi�8ר�ȼ_�$�2�Ȏ#S/�)�U@��S"�B���< }e�h>:�^��=�\F�}i�6��FՊ����NPw��7�N��M���⿰C����f�<�����&�d%���Y�z�:Tz�<��UϦ��_F �ӡ�-��ę�[آ\��Yմz�b�1��-��@/�<�� �`eX�fK���-���4�MH8)�.�G�>h��%{�=�t���oiU8>�Ctf�P��-9`��'����I�JW���O��Rk���-�յ�h$H�0X*��O_KV�|�v*�96.����T|�	�H��|��x^`�%%g��=�r����;�Q�]o5{���0Yr�`��\8����R`��B�|��7ZNr��y m���gn�����/�+Z4�-=�`	�A�b��OR��HV���b���1P��E�((�/}�Rs�S�8�?.��e����)y�d�f�e?M"��7.�B��I��H��q;[3�v���u~�7�H�m4��&ES��JZ鏻L�y�e�;=�d7��T2tJP���#�1����^�n*D�(�SN���a��W���7B�PIjkCK�}GZR�	Ag*��|�q�Iw#˞R�1�����r���]�	o1[�.Z,_Ig���>ήe�m+^O�9At8T�<�s[q��&�7�!>�;�]MC����il!{	\����z,��5����"�z�X,���Ij�L�G�Eev�Q��n��?���,�W �`�Tc�'�@�ħ0�Q��4����R%k8�z�K���{|a�U�KW��k��:�73�b$��pI%Vw��C���b!,ZD��/�u���QŦ����%뉎�=�B�!��gz��(��I�J ��ڇ@�m 
���@L�Y���i��YñQZ������3�g��=��m"��a1LL�'~*�g�$�l![�����^.)�xeG�,֡��l�i\�p��K�i�j��;���6@&�J���ņM��=+�
�nn��t�W|���a�ۂ�;&Ɨ�r�aܧkQ�n޾wX�x���(����_�9L[�%��5^�n��5��	"�5Ш"�fP�_A�lL٥�+���o�h,O��[�wj�h3t�X]����$�P{�����-e]��Գ|%�ll�oـ��fk�k4�=��'&�X���~V<�M�1���VõD�Ar�^�V����Ȥ/�7mw�k�jY(�iȵ�k�W%�e`}� � ���rp(�5�Z� �|�$�����v^v�_
�J���S��~;�>��u�ghE���
��A�0��#��.�ʵ��ڼnR��x0�<��]�ZяY�;m���W���s�PtFѕ�-]1g����ADr�h��g�GZK�N��!1'�Gˏ��?@b��^���1]4(�u�+��;�!�*��.[�]��Y�������\�%c��WX��sZ�&��2�ȡ�3@/�����a��z����.f�jO��B�G���8iCD	s4f�z�
����3'f���u�/�g'a�������H&8J�N2~�����Lm�$�p��GLJ^�I~m��E�<7�"=��TZn��nR�T��x���鿇�n��n�o.��e'Æ���̬m����;�N6�w�ʰ�`��_ʪ"6�k1�6X�p��2y�(�qZ/_v�Rlh�^|��ԑ�Fe��f�Meμ���b�kin���l�a�-F�	��Ss5t��x[:*v ��}��*T��>.%HF�~�XIU�M���XQ���o�Y��M¬��k�$�M�!=Z��^4 ��D���v��*�CW\;;��	��` ��v���zb�hN�=v1}h�dA���n
UY]�=	���/q3jL�t(��5�uYJ|����.����5	g��A2�B�3+�w�g����O��;ݭ���_�|@����@7���bږ�������9;S9_�C��hb�� �â��K�%��,�1:w��}�GP�ކ)|��9��.�'��+�hV3����{s+^��k����]��'u��)�@!l�K��-�v���iu�fVM�6��L��ښ��1i�oTd��"���,ǐ˰�zf�����}UТ��U�b�J�rh�J�]��<8A�\�8�*���:<ǣ3z4�>�K���f����-��o�HŶIJDԣ�����쿫ٜqi��]D�I��0ZL$JXIi4-������D51E�'�[��0���L�>���������9,��"��٨%~Ok�}���n�Q���:x{I�"�M��E�^v����HL�+/�jMZ������BS��|j%�j� ��Æ	��n�4�e����p��3\:��7 R�jf7R��@k�pJG���?dV��u����s�9��2]ыX����D���4��˴�刐��8��"^MBg��`S�:�*�VD��%�Z���Y�9�H ؗwyN�zO>5�
���C&��q��5��&
X2KnR�N=�{ߨ����DnYG�I��ų]!�'Q�q����,��4>�������)�EeN2\:��Ȝ��OhG�����*CXч21��7��ʟ�{��� r����kD���`��
��L30g�?1ͥn���n���*�!�����]u7��ɱ�$��_��X �,�0R�YO.��l�5�*y�oH�0ၪ���T�g�@$�$��TQ=B��q�8��cvhs����B��n�4�3�`K.�$�^.�4�/E-u�d��˽l�P��6��܄��3����� lC��/j��6�����D��rc^i�<���	�P;3�5Qg��-!��~O�ޘ\�vEv͏/��^%��f�=���SK)�C�� �\�W���uqC�c�$r�@\Scckŀ���USQ~u�7a�(Ėn�A!B�g�0<'����{]м�SLz����RH~I�/7ʉRO�.�7������c�E�Tb���kG�P�
\pO�����C�H�=M~h�Ψ��v� "�n(a�|�Y�bA��@�H�P� �<y+�L;��y�zj�F���~�>�t�͗���h�'N��#��_��ר��B��qV���JL��g{;S� ����%�m��,6H�L�ё��@��ʢ�W����#�����޴��~W�������1d������
��������*�Q�~��������x����)ߛ��>�1$�ؗ�K���#Y��\a<�H�M�KDc����8H�K�O�m���������#S´xf^z������鰅'����_�(a��}�8���J���ЮP�_�i������k����SF����pg�Vm��QM k�����p&t�|)1��_&Q�
!\��WO����+J���?п���Y�'��ym��,Vč����s�t������1v��q�ΐL
���O�>�$w��ú�O��X�̇��c��M��n��LN��VΌ��jM+;La��8Tn�:M��s���+�bʽ"^�9�x��Ě��
���)]_f4�����&�En���;��>��	�%{IM�m�I�:C�T���$��43���w�i�ܿ]�kTևb��m��	��j��_c��"�����w_��+r4ul���|���`l�Ŝ�&2� ���.�9�&U�O��_3E.W��5�ܡ�@�S�� .9�P��n�H~�z��n>H��ľ�)-��_�߳�d�����DĿ���Y�"���SC��@�t�'uH�VIv�'m�
v�+�`�DK�A{��R7� ��g5�1&Vea����-w�K�D�[�����qK�s�#��k��+�܅���,�D4��k�����G��j����崁���'�ٞ�	�j���.d߳���r�b{]Ǒ�)
Xj��Y���N������6Ĵ������%�a��O��7�Y�a�u�;Y��?k36g�B
~��L�*ڈ�:�K=���峨���#KQ�E�&��Ң�]#ΖZ˒��!ux֒�@�$?���a�"�#z���>_u��D�b���Y��=4�겨��v��~��Ѿ�mb_ǡ�o�41� ��|)v(c)���K���/R|R��1��ZJ�>,�������[>Q��v#��daZ(V���	��=��xM�`�Ŗ};;������Q��D~,���,Q�3{�1���R����/T��hǮd���H��v����7Q����o<���Q�#�a$��ڪ%�@�L�+	�c�>��_L�TԖ�ɃFν��"��!�s�6���邃��{�	�Z����R쳾�n9ߕXL�;��!Q[ə�T�I�R���#����2za/�ӹ"���I�G��R!�5�p���J�u�v�j7?mv��\������2V|k˔��޸�0D?f��� �=)��0��ajH����
Al�E�n�Q�����������|�+�_ ~^���L��w����WP�E/���)��*�B�?�t�Z D�?�TT�yq�f�B�G/L-�0���X.[�sh
�c���k�L�q#N�e���Y��#zo���:C�]@O� ���Py�[}����Su�+DjR`�CC�ɓ:�Az����3{�겻t"���K���Al��1�MWc��$��}E�s�h�~���Um�ЦYDH��L�w�m�(����3գ}��md�5�z��n�|�Ea�j�qB�H�6&;�R��Kz9��3�H���.��*�GO�L�oc�r��Ӄ��Q��GZ��D�SU������~�~T�+-�d5�%m1�MJP͗gU���<��Ƙ�T�*�T:Hv�S��4����Iබ��8-+A(�s��<�]/�Q��eW��_b{����J�9MZ��|�r
a�L�;�;H\����k��|P��u�?Eo�>`��T����46:һJ�֞��7g��{��C �9pd-_R����>\̙[��1JN����@r��a��(L����4r{�2~E���D�X��e��?��>E�D��sŊ���Cz({�x�D>WR3��ᅣP����Mk	� C����v#�z��Fft[1�``J�㼿T}�@$�/ѭ�=�40O���Q��*���g��`Jq���H����}�w�EL:���/����|�D���̳��^�����g�,5�ow�e��f�DT�����Q��#�(�Sĺ�ƣ�� �c�1 �@8�J��E�J_6�����j�&x�o S��F�^�@אE����דD��?C���X�m����{�Ӣ�q_,����?�f��"�=�*H�e�l�� �7H�X���7���yvr�� �����:������rd�	�d!`67�9e���4ˋ��q���G܄fs1��
�M����F�z��4��mA��r'����R�ciW^��������Ov��"�W�+���+��:�([��q���9� �6���_j�¸4澳���\�g�i���v���������g��/;&Y�{�|G��$��m�&����d��^�?^�\LpWH#�9�n�k`1�Q����ԅ�����V�x����p۲���&��D��1m;D��ڶ\$�71 �q�WE�A�ڒm��G�	��Q��Ւ���ԒXtmv�2���IV�H&\�t�(y�͗��T^�܎���?� �����7:���)_걯��0�sn�Hd@�L�^��tțO.��m@,��K��Y��<��7��H�W�Ě���z��D��������?��p�l5V|&;,~�v[��ўS&�z��/�'��!�(o�t�i��P���\>��Z�����Ӥ����I>I��3QS��c��>E����������yD�?�ؕ���K}�ݬh��m)�<�:	�9��]utn��|�6������c���`��5�\u��E�:�xZ*4�F��b5�{�2��%_�F?�׼b����D����k�;k�-��P��A~����{®�� o^�@�G�x�+���+��;�ߛ�VIk�Ø�~�4m,I�����B5�^��l�����/�ҿ23ऽa4��9��Yc�@`�I��?�v6�37�L��y�E�������K�!4p� ���p����ׅ��qi��,b2\\K�nC�ix��
mb�'m�D3,��Y^'���wR;b:�D4 |����)�BO��.j��O@�؈%��lR�����9��'��A} %x�@a����A����*[��C��
t_�K1��h�5��P��Ea®�DT�Q���7N5��d��2�]��^��96^�jW+���'-:��U�8��I\G������jB"'P��ލ�@0U��7�S�{�}�CxB�; j����m�X�$�O��W��w�WI�Ń��^r�:��߲����� ����#6�(tfǊ�>�P0?��(p:i?^�LR��j�JRX�O��K�D�R�N��G��<W���)��G��Lo�����7��9�5��?BGN�_�'��K��Q"o�'Lܘ����7B���H�*��J2	$�pQJ$�O8Gm��^_�U�25��z�:yݖ+��j�^;�&�/M���c�i�E#�;嫷Uy�L�փ�����Gn,��)s%b���C�4�EJ���/�q�-��S��Il{�P�No���>��V�\�O��*�c<R���C��]�����}�_� �^V)s;�:M�lq9!��w�!C�մXǾ_+{�WaK`jǵ��nU�$��2����FX�7�No9"Ď�7������aƊ����L0m�)��th[=
���E/���j��"��,��藳#M4�ڜد��&��	�Q���7���3>��8�M�oi���|���'p�փ�m��C�O(kX��ۦ���6m�R�1�K�P/A]r�F�>���6xPrLefզCG�����2����)؜6��ћ?�M�L
:P���T�����>�=�,�;�n:UR��aU�-�e]�A�P�O���A�&{��JZ�p��?�X\|��������ܦV�eL����@��$�/���ټ����XHl�=	`��@�N+&9����g�MY���"z�]f%/�h/[J�֩� �٪��%G��JR�vȃKp��{�\^vK~�H�l�tY��$����U�:6�U��"��TAT�3Z�+�\�H�$3 j*K&̓Y_�t?��a��q3d^���52��4g�Ca����_��4kV���0��M�]:g��&^�Lkl�vt>���ϓ	�x^w�u�P=����Ʌd�~���������	��wRn�����XÆ��}{��4&�WMeWPӓb�Xb�,�K4�a�_V^�A̬����4C��W��&?[�KL=ٗ��ف,]����?kY =�=XCƳ�z�܈n�k1/�XNR�|:qަ��ܹa��a�F�Z�&/ S�+�r#P�8� G��nD%۪~�G�Qz�W F���p�(�c�z���G��z����˓��S�8*��f\�<����W�N�pۥ���p�cέ�C8��Ps0�8�o��?���n8�����cx�鬾��N�6�܆a�E�A�Ak7�	f۱���";qb6�a�J��e��^�]SF���O��|!�RK(���n2lü��Cm#у��k��;m��:Z;�z�Y݀��=��>��t�i���)����{���k��/yX�T r��	�������<��,*��0�S>�suac��M��t�%}��KXC���{��9yq�v����̈́�����Q/����¾�=!�L��������dA)"\���Z3p����®"���3!�����Ai��B;��+�ƍz}��<�G{����	�	����$��٬b���%f/��a�J��a﨣�x��Ę&��cw�K�bk!�!i�KQM�B��t�;�q���y�D���W�Pj,EW��S���1tƄ*e�p�jy� ����e5����,�hn����P\��\AJ9���<�M(
��L��|k!W����E�O��P�z��p�!ܰ�9�yml�$� A�M�0{z�i\�s���di0dxx�<ɗ����.�W~�9g �8F��<��"_(C.`S��폤ҧ����~��ً{��J��,Ep��2���_�V4����G�\����Z�U����4B�*<h�#j��O/��/U��kSI����8�sJ���p�jz+�f&�����O��vh�B���I��v6�φc�]�'��Z�A[h/�����%Ƨ�����q�:n�%�w��J^��Iֆ���^�%��2�	�}���ϵ�eq%���[}v�d��c$Y�u�E�c�P�8���i�v���E�5:��4�C�}�QP;?]�"v�y6��/����}��t����E\�h�9
�:��D/)u4'-�\�
��
y����[A�Հ�n;_n\�8S'h�5����b����`��%�KU�X���j�gq�Q����].q&������ڗ��BZ(���퀵[�7>�E~�o��,4@f/�=,*st��/�L.s�1y��+?���(�da��`d�F|ws�!.�Q��2Y3�h#ܥ�����ɿ�U]7��jE^(�}9�ԯ���E�'��{KM�FX�"�S'�`��iK��G��S�h��g��x@	�x��NI=7��ڄ*��L�t��l�c��f�$/ͦ}ym���}��%�Y�֮����^3(¨+�hܷJIѤ��b��_)QW�U|�N�5��%������'ڠy=�d�z�^W|E�]���	�S&A��9�}�qBm]g5�^q��i=�q��z�O�y�H5�c�m��	�t�1R�"��ֈ6�=��/j����z���n�뮱$��OxJ�u�o�����Nn���ォ{?6,/ P?�'9jzFw��}[���^F̘���[��]��}tk�,��'�+�ﰷ
:�Q2
��{-8W��]鈸(a�wye��v�T=�n��ϙH�%�,:��H"��
�m��p?s�����}��^�Y�.�ണȪKk�:����Z�@~���̳̓�㉳9��_�,����m�dm�.�x��=��I�uMe�e�Өu�-;�<
��ߢ�c���: ���y�p|�	n(c6`��VkPЫ��ҹ��"'c�P�����]�����{���yߔw�ă�XC�Y3j�!a��M���<ݎg�l�^�G*N(;q��5f���#�:☉\�x�
cD���#�Z�W#���fc���rUs�ƭ�y�Z��.�i����f���t����Yf���m6dBz	��q��������(F����O�y֢�d"t2j.%�"�e�z.����J��c��&��i����X�p5�����y/�8��~��f},��9�>*)}���;M�)1�z9��Ecl�O��[��*�N{�]��k.�O�ҕ�BOPzxI�b^�^��j��YA�i���LS�#����ӷg�VĽ�?F��r��F���X<���,�v>�A�E��;�ǔ���};Ūp��]������pd�nc?�@����{3��gSO05Q�<#���^����Gܯ q'Y��#Mro��ƣ������M.�h��xe���}ڞ��?����G�N��33R(�yn,����ɒ`���2�^�˄nC+Դ,�>�hd��AhV�Y3��E��
����y�ݰ�b��E����8�Z�_I��μO�[�o�u��8���v�-�H涑y���T����gA5`EO�}���vf����e��B�Ϝ��r�I!� v*���[�I���������|7g�^��[nfrSk���Y���;��#��$#��1�
K�)��Mw���t'#<�%U5��V(|H��;�Z�>��S	�F�Z@*�%��F�0)0o��n���b�����bv
��n�����9Vjh4��:&(U�8�z�\�Q��)5j�i}�[8M@���P��gi�Dd.m�����嘽���R�����Jj�d���ݎ����1�>J������ xqaAPO]Q��FE�I��
g�c���͇O&c,幊��D���N� k�9X:Sm=�<��]���s���X�~7�j3��$�����Y����_z��Z+�D��_�)he��^��O70����D�	vRx|y,���`%Ű�l��+��|���_m�w�I��DӂO>�O�P���c<���T]�t��c�|Z����Jwc6���X������WI�@��2��}Y���q� ������hn<|�+r�:��@w��)������2(�ܜ��i�@�7ͯ=�(O��~�W�+kr�o��Ex-�q��7xU|u�C�����cP�:nm2"m�=���:��a CU�r�7���PF'���I�]��V1�5�fr��}���t\3���K���'�
Ir��/&E��TdMvnj.��np�	:5囂\����à2���!5�����Ȼ�6�Sv_wY]�2��9e��@�m����쮖�!�ϑZ�����â��+�vK�ż
�Z�J�[+��m����F��V�P,���5�����u��-��T���)�y?	�X�Þ,��2g}�J�Ò��h9�/T�硎q�h[��5���=ں�޲86�I��0Z�|齂2�q�L	�3t�؝�>�j�[�+W�Q��5 �E���f�)���w߁eF��Ea����M7��X4�ĉ�J/'�5�N!�R�R0���ƺ��575a���-uM����#��(K�Y/��Q~ɖ%�T�2��M�X�jk������&���RX�>�1�� ��|�V0��'���ZЁq�Z���0��
5C���� ��a�r2��������X���C3q,�'h�X�F�(1��8�7)���v���F+cj�W&�:����T��� �h�Uᥙ%����A��M�*����?��,��Z�ܳ!9s�y!��r[��wڭ]�b��R2B�4@�&V#�������<7}଩��Ϯ�\]u�/�/¹r��U�e�\f$
~�Iu�%�-�zm� ��np�t�b��\@mc�����J�K�8�5�/�ohO/>�Z;h�^7l��0C��j<��̀L�ʯ���t��J�z0vǬ���H��s�X����!\,[��$�p��t�������s�v
.-�=O��+��b�H)�]�
��9�G�'mӲ�sY|s�S͢]��d����9՝�v�6��	�fؾ��6� (����o�h�	�$���C:��mFͥ	��V�����no��[���&%G�l�7��>���xv�MKDi� ��<��� �t��&I�*a���U��g��A��w ��zŗP���CV�&���6ľ5�çL��4ωj�*	����%��(�R��)��;��P�r���M��9�r��y�!�Am%2����\��h� �A���a�����y���h��tJ^�׉&{�\N����{Y���ro\���R��l�)��l���2@��sg
F%Y�@k;��	�;j�{�ƒ��������/J��!��LeOmb̻���Pq��4QUtOY��O���`@��my"ys7q�p٘��/[W�c]�^p]&�3�G:�7ݦ��&k B�~����"�X�HX�_*=��޴��Gk�f��ˏ�j���L�^ ���l�\8/�V�_��K�%q��6�~7o�&�B� =�m�N푡j���Ң^u����M�.�T�����O���r�6w���>L��uo�u���Y^�i��@�O2@{	|��j�f\,_UN���|G��7�=��g/������z�Dr�?$��h����!�*8n�U�ó�ph�F���=q."��,.���hb!�g59Z�˰'��Ð{PA�b�I
	H�)\��s��#�a���MB�.��/��9��]
+�|������ĘR�V,,�ʧr~.9kx_�I9\�t���p�D�S�Z0��#��X'��l�e�5��C�<Dr�M�](FL��kc2t~ �U�}69���tk8��!�Nz�w�U�m,�w�=Fڰ�~�<�&˟��Z�SկY`c��9�����y����但W��q<I�E�Q��<e:�c'��๠��� �����_V�ʕgq;:(�9���pCH�i�|pO�������z�ɿ%=�x-Жh����T��&յ�5v��q
��������x���5,�����~�o�~�<.aՙXR�|W�u|�ޕe�h`� Q���Ⱥ �Ki.Ϥ�!ֳwƒ�R �|�_�e8���Iuc��{L�.��Xy�¬���*l!�W��bW²4�d��K����Q�)���bӲ�����z�?c*�>Lc��� ���XM�N���q0>/n�Q��<%�tW35_�Ido���������y��X6%0��sI�	ƥF�����ԟĦY�0�)��������,z���d���Ok�j�֜���wL_c��{��Ĺ�2m��::���2k�s��V�Օ �/��OM�����`y (�I*ߜAu��QA��;�i�!��B������Q?��s$��� ձ��B6����F�+np��Xވ�*�Se� �:��Җ�H�ou���amn	 g�c���kuIb��pST��#�f�ՙ��Gc��z""o؆r(�����#I9�5�m<�u5�HA�3X�+c{�{���x�rg�#��Y\�6|����-.hxϣ&wUO%��P��MeZ�gI���CE��#��3v���]��8V�X�3-�v���l����;`@��>�/,�'+�+ט��	(Ͽ*�L�I��5Qy��{а|T��U'
�-�@3�t �����(�7@$
2��K@�e��N�s{x�ރ�����t�x^�`y
�I����� ���5�v��[��W���I��bX�0L�&����������aF����x��O�eޏ��o���q�d'5֙Y�g�����	�ߤ�m� Hzo���ue٤�OMy���2��*xK9��j���_�(H�w�������2�d����M?]�A��ԓD8���R���S�`F]٬TB-}�U�I:>Ҷmk�T���a��}��΍
2�U*�w�-���j+�T��
A]�1qD� ��R\Mc���ȯ-K\�[X���%�˼�mxO��R��C���})�F�����
�d�L�ב�8�fj�4�]g���V���{�A�26`W�-k�h�C7����n��7ܿ+��Gt�cVk9wG��':N���Q}pNWT[�4k�U���ݠ���w�/jM�����h�Y�N$��W�!ю[V�s�z���7:!�1���~$������= q��qej��d��zs�.�x)S�[�_˵�/M�r���9J��'��LS���Y������7-�S@j��7��D)4��@�Es��NQRL��&V��(������G^��j�T~��g���>z�_�U^��Kb�*��Q����P��u�A"F}�;�����Y�R��G��0��]��s�w����Ȍ4z�N�-Y���%Z ��G�I����6E;X��56�Yy! �5����������H2	��ܩ��� ��5@�1R��H����9@azo��ڲ/�P�!VJ��آ��'S��7C�>]{@|U��]�2��ߕ��1�����	m�$��)�:���3�~������m��6X��I.�d��9hj*vz��]�_�Q
����ԏ�6"ӈ ����;���_�JΡ��H���۲Pꭠ�`��R�Ik�jW��X%���ޖv����`C,��o�>p��cz��E.b��
 �H(��G+�0x���p�M��L!:�ѷ�s�Zz�<�o�o�>�FY(�����0V������'\)�	���"#��9��:J�%H�g��QtUf$�&�\�V��5�"͕��y-��E�*��df��f�"tdcgW�J�.�\�7���K��n���I�'A%�P�vL��H	�`w�a13�.��g3XI1�����-�\#�Ӑ2i� �L�E�u4�&̙yG�ӽ��Ƕ�P��IA�*j��{G凌a0<�HQ�N$f���F�OqB�ɖ��v1���U�5&>�p�i��SřM?����8����8\���rƽ֥�yl��o�q�Q���y�����	(�Gj�z��%\AG�{���]z�)�o*���+0��>.W�%Ua M�p����y��2^�Na���
��b�����%c���?/s��SQ��>�׭//oHhAύgk��U���X=���n��o)z���S��*I���;d颿��MY�jj�sTj���	�ZX �E��<nu���w�]s�w�E/[dc�5	n��	"|�IX'Ӆ��?Y$m����I�bg�<e�w�<<�JRQİd;�n&F���hq-��)�s�D/�.��=��~/�Eg�ٽ�R��AB�}�xf>2Z���v��<�5��|st?S���T4��,Lvk.8���-����u�hι��BG��:�5��]kF�r���?����+T����\8Oz����!���w���>^tZ2� C'�d� ��b�c[!��Y�FB�����k��:;��B�1}q�;uA򃟦������0zJ1�1�|XP�#���+�4"�s�*�"*�gAg	��G�`3��?"�Iي3晉��ij~�3��J�N�7�(�I��dQ}�GqF b��������Q2�N�t5v��k����15�5O�)#h����������������d����/}�W��ŝm�WjO�!um�2�`y��V��S]ũx��H&�=

��Mo�ʿ J���y��؁�)�+q�͎�Y�X�Q0��I,���eW�=�N�����E�٥Kkx�~$J�V䲙4�����9oN���f�K�HJ$�o�ӽv�?`�rv�f�-'��|q�~����=�֭[�΋�+?޷�R���w�K��a>S!`��)�b�_Q���E�&'"���?ݫ}�i^�E��3ur���Vc��To:��OA��������5\�N3��)���$j�5��-1T���]�Y/�%��B��F�V��U�I(�.`ڳ.��-"�1ۈ��;~���K�8.}D�?��"�JQ��_7^�L�����}���'kCh��SM�g�!P�ҽ�O�$��E���� R�5s�W���4Ƒq����/Y��.M����*�@�޶�@�5V앢-m5?DrU�����?���0[Ʌ�hxf*��+.���ǋv&�[<<�K�A6k��b���{,����r]0��*$�&HT~g%dVMF�4�UP��j~�A�<A)R;�i�DV�8f��������Pч{W!}�yc�g�ˀw���Q�Һ���O�F����1���X6cWd���j��V0���A��߃�Q(�A�|J�U�$�3�[
]ğ��Gv�v�o�Ǥ%ü��+Z�d�Y^��|š���1-���������s�6i8?�Y��[e��Fө���o�;��i'�0�YM�0��f~3�B�olt<޼���%xlSaU�<003����c���!�愭�% IB�̡w��AF���/�M����/dFZo�J�
��C�� U\)�r^�N�o�Mӳ��l
�p{�ݛ��f�E���(?<�[�>�w7r�GWV�F(�+�R�ğ��#&1ˣ�00*��@.x�`a���y����<��:U��,s����2x��l7���r���I�1Ѓ�Z��;蛆b�2�A���@����%8��BU3��.,Ej�^�����tdx-��?�W��<�o��������JLX������9 P�=�"����{�<JB�e��K��-���"�X�>ޫ��K�]Ylh�JҀ���*f��{���
��:GSLVB�%f��\M�O�q���z)I��&�\8���f��r��M���_��  "�_���3��,�$�|K}	}�*	�y��;�&�>���8�2�[�pB�m����[�����M������o����wV�I�G5��6S�>�cȰIh?cw3�tA�e�S�s�{?t����`K������`��w#�n�ZMJ�4Z|����
級JC,��G�f)~�p��o����	T�^!}���o�̐���6F�+;�Ų�Y'9RbI����U�lE,�9��TRX:e��G��B5�<i����l��+� �<���=�����l�����ƣ�F2�WT�\#ewAE>V@>Bf��%�/���]�A<U�Jܩό���������N�:V�F\�ϼ#I_��'���!
��0b�����}�1��p����G��0�+<��VV�X��]��<l���b�"h�0?�'���	?v����vBP���LH���x+�OY4,"��FT�;��P��L!p<�gF^a�x\�8?ڥ&6j��lJ�vD4z,������~�Y]�#��Yn�EtA�	�2"4$����FA�eq	���	��f�m4�@[לE5O�'SJ5g�0���l30(�q�e���J�w�*�����g%-K7��5^Ý�Ӏ�*Z�I�'Y�^���^�`�	ς��;<DWy����_���HQ<a�l[�h�	!�R[��v:�U�?L��ӨI��k���̀��?���z�zG��щ��u�R�r�7
<#�t�SO�3\�N�7����N�}����A� u<^�o�TW��Ж�뷶���(�����4�������<��B�[Ӱ�{��/��2�u�{�Thek�HY��U��h��R�x��q�*}�"Q�|�A�'�y��4^ M'�8��6u��do,Z�lKY��"Ϡ>�4P4�
�AN�4������
�d�Mv��%$F̂��Μ�-�Eږ`���U ��,I���9ʈ���sq�B��N��C��݁V�41��G%���'i�=�h�#�cA�&�1LBnܫ:!]�<12M|��A�f�qG0*|�y��;1~A��8�^c����i�%##�0��؛���ݡ,r/�� +�h7>	4������b����ZUT��&���'`h�Wf6C���$v�r���ޯ��"��M�F�H�s+�@b�3g���5�2�g��n��\��n��$~���z�eV^����+�I7�[٫�i�jê��E]G���Rw͎���R�R�\k��,$կÝҳr�2�\�KN�s��>���h�yN�jE��ϋ�Q��e>�\��(4�I[5tυ��5 ����[��"
mb_��gJ��C"�i��$�,*�}T#�@�z���2=��`�\R��ҼC%qft�P��U����:Y�N}O�o醷íx-�4w�D����U蚻���Q	5Ł��I9��$����q���X��3�r��e��[G CP�iH���}�*i.1����,�=��V�]7�e�#���6�: UpG�6p�jȆ��������Btlݫ{��^~?��[���h���:�肶΅���]�"^e��h,?��x@��l���d��k��Ւ>�琶���@j����0��>� ��+W�;�n𥠈��[R�a� �4� q�p]w{:��5��+�+������y��~�~�zeA}���Y|!�J;��(�M��=3�&�ӱcG���e5���$8}E7���9�X�Nc\�HYк!H����ŗ�t��S�i������Sq��������E#rE�/�[A6>a��`��ҩ@c*�p���À<:�ƚY���%��]jˋ�6Ǘj����S��@�w��6F�l?��c�	�+dE��]u��E��-�m����TQ����zK�ke��hN\�΅Q����^b�Jb����m�#7a�H�4�Fj�F��'aK.1RE(E�'�i��$@̿�<�;,C�M=�����]Bs���{#���'fP�����
bt�%�%�?M�i�|�v���lFw�8�8�(��z莳K{�^�b�*��rn/�޲{��	���?�F_.�RɿR�����vt��(:�hz��f�Y$���)�W��]_��M��Bgӂ��$�zS�i��Q��#2������F�~� oᱍ��~W�!��b���{�]��q�s��,��
G���t>�)�.��呾���.�����q�/����ׯs��1�3"����x�0��,�� ����&{�6�x���@�Z6�P��k��?%ɵ���|�4l-i6k;�����k���سsn��+��SFǜ��ݮڇ{��%[��9�%;��ň�يxOl3
a�MW슖���y�K}6:x����|�s2"�^����b�_�m�/����h缪��|��/ꤦ��������)����&��i�L�,������VI:��u�v.��z���p���up��l�jJEѨH� �J>���ܤ@���>�V��L�ဟ|[�z��f��Bc���Z\� �f�$�Z#� ۀY��Xti�2wȼ�Hw��ì4�ɡ[L{Tm�?��,�jtsC���������L����<��q���US�v�f�`��M��S	tYW���U:��N��{�|{�M���a���+dm�k��Ζ���)�,E6����k��FQ=(jO��Ǉ���\��xM.��[��r���k��K�����eF��A�f,�{��&u�TY^N�J���dy.it8M��Am��OoF������>jB~'�bHy�O��^�|�(dA8yK;ng��{53��\���`���$�
M�!I��_�~mre�Y�~�I��2��^�a�7��y���R�r��j]̛Ђ��x�����MI���BM��~jE��#�:R���jgav����"����~:`�wpa�2ܮ�Jp��1���,yp!��#���������M������+p��݅b�X��y&�9.6|�#�
s���
�H���ˁz�})����6�e@��$���m"�n��T�V:�v������_��WT7)���r@Zm�nZN��o�j`��4�[�&�(�l�}T������ZD1�c�ќ����n�,+���������+y�cj!�6�V�\�j��oS�/34�aK*�M���h����s{mCz	���b�n1�g��M���@�����s�"n�SM��U�I�h���{�J���i3����Ys��,bE3���: �}�*M��~۠MM�Wm77��/4s�W��~�x|�;���N���1�\�k_&HK�� A�>��I��׆�/���O�b��'|tr�9�7��y����E<��#4�6T�,���������c�K�����)�)�Ո�V�s�6U" �
5%H�;��Z����u�����eǈF�J�}BpxQJ��	�%:f����蓒2�Z����y�_*���g���[o���4*mz�=�鯛�]��X^*bo��V�El��f�MU���b�u�t�s�
���͟��X�� ��X&�yrU�(�pǾ��DШbFz�)�m��Cm
��Slt�n��4����D~�7��m+ n�&��g�m�:Pu4�d�����٤m�,�q����q��ބC��F���U��򛼳올'��e�<��&`����ciRN�-��`��o�����Cݤ�k�/]a�D=��"���J�Z�׮pg�]ç���yQ�N��g��TR�� �8�J�p��_�B��q$7�V�l7��������3H2�qv�nI��t��߂Ǒ8/ǁ���;��/�L����8
Yi���� �S
�)�v�up�Mcwj�T�X��t���%����>Y9o �3�3O�}�r�+�o�s���tcЍ1Z���BԖ��t�B�v6gЭu}N�0BEr/�Hc�<&+����lY(��+N�7���H�M������SPmoL�}�a��)���G�k�u/j62�o[�����6f!�p�v���T� �z*w��D��Z���L��SޟO�
�GC��W�<��kBg�jf���⇹/Lե�����i�<�*ui=
t���^2�b" ��j���=���"�=��-(�*���|X�cf�g��sT�����R�OQ0:%n
q�V�ժ;���:X7�"Hi�o��@Q��\ٹ�z�;j.�I,�ZF��Ov\��k��1'2{M1�Ȏx��?D�ڏ<��� =g�-��
O����(�Y�;�g�ݲ�����'�.��uY�`~�\��3ҡ,?��࿩]1�����$m���	zm7#�mu��kf��ᄮ��Vik�j��0R2l2���ޤ��A�~�Sq�߹rM��J�|,vWX��s�[�#�<�1���8���b�U5���C)a���.
;a�rjh��(�����"� _Q)�P]���Ӽ�(1��+3~>��g/������^�W�Ҕ����X��hz�a�2� ��:$�-w��DZ�y
��G��\G��S��5���l!LT��`F�%6���|=�x��}�xM�� ��8fL��s{�_A6[E2]q�JH��%�Ӹ��ӵ�s�W���١������o𱶈�崑�`�C��\.M��o�fX`����B���M�Ҵ��&)�E>"ܙAc<���^���	��z����/�f,��ME@�����-9Cn�3|�oiI�����Ӷ'�|��w��j�,C�zμP�Y�͍`}&�z��]Ύ��8��d��n�ơ����e�w��.#�b��=@��pbj"��D�Y��u�ٺ��n��zsܖ� {ku7x|A�J��d,��0��	��}j���C�gȜ'f����{ܻ	��F�����QX8ӏ,DBiB�CNI���(1E���?���5�nE�$��DG��{�P~U�u#����<g�v��;=���2z��jZ/}	���8�j*L�w�9���q����*6�әԱ���d�8e��Q�P�Ԇ�@��ܐ;�*jfV̽D�{3�s��z��P�����_����&o��*�Ez�����A17�7b��6p�1��Up�����M������y��r�����}�?�>��R�,�������QgC52���NY�R��e�V�!�ݠm�$��
�~�6YY� ��|�-ì�-A���U�-��_���7M� �ؼ8����7���C^R=Ny$�k�YO�i�
��G������iB�z�Mj���Ĥ�t#on��I?�*�;�1�)��z���c�T�s�`�t��32$ �l.����CV����[��vcmZȆ�Qgv����"/N��O:�.�����FR`$֋St~ʣ7G񁽃Fa�1Gs�4F�L�Y}"t�+	�N?U@a]]1;�?{k���!�b���˨���-�,��Ŵ$�mP���]�PX�9U�<,�1��mL�B;��<qE��k��j�����j-��U�w�jBUZ{���p��WC��\~SM�]�O.d�^`�"�qV�kk���f�Hq��!��g�JTi��+g�w�f��txR��SWl��GV)e^V�\{���.Vԓ�O��
DM��^��C{���ːY��w��alX3�	G��-.<;��)���&�E�#���)��\Ȳ���d�Y׍ �R�U�13�+]bCx�&c 3hJ��H7w4�;�Z�@~GgQ� ��AG��:�W���'���ޅ���P�R�'����/V�lfލ���cf�=���P�-�K�>�@����;���_C3����!����F�g��F������p1{+��Ȗ�K�f��B��<DJ*Jk:��|��`������������IK�LP��.BCHPW�;�<��n����r�����Z1�EOR"�ȹ��xl� k��τN�Z�������e �"7M>�����A��;�[o���0�R�S��C�`W�$g��^D<~&bB�A�F)˟�������������2Ce$�� *&_�iZ��ϸ�ҋ6	��h�Rg�@n���>="���XU�V/����9;�*od�#�WCUx���t�� :Se8HD��V��ꁠ��5`4%2� �*��+�_�	�z�?��8��UY֊Qe*Ȁ)��Z���a�U6��o]�	`׃XP��u��E�)��EX�ʈ�C�)*f�`��0/��q>�5%w�F��݃����Zn�v�<����77U��6����b�)�������ġ]��(nQS�E-�A�zy�9}gN��mM�7%�Ĥ&��¤��_�9��cc��<FP��h�u�&�U��Zi�r?�J@��k�s'&ֲ�{�r�J)ݐ��w�_��<�R���{��Q�u��R�Ꟙn+Ȱ���Y�33���K�&�gD3g yH�r���L�v��N��&h0c�X��7@3��3@;h��������R,�����d7{>�jm ����:��MnXƳ>[C����y���7mo���	����Y򴧽=ڡ��5�������Y+���ӾҲ$�u���^3����'�jG�� �l��P@ȯuB�LuvLk��s��U��5Lk����'�\r�;u�x�തh��<g.�����q����BeF�0��4���=(��B�/�D�cc��z:\�kp�:/a�
���9ğ�d�Vo6l���|�1�2�uI/��4�W���`GAw�Qyk3�))���C�xA'
4��>&����B�{��K�B��x�����÷������V�ҍ��B��Mg����wBB�jG�'����[R��X� 9�S-qt���% `�1c�ߚ���Z[C��[=��i%�17�:9���I�vl��a��� �$)�1.'g��)%�K�<�5Q��d`W������4QJ|���g˟66:j=�	�v�z�#��i�;���������{�4��ӝNV���^ "�.��Pu�䖇�8�U�R31eB7��>�����82jgnT@�x૞�cWz�V1�9����:��?���R��Y7�|���8J��K���n����_AN�,>�.�p[�G*�7��E���:5`�sџЅ�^�ܞ��)�*���׏տ|�Hm܊"Ŭ�j?*k��1w��G���z���:�?q'>Zn�w.�o������`���w����r��Tr��{�g������EYl�[�	�v��e���d����9���u��a�WV	�� ��4�^^�@��5vɟ�	qT�37_��k�7��@g�$ϰ�n</k�I��X���]���`5���b�0�X>�}����zs}��̵
��1��}m��\��V��д�;���̂���x��
�?���2j���ov���J�@����b�Nm%�o��U恩�H�MI��O�쬒��z�o'9]���v˝����x��=D�Z�����Ǐ��w�_�R��,��^����g��zk��~Q%Z�m�~Y���j��d֏Y((��9��k�6��M�>:��	������FZE{i0��}n���a�?8��MZ(s�d���yǂe�o��M\�%6�rx���V���z�7P"�@8��S,��a?�jer �:�+�Q,�lR���:&���Q�Xѧ?�6� �e��<p�Z��-�!�~�v�����ƞ�afdߴW��5�e�	c|I�O��z�� rdiD�}��6��Ty�N0'������"Omյ�(�۵���/"��G�G�����IN�Z��lX!�D[H�/���PcOo{��+|��lۛ������b�!���ތ23(��;�~���mx���r�Αt�>�e<}�yU��O�g���.�g��sF/��rSy#5�9�;6-O>�Q0�9D�>���õ�a��� �E;����^�c��9_y�l0��Qqދ樫�.�h��Q1(�n������E�i/�G��A�i�ⵢxN�?1��n	G��7��P@���һi������ԋ ����*լ���+�H�ئVP��<��'������%O�;6W��bF�.ڝ5w�Vx�Lo���By���{�5�Td�����������!w�#?H+���Z�"G�5#+�|(�B����=�0�BYM�p�q��w�t� &E�Zw�+di���jE���������0Z-�Q��jL�fL�����ʷ�ڮi���K� �a��\�#�<Ǣ<�'����Ɲ�$�^�o�#�!��G��qK���S��b�iN��	�ӕ��FXuoN��J_�~S�B.�}Ϻǣ�J#��.�3|&K�W/+=��KK�	��z�;� ka�l�Q�J�k=�+��S�#W!y�г%4E#/��j���fWA+���~ZP�'0��f����`����fH���ľ<z��'�1�y�V�-��JV�{=d97��*� ā���?&�)ѝ&�Xr��6���	�^N��H��L�f��>��f����(�e��`zE��J��~�V���Q���ܛ�?q�qsI��0�J:����k��[crCj��>߁}D�ZZ�Ԃ#^�m����C��ƣ�퍅?�:�j���M��IQ����#�Or�ȧу��;3��5Z�쀚T8���,]� ��f|���t���0F���)T�<E�:�T�!:���@vKKY����������<�`/P�G���c5c��8E+b�h�X#~^�e�s���B]3���/�&=xdyzO@
�����@�yH{�E)��M��ܰs�@z�0�^G7�O�@��gqgi���_:K�5�::��� �{�����=T�N�7����\g��#O�в��D(z󗓠�NW�fBt�6uLc�R8�65������:[�Ȼ�	��Hq��|F{d�x_Z ]%�� /ÞH/�v%��c�c��M	<N����U�,?Y�{y�Jĵ�/T�`͉��Z�����d�A��|�fFNً�Ʃ[{e�08��UA�΂z�k����S�&Q@PwYC��64-_����o�+"C6���5q�S��ٔ�������V�>�;D�9[�V�c,2]m�m
���q�97O���dwj�d�:`y��騕!46�3�u��j�Ơ,I�e�����w��J���,��\(O��J����u���r�b!��
�>dD3 ����֨�CH�OVa���|<���E�m%c+r0��c��U-P��c<��������'a���"�*����O�g! �@U�p��	�P�������T�O�̼���Fo�q�*��_8|��Ñ�"#���L����7A��W�+�������D(혓{��3#olv���qH�<��n�N�l
�&p��X��8�u&���g��!���v�Կ �弣q���� �}���i�yC6K�Q�T_T���k2h�"�G��w������"4=�c�n�@�܂�|��=j�'��3�Y�a}ڧ�&���v�`��H�(�������g=/���Խ�k���6� A>=,�Zɬ�]���޸P���"�f `�ޔ!LD���Ȣ'z�,pt��k�)n�z�"��p2�. B'��T7zT,� ��;�H�Q��Q�_����D���̄�S���^@�����f��LO�ג0V0MI�7C �{
]��9��К8J|j�n��DX���/���"��>�~v�,Y��9#�#�#f/|[?�t/�U�,�>Ub<+����2��>M�갟�!��;����Gnw�P�/�ϴi�����'5�lM�>�J?q��D�ļ�$��,���u�N��p0�kdD�Z��uO%�ƍm�cn��@j�C� �(O��a1P=���.��H}0�mhԤ���&{����D�a7z��Z��F�bNтfZ�q-0.(����S-�ry8�B�X�s{A����S��\__"/�L��Q���<@��Խͥ�~�A�3G6F��"? t�d
�p���'���.��e�`����HX2�ޔ��s��"�͞頛�\�^Z.6�C�������'<ڣ�gfAx2Ӭ��x�叨�r�9��kʨ%]�����8E��<�?��;��H�B�Q3��� �]�8���
�~�}5\U7���ϑw�錿�(4�	�m�4-��>�%&�gn >f��`p�}<�
��Bh�	*s�w/�u���f����m��[���Zwx�,8���Cx:��܆��0�6�*���X��f�Bp�!>�s�V��Wn�?��Y|}[dTY�%2P�%�Y�藯x!��9� ȳ�X6���҇����Jd_�c�e�}%rR yI 6o���G��;l��Y￷?I`���j�Q1}\��t6���<���R=X^�Nˏ�ГKjYQ_?b��D]��}��uy�6���=P���� 1��o>���뢘�{�/j�2�� ��f��
� dʿ����S]��9B��.�O�?Ӕ�D��ף�NC��(=(�0Z���]�Z�?C>U�i������h}ɷ�'�rl���qO}�`�4��|=nyee~�@��}r
U
̮�v [��>�p'����D܅qs��FN�ex����3�l׾�=*�b�z�>[Tԉqb�Ƈ���������֎�Rc���t�k�kBN��p�_�^���PX�8�P��G�.�M��.vt��|�qva���j/��F�=����ĵf�6�������u��u9�f��4�ks�����ֽޭi����3�&�y,�/�~�e����
�Ǎ)��v��}S�������l�H���l*�b_d�n����/G:�K&Ϧ��?u,������7��ǿa�)��~�	ѐ�� 6x�i!�I��3�vpC]B��["��(����:�G�f�'��������Qs_�3I�e�X����	ԕ`Md�~�t���;M/�Fщ3��V6.#�՝6��?�znv���E�7a���3c������4#�����!\���X�ٌ�%Ͽ13�n~?��<�a�va�a�m
�Z�W��`Ж?�Wۓئ;�퐨��䖲a�7������9�=���MϡN�J�q��xQ�޻gς�����棒-��H�g>�o^i�ݓ��Qr۾�	[���$�v^��TiV��c_�/��!�cihF	��8�FB)�r��� r�J�� v-P�jf�"�߼��X���d=W��\����U��W���A��[: U%I��/i}-qߛ�}>��p��l��l!9�+�d�R�R��<��!�X4�R��E��y�J� _�q9����PŰ�g��5���SN�1my�q�3/&���Dh���/��҉$���i�',�*�U�E�����[�t�91��6�qd/�&w�v{���I�A�H�<�Il�]�t��3�Z�,ڟ��ܓ��`���}�ub?�W�pr����b��Y��i�	Uey��S ~ �Ϭiz��,o�R�QA�չG4퍔���ofX�}�b�Οy�X�<;��q�Bw1�A󵶗���|~���}@� �Z9���b�T�Q|����g.ź��0b�Gt�#irr�g�p�q�8�]��I�ǥ�iǺ@B��?<��_���
d!R71TW����{��(L�vO"%~�|5��5�GL����EV��9��&�:^�ʌo##wn�����s1�=�v�|�D��i��u _���T��.��dQ�)C����׷{�U�}��C��i����H[~5 �&�>��&e�#�R��V�I������韘uڶd ���ds��7v�S�Vr��*�w��	���ر�[����y��80��gA�d�.���$�|}�Yc�I�hf�����P�n<ɷ
f 9iV��S�b|�4��3��,s�b�k��6������v$��'�5��g�b�� �F#�D#���'_����6օ����~*�l�O��p^��$���7Ȉ�BiX���H�J!"�GV%S��|����۪���Q7;z�rP�L�V/^<��QYmqK����aΞ�3A	g#�r�LE��s4���y���$�BX�L��T�r���`&m��+���A)���fG�b���"o(���뎿o[(� �{�	v�FSL0&g<sa�8C�\O���R����۶�e}�	ȹ��Ey���|kᯃ���Z�+�?����.juH��&x�|���O'ђgc����yT!α��d��CO�3����Ab�����je�|�X�a��x㔨�R�M�'�A����C[ji��P=��j3�u��]�#�����p��Xƶ2AkL���q��Qthx�W��SA=�4-߁���1^ư�K��u�3�)˳�X�<c�7���j�k<lİ��p=n�Hnf��j��w`I��q�@!��~���1G�FW���!a����f�>�3�Ī�~��������q���\�Lt���hȽ�xH`	y�s&o@ >�`���s�)�k��<1�"p���i%�sw��N���e��i��Ǻ]��E ������7۠#�o���ꅒ��80��x�[	hN�6�rN��N!	��@�i[��e�ZR������[�\M�͈&��+��H���֧3t�&^JkŚ��Miݦ�l������0�2��ΓvE �n U]5�q�R8�0�֡u�i�Hc@����K�V�8�H��n���o>�	��/}��"@]۰���h=�'�*d�rW�g������]/�}~������6LPnV��87s���L*$��Qm��G���b���,���_�z��j���Sk����Uh��kg���xM`PV�̃���<]м��~�<1VJ	�s��5�O�p�󭄣�7���ɰa�g��*3��XsL�澁�zI���8hZ�@���7tn*
P�K�ƭ�h�aږҔσ�֥��N�x���V��q�Z�2������28��X�9���i���N	M���<ل����4n��YP'�~���" ��,/��W�֠��yR��0��ǔ_������ա4N�d��#�t�mj	�_�������v2�M.�Xs� ��	l;}�aZ$�of鳟�R�J ?��j�/�2g�� {��G���{Oy��>d�_l��s�Tܳ�&�֦��8<}�##	�KO�f��o �����
l��4f6��䈇?Ն������˟<�k�y�"	w�YC��l;���U`t�d��՟�;�׷��X�,X���4VD��\F��9�=����wc�X�)X���r}<J��+iI2��z7�˂+D�N)"����C^'^
�fd��#C�Y�J�,��-�^Ø��>�1�#��3jI^g�ʗ��~��g�V�A�@��j�?�o���rj��),�|A�`�\�Bv�����Fh�]÷���C����Tq4tc٥�*#/�.o���PKxO�-p�0��m7����2�{����ذ�|v��-S���6�L/?��U�Z��䃳�A���+}K��,c�w�k���5t�dT?I�^��X�j\Gs�T��������6�ǝSQ8-L4������TA&��Z�<�[��&�NW'V�,��%��bڂ��
�0�_ҹw�!t�6����e5�@ˠ�6�l6��M��"��4��&l�I~�w��C��ݼ�-P���kLwB�E�̭�k��e��-3Q��O��º�b�\2�0�Ƕ��?�)m�����x1��H��G wO���6��ūS��X{��(w�񧷥�v�/�O3=U=�*��E�!Cu�\XB�DL��;��=����;Z�$0~���0d1���߅U��@�[���N�Q�D�
�ףq�3�E���}>�bJ1��a���#��7�:�[�b�dc̰53.�{c�.�h��8:H�)ǵ�g��%TYz�>v�&��+%�q?����Y&A5�~�_ơ>��"NZXώ���Z�*<��46e�D�]�x4�e����j��OU���D�F�Ӛ���S����og{�qK�0�.Rg��SǴ���KY���]����a�\��CB���0-X�H��3�AؖTL�����	:?��Cn)�<a�w���;%���ħ�aḔ^"]h@�c��c?�_	h��M��~�'%�W���ᴁ!}���8�Eu�苑Q�?��B��r�c��j�� KV��_�9kO�D��):�W~��=@��c�]���C��:)��"#C�V�6��l}��������x��ޯ'�IM��4��p��(�4e��5��a���R�6�N��N�����T�6I����X��[K�F!s��������hy7��s�L���c.��R�fM��^�G4Okj�P�v�H�i��{N}ѻ�����aHv�����⸳� ���.0ڸ7<����ȑ��5>f�`D/�L
L��9xu	�,j���SRBQD6{f���e�?�q*>��<4��p�;8�4��2AR.֓���`)���"����O���n̷ ���G��v���˨�������m�݅p�{��o#@�Y��X���H�H�;;�h)7aىl�3W������|��1�~c�Q`�����ם&�|�f��ў�����b�V�UO�8k}�Pߓ�/d\��qrz�_�%�cd�0�s�z��J��j��j��B�>|e����Ƀ��NG%@�x�c�.�]�cs��]�/�b�Kz�����$�r�F5�:��k�]��lq�t�+aR��w��*�_�s-R�6ඏi����CPw�]8mu�P�������_�-�l��-3���^������
Z&�Sn\����mv��bH�5U���Z��r7������������2+:�Z���X�s��?!�{;!�a���Zkz��fɽ�j�G�Y�)oF�-V�V	���t���z��-��  ݈h?]��V�3��tVy�%F�-�L�`I��'�����x;?������D�T�&����&� >�$�zq��{��Ƣ���E���-����[���'�σ���)��&�pgN]W���BdS2�v��_sjp�r���jbӳb�Y��)y!f�����H,|��d.��Й�r+�3�6܅l����٪j���k.9P�[�}��o��R��o�[��t���̤�K���Z]%F �hX,��'5�qW��}�U������Q�!r��`�	}�G8���'�F2�N��- ?`Z9�O�\�J	>��.DK���ɰl�qgk�kd6>�F� ��@d]O�?���B�WFƓ�<2�}�q�rݵg����	i�\�-���Чܲ�b
��@AN�g��c@���Y!Q~����KŐv#!�_�B?5�~�ƩNʛw}fw�쐦�ڡ �#Ѕߓ��
;}f�g#2�$�Y{�j>�ì4������7�����}�]G�̼���Sr�ە;���b\3F��8�M5&����|P�]�k��L57�o�G�x�&��%&|�k�ЮD����̬Kn|����$��p��඼�8.���%��N�c_�9x���ٜ��V_J�����kv���˭q�����B�E_ZI���C'i�Ǧ�@H�?*�F�0��(��"��N��
Ό���q�����lV�j�֍7��;��#������4`X�6��T%��.?bk���z�r*�-��<�|)���	�#-��HQ�(���e���К��j�9:���j�B��"V0�����������[�5�ˠ>}����K����UY���-^c�q�St�t���?
4b�dI���8��!�ٱ��"�]��Q��z\LXuiC���V(u�*%Lʴ"}���;�X)�5йw�ey����?F5�����!�	{�/���ͻi��M��s(��H�+�����	G�O��3Ϩ����Z�S*˚+�	��L@'_5����rC'��$��zf��c����.�3$y�����0�zM \J��p�����a��m���>w�&Jrp"$"6+�Uw�;Ϛ&T*�:���?S�oNf�5���s���Kv,7.u�u3��V�w�NOk�_��H?Y^����|�>�*vv�jԏ�6��K����yA��F����N�Y
j�VcLtV�Z��]���s�>Z(#����g�K�)�T��GFk:]�%�w���6���L�ט�'R�T ä����up�V�q/۷�}�p�8�d �<�%�g^���~��n�$�"��jm.�$$XE�r���{<���r��D�>+^�7�/~4��^�ztl[1L�����;9��D¡GOLe^k�a՞���h�)�E]��L�s�uK�Hk�O���_�%a�餏B�/.������N'�d��ϝ�VӐ���W���C~Ѓ]W&�E�ψ��0�Q����h���o&�w}�l�{3nmk[��"�p}�:j�=|�{q{�@�!�!��kY��F���v�����5�G=�wrJF�zm�@���ɾ�&:����Ȓ�ÀLɐ;��w�IHk�C��p�U+O�rJ�Uh��]���BL"���L�Y&Z;c�!':iO�S��C[h���n�i��,�[�#��Y�~e�Ԧ�'R�wԾ<�VK��v�� ��G���ɫ2�O��a���1�o��^A���E�JÜ�ψ�� Z�֢�U����	ξ��U�q�i��<dD����x��f��.}�P�˖k���}q�E(v�z�X�[�<�#n�Z��zÌ��U ՕMm��J��5��]^��y���<+�/�����0�,�� >��m.�tp����B1������#�q&�t?��Y
��s?��cl�)w2��}o�Ϯ�j����:�i��|�)�G�.��Q�ku9�?B0�s��<�iL���\�.��A�F�R}7�v��OB���R������!^GsAMO�L��s�֨I�t���P�}ޔ4U�[)w���n�&�n`8�/����EZ#�iAȬq���pӆ�����ġ<�i�*tؾr���?���s.=S+���L���-�kc�d���R�J���6�%�S����|�n�]�7u�MǺZS�y�'2�ߏ�����s����م15ftYW��3��h��:aL65"�ɨv�7rq�J�����jTVw�o`B:�ũ��֝�"�y���E��J�:�p��&�c��8���]��&T����/R����������[,��|zs���(u��o�4� z�?����!�>�Z��<�]���v����d��#��8�a�-v��0���<y���C�B+�q��,}V�
�|��"�wi�þ�3�4gȬ���������s�k�ɩ��V�}���n.1���������||�&(&cK�'y ��s���Ŧ?����1�3e�
 �NS���|���q1��(M�������tޢ�BPĝYÛE��3�/�h?]r9��0�P��vz9-�#�
p$8n	��e��)��>�R�5��e>(RO����-�1pqe&Y�im��4ԥ��Sx�rT�J���o�wf~zP�cD<"�5����`�	����R��.�0ފ-D>	�˸*�5O���%m�,F��)�/�O.�&m�b]I�31ڕ�����p1�`�kmMվ1��x���C�`�Ӧ?�P��K�+��P�na!|P>��fq�XKP�C��:�m8o#<Mt�;�$4�J_��u �C(��l�ꂵ���0f���m"b�z<�h�Pһ����*��c�Dn����VT�y������5����q�l{�-:x�3�p����A��	z�7eQ�^��C�BZ��k<����5;�R��:��v'�*���������Bc�H���LQ/�{?�� "+���[*�q��D\
<3�_a��D7��e���X�%��L�?u���5��V�Є���N�Di���}��q����\=c��B*�{���.m`�P���&���BkFY�V
�t>�J:*������[�7�pW�/!�#����m��Sg���V��jlBU��#0�74�<���J�����.m���#bR��P����f��$��aOZGRˇux&T��d_o��2��?9���n��Z@�mKM�PX��~˿��:���xn/�S�O�% �*1k�;3\����P-��k�������欓�)�s�V�;\�n�%/:d���U��U.Ǖ+μ��b>�v`��ׁc�u�٧�5O��Q:�}7�&/F���W������O*�/�;�������7U�9��*5:��:�6�2t���L ���AW�9���*���yNI�{��8�P� G�l	�FZL�k0\�9o-���D�'S�L=�]Np��x��d��,�4ۺ�5"��?���B9���N����|����F�%���8�yy�r�X^�Kp�uOt?�:������~�YUa|r�Q��(=����[�3���#Z�m�}Gk��,�>�$��'�ʎTD�g98��N���u7h��ۇЕ�@��Ȩ:�:C�ӆe�A��B�ƶ���kv��@��������d�<�l��G%
�C�܉�hZv6�XٞH�%{����ѝ�؟�a 1�.]rM�d'"��,����z�Bb��gbX�_�EM,�S֓�f�4j��w E�AFH��#�z�H�t�V�����j���YCZ�TkŔ(>ݤ�|/8d����}��S�����_�V}L0���EíT��	��w��r{ۨzl�Jre,/�T..d��_4�ZN���_�'�~
nc\'3ϡyv\ϊ>��롐pG��fő>H�M���3N�t��f�7�|#�~�F&��@�k�@,����AF��X�̷;���ޙn���В�k���R�h�Vԕ�E����E q���"��å����rg:Y�d�R�[G�L=��[�+4F��0齴��繉�B
H�Hc" ʡ��̰�.I}��\%�  �=���1�$к��ei����X=镯�eOoa�C������vP�y�<z2VϬ[$�Y�6tXښ�-��ZL 1���CÙɒc�:�j�{4.����$�l�3Y^��L�����PT�F��(�������H���q{>����=rVW�V���En�o�|�v����*VM{ަB������Jɞ[�4i*JS?�SN�J��A*X �6Y��*�j�qq>���"�1x��m ����z;�!ϒ���a{��_���h�S���4*��iwp���;n�4��Ԇ�����H��ׇ��(���10�Qc٦�8#:�}S����_/j��m�����w���Û��k4Pϐ����6H��y���3=�y)^����u��r"5|4kDF��&�g�<E2 �I{��ϟy*~b��],�M����5]�֊p:T�'�4a(&��*�6"��A��r>JD�oC>5�Tj��=��#C��婰2.ލ��}L�Z��m����Uo<I���$�������Y���j>�^��#?��DT������{�mj�M���|oD�5�f&¶x��0��X��í7��d��L�<�-��-�O���~"\�k]"F�w��yX�8�G7���"��r�-�P���U��d���r�p�)p����)Ss�=�9��^�/i>�(�ƚ��<��'�;=�A3�7\�*ǯ/�T��䅻��x&o��r��"�-iWg�82.�1��0hU+�y���f�3P>�Z`X0��)"�>�S�˱��Bcp�^F���W�ǴiD�����i>o���d����5/�"�ul7zj����ViYQ"��ey���!2�	>zU#��-�%c� �,�% q��~1C���VlR�"rF�-KO�S�d�
��v�B`��������bGQTꉶZ���������4"���׸����`'^HT��	ԗP��-|��--�ew�A� ��־�.Y�'�#�$W�$��-�eKNs�4�GPGL��[jq��/�Rx�:Uf��?�@�6OK<�������}��B�����Flc�0�EK�KJ!r����N�lg&%�2���˔IH�����%���3�Z1k_��d������ѥ#!K���}�r`�>M�V�M��/)���S�0|��u���{�؍�ބ�gbH��U��)g����{;)3d��L�Y�FT�E��u
��ȄT�q��u�y%� |�|7S���'�T��L9M?6��6���ԓ�:�t _2nc�J�}�S�n{�֫1���8���0v�O8�ɣ`��lwuT�u�LolH��%Uh�Z<�T!�ck,��\�?i��x�%��߭1S.���H���U��DV�:�{���j�~�@��Zh�,���!E%��y�}�9�}����";���	ޠt���~�[��m��
zL��8t �	n�X����6���9n�W��_�p�g���&uSK�	�I���-o�-�S�U'�*�����UI���9$s{�rz䁐�m1�B���4�Dú~�]����&�+6�,t��`	��,,��2-���4�zjɘP��\*89�r^G�[P(j]оj�_�)�'1� ����	���T]�d1o�Nn@!Xby7��u��ku�H"��`%���a6�b��-%�R
m��3Pq����h�=����9l�C�n�<ɑyŜ��o����"U�e����X���Cٍ���k)�JB�}0��iX	�����đ���!�4Oi0��[߇��
	2���A ^ ���gsp�9� y���B��Q֫�5ۯ�]t+��IS��*NJJ^�VAf�� YS�	��б�W2I8r�Tg���$\���r����h$�SZOx�'��sC�'ѯ�;<�rX��V�@J�]������5��q>&�|��*�
���T��"&|��2��k�_~i�k-t|Ղ��;�n>4y`��]T'��Ӏ^������Ќ��`=*��5K˅��
�W�^�jMSI�0x�������0�9�x>5
>[]K��9�3��Q�Ӂ��X8�f���i}�^m油!Kk���s)��E�(�������]��Q�Ԇ�yf���
#�����!�Ϩ�2��b�,��sp��z���x�;3�Q9�ΊOޤ:x��6�h��مpi��1�T��h�a.B��Z��ioVp��}f�d!a��s^~5q�!�c���+�26χw�a]s��`4�����7����J�"��h�y5�M��,&���Lx�Wť��n�<
��&�Z�;aXb%�E�6`���~d"�w�7BUS�����<K�
�gwj{IR9�:q����eUs�4]�А����bp_��\(}�@X�o�2=��^�m��!�E�j`uW+)�?�JX��#��}�e�	���Nl&Ca���@: x�jw�F�q�	�z��f�!�Nu�l��sJJ��w�l2�|�.M�*'����*�q�R����
�T�;z�~�K���MJ�?q<	ﺢ�0���z�|�y%u�b��w`�ݢ��aGkN$B8K륨T�n�UF��?>/xY� מּJ
��/Ȫ�(���Z��sd��9d�0
��G������JJj��O��Rft��ȥ��w?aY��0v��~Z)N�o��$��k%O�|�
��8�6M\�c��?#��1�������o%��EҜ_� 	����+_��"�;Q2GS/�
?Ij��-K���wjLP�6Xf��|t �]|&��J�}���߮�]O���%�F"��(�r�~��*����±.�q���ۻª��(�"�Xђ��+�'n�l	<����T����5v�q@�K�lg/��3��)+�6D<�},6�7Ux4i���TjQ�����c���4�qE��6,��m�b,��r3����Y�'v��	������V��46^�龇2��)�͓3�ya�ǀavs�m�a���F*�`Bf�6K�Д+C99�EP�,B�&�j�R�#K�x ��|FAHt;�q
1�]�>(��5EL6?���7�tQ�x �[������X_���S��	1���L�(*u�W�#�ߜۿ�}�� ���g�0�9��<f��jRj+��6"m�v�M��Ȍ�J�?jg~�vd�������Eq3/P�.�<1��1I������{2-r��n�l�R�� ٭�P�-�Y����3��79�5�}Vh��U�nk	��=�8�Jy���y�^6�v��/ļw����?��i�h!ւ��#�H���	�Z����-A�<�gQ�V�!�����}�%�8��<���ɔqy:dbg����B�n��+�ړ{4��<�j��z�Җ������(31Gh�����[�?�al1}��&���P5�$Ā.)����;HL�>�E{_�~�^j��}f��e(�� g�|�aՄ(���a�G����9�Ќ{�u�y�<
�s�5���Kʯ��l8��YW�m$
i�\�B���S�����0b+-nF�U��k� s�H��Ɏ󴴗,7��� ���n�\��x� G�����U-��)t��V�o��չT��O��2��mæ!�: 1pl؍�tZ���x���G���9�#-���ΐ>���o�y��{7��7X�OTF�AidFxJk{�t�?�0�S�a9�D�������(�
�*Y�'FK?�{�7�?��Qئ�%�xb�M�զkG�b����*5\�n�Q~{'l~��w�K7'�P�đdŅl@�՚<�wM85K7�8c�c+�"�A���L�G�|�I6g��.�,A�f9�Lߵ����A�w;aaB��8A���E�ɩ;,�=��/�E`���7p\1�0�fN�������~Y)��Q{�8�����9����r"%��Q�����/�X�w1K_#2��S�����E�*��.��0SC�՞�Z����8��'(9��n��[,��������0rb�.I+D�\��ɣ�k���K��mE�8�^8�_x���-���8,y��Q+JƜ�g�/�N���z�X��d���>��!��k @�,)�"�&�[�+��x��zsXG�9��f�t��cw1���x�T�VǏ��X%~��T��C(1�:���@d>܇%�!��M"�D�����*�p8���_jF�w�#�$��""1�>��-P�B�������W#;�VbB}f�L7v���@C
};6~U���t�Y�JT$ÿ��:	�}-_X��F�j�&��Z0}b���A����>d��[��������!2��a  l.	�:!�,�Jߛ�|@��c��)_�r�?��9׽'|��ɮ/�2�׵�#y��&���i�^�o[�]6V(t�	�qȑ����G���>;0犢��-a�W���9F��p�Ô�a�������J:P׋݃�o���sy���~@����'k�)\,�G���l��282��UB�η~ �I< �K���C# ��}�E���qSW���(��"+=E�MʺM|��u����4e�u����~U�Gڝm����NM����V�Cd��t��ׂN�rt�u���N����_�r2�����g���^H��B�2��� =P��6��e�S>!M�Y%*7U�M���*z�s��-J�	ڼw	5þΌGX_��P�1�K�5�WE�{t��9�7�� �:�5�����KM���/�c� �{\#z�^�-NJv)?���:z� ��)�.$&Gs*�{Ջ�$G��c���"Fnd�i�m����e<�(�?��Fٮ���T�8���f���5�MWG'�.Z��iȈ�V����{\�L��Pw����	+�����K��[p�.F��U$׾"^��"w�hL�,sg`jW����;���4���(H�E�3�,l%�,Feѱ��Ҵ�7?�:��xXk~s	V��u������9�4Z�Xӥk�B�,��0�eq7&��!�w.�q��?�1��b%��hЊP���/~.�A#}��Mc����}Wg���vO�r�y~5�m=� �ۉi���>9��	��"�a!j3�=n����3ӵ��A+?��tK�pӝ�/刯�?��y����U�%������EV#g����A�]�YU�N��.]� b�Qᾃڣ�3�4<�O*EźBk�'���H�T'L2]pPT{�=���?ԏ׈V8��)�9F���V��uE�q�:�%��o�P�_��x9��� &azX���YمC��2Š�Y��Db�4HȞ�&��m��w,t��a���ݏL�B%�*h�R�'>,]�|:&B(c�_�W��	kĆK�hV�6P��)�%�g!���6�����[q��)�O�o�/��zX�ki?���^NX/�'y�W�1���+5sѢ
?|�B�&��/�&<ȅS�!����0�U�O ��l��\D���K��O�m�Kl���ۊ"(1xA��t�k�|̓�W)o��6����y*�"�v�����RU�Du+�Kf`3�)�ȓx=hU�/�j1j��p����K^N8mg|:���*X)* 0V���^A�>�NN�M��0b^�l���Ɲ1��e�ء�[�s�D::�䙚0V�F4��q��&����^��lo�3B�ė��]��kR��|���,u��������?��~?YK�77������nQ��v>YZ�
B�d��|�s�=�x�C\���ik�Ŀj�Y��uQ���}%��*�G���b�N�]�a ��;�IIA��R����^�(v-��N��4lҗ`��$���6��P}�ԇK���K�ߟ��r�dZ�6Ե��6��J��A�x��mI�K�@1bw_E}�����jυ;��w�����H������3��1�Y����b�NxRH�sO�7��\�r�*��P�-��̄��ɚ����:�����`g��1����
s���_m؏�>Ǹ�"�߆:,�����߇��8[�dτ`A�h�qsGQ0E��7p�Lb��P�}p�P>�Iѥ�A;9!����C{g�v-�R���Q2J���������%�NZ��� lB���A����d�5k	}&���x�et-�vsQ�?G���;.10�$�T��녊W�,��Nۡ��5HMg�->���1-k� ��Y7��I���{}y�F�9��d�o슾�~`(�B˭?��H�>N���.I'��)�ڦ
g�V�#z��P�{ʟ�
�1�j1�A���W���Cb`��Q��[_��F���mZ���y��@\�:������?���ŕ���E,�e��X<1��0t��qz8�`<)X��2�����s!�&i����тz:����$���M&��~��.���?�Ӆ�;`Rgo��xO�Qyhܝ�6G�����w��Opܦ�ZRV�*�"MTu!zM�3�V������Q%�t4y��H��֛�x�D'��I��n�6WW9w���¥Gt-��@���J%b��;�C��nJ	��Z7S�j,i��@�f��6H�I�`��K�K�s��#-��ٖ�C��8��7b�K!bՃ1U_�s  ��=}6�YH���b�_�{GУ;���������jJJ4E����Y}
��|�;`<���b����d���biWD��	R����}���7��=�K��.��v����M�Yݫ3A=����"���˲�f���ޙ�/^�����Qdb�}�7_+�{tE݋&ޮ�)~\�6���O}�Ru'���8���>�%��d��{ uA��G��c˪����m=���������o}�J�H=��Xͯn���������'��ޠ���7W�*m�5׫�oyD��W<�T����"<C�S�}�ˍr�|�Z-?�o��=���\�	=���p���c����^,A�B����)KT��ƃ���Hr��t�0�m�h�k������B�`���|����}ڈ�~9�	�0�|�mC5���"jb�2V��s�dĞZ�@\9F�V�Y�vw���{6u��k���B�$�֧^(�%o�r�
��4��3��ʟTq,8�aqr�,�#U��~��*Z�;H]�� +����JO��U����N?/nƫ*k�\����ة�v�[���t�u��8sH��}޿�Er?l�6����!f>'�ybϸ�Zm4<���QV���J��9^�H~e��&��+#��|:���}Ͽt�V{),wG��t�_�b>>TL�7��qR�¦=��I
��(m��`�dС\���(�}����pT_�$�i8:�A��V�~�v+�|�R7��Pw],U��ژ�9����)6���cD�TY��D��_��3mMf�ܕ��x����gn��:`(�H"7�1s4٦;'�l~�� ����]��;	ykO�&��׃;��>'XV�{v6RQ���ʬhG��Oz�0���%�	��u�Dڏ�O�H�<�˶�Nʚ�C����X�_��*�(;�@zM��D̜���{ɂ��b;�	��蒹��%�:��v`R��Ƭ(�;�p���R��h���C�d�H�Z��2˭��� �˅y��^��6ojrs;�@��ͻ�JC*���Lr]�? _��ҩ��CAW��WY�+��M] ˡt��� /%ʋ10�(�`/�%�
�����ha�yV8f�,s7q9���]|F��qEs��ّ��Z�ޚ�&ƻqҗ��[��[U�W��!��IVd���:��S�u�)�T�x?�0+����o��	1�=÷�>)�[���Z�һF��t�
^�����J�6#)E�7*�Y�ӄXӺ\}�|�؆j���/�2����y���&�m�f��V�-�~��.R�G,��e���CS�pӯ�H�~����./~�z���$ҽv1���S���>���,�s�,��>?�����G�H�Y��y��(�Z�S��_&���d�����:���X�+_���ް.��	����fqh��&��j��� 9�A�Hq�Y���K-�a�5H����;뢇؃Fӝ���f�.Į3�2�v�3KS��d7��EA���lg)�}4�x���I�`����<6���j�ms90����"33��t��a����vۑ�	�W�z��<����Dr�j�\�qi��*��x%��i�o���CtΎn�e�sh�
�܌�Ȟ.l�BrP��&$�<�ЬBAa7n�\�vy w,{TC�Y*�Y�\����ME慚��R�Ac�k?�����7��ǹ��5�p,ee57����H��+��ٻ���hP��!g��c�m���|�]l/d����[@ࡶ��W��VC���i���@��-����Y�/
ۭ�g�d]Hϝ�l��	]E��2f�U>P�k�����'�pR�&g�EC�'�3��;�Az)�%rI}%�&]�8`�V��a�������~�T��/�ꍾ`:�rI��'�[������ ������'Q��3��*Q�7��
X	�: ��"�J��|���>�{K>�f�+|BlkO��Q���x TI�0H��,:�|6�n޷%V�e��h�$�e��ޒD^*KW�l�m9
h}ia�6��{�L��Sv=�Ǒ�S����I(i�@x@�w�^\��E�OT�g�]βb�&�ӈ�����)��v#�!�J�A)�|�����^����rl�Y!�]��U\@Ӽ9B�{������ ���47Baj��<�l58���A�4C�\�r1�Gڙ[��m�׸SnttZ�'U���h%�jh�ߛG���b4q���H�����9�力ع��ߝڨ"��,]�o�@K�������.�7�`��8�*�߿b�b�j�l���H��K���J��5�\�0Y��b��;C�����c�Ҧ\��P�<�cQ����g�k%~�~���ZQ$ڐ�ڞ`Ϛw=m�>U�� �B/��z�ar����X��4}�
�+�jhx��a��0�-��^�˴��9)H�]��(����5�q4a���1�1��}�oS����!�,�oל�D����K�0	�+��ü��1>�%u��`��`�΂�`�OL��/�.���G:�I�����p�Y�',L%Y0ޥR���v�Cvzb*�HǢ�+ X��t�®4x�,�.wu��z�.�����ڝ�D�5KXh"[�3fW����o�����A2�D����R�^����Jw�KD����7��-���ty��!U��.ٙot]BH$��Ǫ��U���p��h_0���|J��?p�M��E�̫fH	y�c���a݇���Y
��'�3�.����4��>G�7h*��
t1���ZL�X%�� �O9G����J��g-�T��n�A�}�itB�$�1�ɞ�]��D%�Z�nB$({�1,m�6z� 2��fE��щ���k��yw�Q�;M͉gؒ�px�/���v��7�o�P�0��y���v|�jsS<�$�;�j`&�u>5�B߂2��<�@W��&��/���e�$���i�e;�q�Hqj���%�#���I�&j:�Bà]��A�r��4��W˄4�)�,p!dsu�1Z��v�������x-M���#hv=d��H�&�վ]��@ơU�3��+�N� T[����n��{ q�x���{��Dfqz�ƣ-��R'> z�Bɫ�L��М�Ҷ:��Z��x����_Y�ќ�خk���E���|hB�@��^veOvx&$U�E���A� ��"4����-��|v [%s��k��g�+�3Q$�.�|�O��]ƪKb�]���:G��ƀf�@����O��_���LΧu8f/,���6��l�_
/`�K����sFk-��O'ȴXd�6��:qb����NGՁ��?���j�|S�����r�*`��|��\v�$L�h8�F�x�"g�`�ٗ����=e!�T4w��`���"���'�� ���|��GOQO[�	��a��/3N�*~�ƺ��a��Lԥ���8�8���|�zn�ޓ���,�����z�j�P�\��;��$����h�o�{j�o����yt=N	�Nh^wǄ��%?�8,�V N���_�����VT���a
s5������µ���X
��p��C���3�_ ����s�P�Z%���Բ/X���9f�c;1^�|O�g���}%gb�ߏ�/pW&8�ú��8<���X�4J��;�C{����~�n+�}�r���)�Bp�����I8��DA�b}��A&�Ӥ��c�ó�d��c�zV��[�|L�LR鵀p-R�4liZ�٩��ٰ�f)��z���u��2�_f�*�"����2[��y��f��_]�XpJ���\I�sd�QQ;>�@RB�����x.�\-��J��-�-7-��?��E��Q-VH�Rw>���O���[�t N#H46��o��?Ʈ�KJkrm���̇*�O�>g�	C��[�E���q���mR�L��q���*�F:��M0��njFw�!�d�K{l>��1�oD��p�Ow�j�z�4��pe�+QK(O��L�`�wYى/�A}7�5����3�h�Ђ��I��^� kH�ߟ����v��R$>�F����i�#;o߲Ne�6��)l�0�q�Vr+3�^��B��� �v��0�x`�{O$c��ׅ���P�+���Im���{{�O������x����h��'P|^oǯ�H���c
ng���wq�;띒�X�W���@���w�ᏨĠ:�0#��#����/|0���L�kKZbP��rZY('��-V:s|����t+�&�Vj� ��D�s�\��BH�l�c`;�G�6%r1Hw7�g*?po��S [.�1�P������}��w�jp��=|/bb-���Z+�>��!���8Z�&ͦiR4{��6 Dd�2�6O��"J����H�apr�!ϊ4i^3߽z��# U��(Q�ջLމMhΒ�?��j �[��}����D�
_}���ʦ��C�/�#���YyA�x�G��bw���a��vF�T,����E���W���o�]�1@�E(<�t�'�x��D:Y]n��l��{�U��3L����!�Y����ܙ��N�]�t�3(@m�������������DR�tP��[�ͅ�L���qD|��{�2}�п��pn�_�XbOy&�%J�񠭝�tȳ><�0�����������Mv�Q/�t[)z�)�o��ir���!��a�ئF�ȱT��M_��B�� ȉd��C+$>�	��~|k�Ų��w1��+��'�����0&?=&lD0�v2�$S�s!��7Ü,�N�y���� �iP�&���_��G�`<�6&���\X{�j�:��r��(� E��T"j�`k9l�Q�2+�
V������Vc#��E�E-��<`f�X<�RP�E_���j��$��I�"�r���	�l������
���7�a9�1�X�5J�q�J�xGOk���"���D�p�6�|�V�V7x:�-T�U�v��[n�}�Zs3��NE�J����
Kf��\���-�Ǩ0a[>�ᜭ H�*�"?�:�J,��Q��o���7+�Wp1/���Ek�ե�θJl0vX�:��&e�G��/C�d�����FD6vz��-B h|t����D�:�&4��d(���tcc��ܕcg4�Ѡx_;�^NØo�:]�K��y�XI�������A;D�8�N��]�w.�rv
6v~�Q}d�;O�#���>��s榌���NΚ\(��b���#���K'MVB�	Uǫ�M��oVz��iBk�4򳏳J���<�C��	깭#b)3>����P���>i\q��e~s���Ԙ�#�{������̀�쵤�AP���s�Jl^���c�̱�����B�����D��z��(Sē0f�O)���Ǉ�0�ˍ:a�w��?�C�/�u��F��\�bDZ}��o�=�L\c���G��$�1v8�7k	�ԋ�uo�;�̿���:��c��#�L+ `S0tQ��N�}� �������x�yd�@� �tK��%.o��Nڵ�'�X\a15��e�:D���F�d�[)zUd.�/��ޭ�~��ʷ?��tSۋzKQ ��uL�	k��@@�y+�hg�BhP̞Z:�DY�1��s���KE�p�	��ܭ�tC���(c�G�E��8f���tJy2��cT/����W����]����5���m�$�#�)!����zX�f�̂^6��4���n��\�^�/���e"ͩ��Y���%���O42��f����8�XΔA��/K�$�
�Ū+�3��u5��:��J�]�a����ӧK�d`�}���1�)D��9�|�^�Gp�d^�e����?f��u�?}M*��kV�i���:���Խ˯�� ��8���lH�>��8��С��@7`[(���A^��d�0�7�.'��<!�m��p�����&�C�+��ikh��0G�C0:;c�����t��5Dm��ښ�(f�ύc8��M��Y][�~h�[� ��R/f5�k\�)��/��v�}f"����&��g��ʓ����Khw[�3��l�Q��h-M��HC�dԩ�{4��&�B�ߒ$uƌ�@�H�v�ښ�2Rp�����"��2RG��:P4u�%���phU���>�������|\)���?m(�FD�g.D��D�x��w�։+E�\�����^�ݘ�u���#��"C�A���zR)�
�Z����e�O_E1�ݵ+�M��Kv��y���+3�>����p�Ѭ�.SU$�� ���	�h?
,]s �Xf"˥��#t�p�y����íI� ���u9I��4��uo�C�фՖTN���y����Bso�����sb'�?\f�<�%w�����h�Z^���V+i	p俅��� �8��#���:��ٺ�뎜���g�C]ܙ���6���P�����4������G�J��v�D��|+cu%99o�Q��p�؉��V D��d��<V��|�l� ƞ��]������-��SW�4]��:%(V_���y�
OsRn ���vb���h�p���i�㏷���C�
���;>��W~�7�:�O�f �h̞N҄�.�G�����uG�f��4��>��{�	|�D���TYw8`JB��}��SL��>�4�`I��@����QvFK��䟴C-��73G�|SДw+l�h�}��F��u}��+�:R
���r��<��:�uֆ�!3��?Uf2�@�H�¯��>���_vs�8+4$�T�D݂�=��WTLi��ʉ��7t�\�~�� O6���R�%-<�>�<��y-C�m�ϮoǤzď�������-q�`Y�錮���"�����E��s�x����g�,4o�$x�ۚ�dڦY�\A,��9���A��4��L�_Ϥ�g�)�X�YqQ(���i|9��z"W�~Y�DN��$��.���ث���TK���'*��$���֦::ǚ�qO�;���_>[����_'p��CvϲU� �pIj���62ׅh0��Jfy<B�p��쭸���}%���Б��I�\AV�����]�NY� <�s)rh�I杊T�}u��V��/�����(p4���=�|�J��]�"��*H�>39S2��q��q�Y.m;���l;��e�[=d����´H^�%�M�B�U��V`R ���ע���&��F��@ا�hZo?4v����I"'K�����8 �������M}�XeF����:±�ؚ!��4#�.�,�(^�������~l·�<�n.s>����|�cAt| �TN�3$$�{��qn�$��z��V2��Ctɵ)�N�"j��i��-v=	ͅ�6{4^�J��O�{G�k;����+H?�+Pjz�5ء�
�zGo�U����^PB���׀`����~?Ӛ�L�G��Ϥe��i���AWi�?^#�d�]I�Ty�f��?QY��{+k"��J%�T�Y�����$<��[�r7��gZ���g�G/��qnHoy�����N\^��3w��p�[^�%�,v!��0�3Tl`�2���e�+�&��0�l'p��
�y=�HJ��zu_
Ǵe�&� nzw�|�K��ˍŻj'.n]�/[,�m�X���ɂ�����?1�c��QSL��=F�L���:�˾�G˦��v�d5sÞ1��ֱ�����ʤ�]������u5��i.+���&�Xc�3��`�g^5�(V���+m���#^��� �K������:��QAܳl>U蚜�s��Ka�CLyV_̓Pҋ J���`�x�{9o��Z���*+���g�����"��`���KBy��ca�gS��̾���'�����\�t�v���eD�'o��5�� �������� ~&�1j���VHB���ˣ6�-��k�91���!p����t�[����4���$C*%!�7�>"�cΕ� �@e�E۝�'�RyC��35&P$��<�`G����}�Tg�D�nX�dq�M�p����`��C�I1��ԨD����3����a��-H@�52�;n�eT�[/��U��f�$� �$�lS��<U�o�&��a�*C��|�p�Ҕ�1���"�Ha��<?��4Rj�
�;�I��^��ݮ�ۥ{��}�\����5��7J����B��˦�9���J���)�ۍ�^��A���,p�d�����F�#�3��Q�=-*bx,O���d�*�4C�^a�	��J�b��J֭<JF�7���X#0��\�GSintu��ղ����6O������ݠ�Y�959���h/����ix)�MO�Og8���}�ʁ��� ��f2��f�^��>�'I����l���lȖ|��>P��m�oV���=��G�
;;���fPi���e�-l���	�.���J�r�r�zq��t� 3�U�ޣ��<M��.Dl��HH�[/g�K_�� s�0�XQ�@Z���^� [Ь�;��D�+�u�~|��U��Y��1@>��4 ��o�� �F��7�S�,;�;x^�`C�	;@]��[6Z�4�> 6�ڰ�\Hl���Z#��7�A�;�XC�H�A�x�`R뚐�� ������ZA��}�y������q��^�G�@��ʳa����}B3ܵ�\E��\�+"ֵ��"YA\:���9�G�`�����[�7�_�Ι�ﺗ��w��m��ڥ�o(��Z�{I|2�H��n|��l�9����� `��)��G�'��YX���ԧaO���z��b�L!QThQI#�NgC��ڜ<Ev;0Yϖ34��p��ey��V�J���𫚔�ӤR�)L�9>;�Au���Z�l �	hr�w�>��x��|U�с[g\VlnHV[r�TNK��:���)���	�B��d��>b^N���>��	��4�Է�s�\�ޤ���W6�o�s��_��9cx�m�pB���
@�C�2jLY֧8�����+�]���	M���W�Q��xAZ����.%_Ĺ��#�efC`"��~]e~����R���d²���Wp|fyE*U+'��l1[N���!��*�����h+P���,�4�m�!n��"K\z��K&��h��>���w��$Wp�@�Jc��Gc��!�ɼ�s��T�}�U,]ಸH����J�Qʛ�K+�W���/
�2�\�^�ŏ�㱮P�AX�v1\�;���z�<�b۰�j_��t��ղC�C )l�T p���g����0pΒ�~m~��'" �� �Q�K�=0\6�X�u%�4ZP+����]�*Ω���P�f\,�̬1�Y� ��YHؕ�M��*k뜾6��DO�=�k��ژ���_�nZ�zAQ;]2=87��-��pi�X>����V���u)�5Q�e ȆW�j�}&.c&����׭V>L0ZqC�Ț�p~^��.5�=�|��17e�XV���u���=5lGI��I?y�w�Knx�����B�qX9���`o�A�m.����� ��jZ3H ����r�-7��7��V��nޘY4����DcYΎ����<�=�����������4���>�Auδ�	�t�[Hݺ�	�L����r��������(��RE!
w ��{滏K�,�r���P���4��|8fu�T
\2y]�1: "D����O"���?��Yƿ�t۱>�M#��!k���yw ��G��  �<�i �EL�{��s�ߤ1Y3�.S7Rך�u%����g9w��Blvȏ3���]&��ǎ�C��V��c8�_a���b�75v!"��`��H�X�{��Z����br��&�=0z� �*���F����߭V�#��b����r��-a��*����4+���ōg��7�K�?��H�7T�7oԪ���^�)����:���f�$EgV@��`38LZ�֖0mSJ�9��%�kA�G����j�,��
��ٚ״�N�Ͽk��jJ�����}Vd���_CA�YpǶh^@�
�
o�i"Zʩ"?o�1��v�Z�h��#�vU��<��ۼ��o��ݾ⺠�pǗ��^�~>Պ�)��]-�E�4���}!5\`��#�1�g��j(&�}�Gk�[����ʬ�[Q�Çm�r�U{�� d�j4�����-#���
�z���;0=�)7x*0�6�X�Vvs�/eV(��w�̰���+����\���:�l��CðrWi��5���hϒ�U�&�zSԟ�k�ՍQZ�vF�ˍ��!�3Z�h�L�H����0�_�r"%nW�Ź�=��+��OX��
~��M���32p�i�|qP��v�R��EU.��U��S��Ԇ��hb-0��!����<�Y4��|O���u��e�46��|��ج�ƀ�U�.5�я��n��~�cX��A�����D��J�?���7����-6��R�+,�n�.>A��������5�R~0�ĕ�Ú/�b{=�/�0��7�I/McK�U�ExH�g�T��~X��������6'y�n�t�oPuM��j��;����e~*2�"#�vA[4�<O5A�`�����Ǣ��8a2Z}R��\6� �?�+���=�zW������4�_����7�TU�
QW�%�%���F�<5����àԔ�[��x��U�s�)�ց*S�S��p(q6 ���*��ck��OB���lH��1wukl��nX�?��R"ǃ I�3n��L�Uf��O��߉L�O#����39�ڪ�	%�
��f��F��e�|vЇ�?�R��q�/�Z������F~O���yY���6��C[��pq�$~H���!	��,
�B���9l�OV�F|�$طBqD��(Zj"�?�i>������ 7�f���z	�t���s���!o�h3ۈ�UZ�s�
�,�=�I�_�Y����o��F����ղ���ܷ2�3+��L�����v1�sX�8$C�*_ˍ�2���HYxYء�7��sqEӷru�-�T�qS�wo�3�K'�p�ÀbA�]$�P�]�:����4��1$xV�V��;��'�m(�-� �?�,�@ Xu�*l�{����5,)�E`��_
��O�ǫ�1�2`����ңE�)%��4F�驡^���ř����]y_:(#&��C*<���fO�<�����H�U/N{��2���T�4�'�H7)kW|�Ԇ��dm��8[��:��I��������_E>K��ƕ�12����u֦`�U3����Z���r��w�:/�m�+���uU������x�\��4S���m�I��[{���^�*�K����k3�����f-���Z �El�o��o��3�K���v ԘM�����S�`�j
��^��(��Y���:֬���+w�(T�<�V�1B}�Y~�p��3i.\/�Du��8�PҼ\!#kz��R$��k�Y�1ն���'�b-ICԎM�>�Q�A����={�I�˳H}��-'Xӹ*��X����Cc;q�����'�2�c<��S�_��y��T���K��kvQ�Q-*�A8���=��WO�H,�z������7ݻ�� ���p�MmO��������j|��*�H�d6}>R��<߻�����M��*�����?�\���Z�D���	�����]�j��?�Y��y�ÏyޱW���\NϦ�V&��Q����P��u�_1�.�@�F\�V���4b�5�V_��V�B� �80��Y�'�V�}J�L�-�[o�s83\�03���SU�&�r�Rg�bb0��.��[�H�O��gľ�,.��br6�;�D�N���t
^��F��9«5О��V���к+�KE�f���L�4U�J#�;�F�o��Sa��H�CĄ�n�k��׎EZ��,���`�!?���z
��{{����E���I��*����>�/dgDF��t]�USژ�������]tT��d�Sn�1D੡������a��L�8�\?V�������W�}J�Y�3g�O+c�¢���a.0HҶ���pY��͕?F�.wֿ�ک�<��z/ȴ&c�<�,"�U���u�N��o���S�Qqю�v Vd�c��*)*����ג��c\�Q��c��_�-Ю�z�<e?r(���!9X-˓<�1��,H�$mѪ�1m�,�B��6y�o��P��L�ӁɯܒT�4�<ҧ��]nT.��4t�"
��މ�su��xٓ�3�Ʌ�nc�H�_���rK�?�k�g��bv,o�F��h�AR\yڧ �r�綬�L|@r�� �ɦ��8��R��#�j�.�w7����jf��a��R'�#�K����ŏt�q�q��S*ea�k+�FS�ne��u��&6��
���F��L�wFx��܇�֩h���P�Y ؽ��>:�6��k��?�e������S<}�.�``}Zh��ZIN��'�q�߀U�93y�/R�K�a�.�Jm���٢�������śN����VO��� �����܍^�P����w������`�ZۜY�t>F��U���;���L�{,h��4��tv�������t�,�v�1�s*ׅ�@
C��>�� `�T�-� #��>{�Y����U��heN�����w||@,�����Y��$����<Tj�v����H�|K�mX#�;E,y\�eC=歘������HP0Q�q�-�u�<�녠J�T���WZb��?�`���g=
�W�'�uo����|Lo_õ]^ARBOg�������X&�ڃ�IJ#|����
vߗ�����Xd�]V��|�般�i�y)��b��s8�h@�ًn��?��i����'2va�;_5���,u4]���ض�V�/Qo�X�|BOiK���~��) ���
V.���=_��uܳ��q�ih��*#?�f�C>���x�ub�%�M�
��K������u�Y��U��v;
�^�4���F�\�P��������Έ��Bc�([i��L�܋c��a�-�$�Y��u&q�����c�o�b��o�Z`H�>�KW�CᒘS�-T�p�N�iZt͐��l�z�!��OtuH��R6-�U��� �]��$Y���g  v�����l^1��5��˲��Op3qw����f��:����9�[F21��<<y�_q��=v.��A��h(+��|C� )�|���=.�7�LE�%��?���>ߕ�L�|�V��F,�r�D?=�;o�(�q���dO�����w|�:���v��h:�7��˽�T�a�$�m�t���W�� �Ri�?���ׄ0��p���Yﾯց�x�����-lj�S��jf�jEoh��E���a�ʔ�0M�x����B�(�U���4f�V&�	K��_�sg·�u��#oC5S��
:��_���sG�t�t�K�rw#�������ig��dJSdή����P4Q���pV�X��~�K�՟<䵉k����l1���}l��hW�Đ���V:�m���*t�NOnWm�S�|�Q�.�z��8v�=\��:�4��PLԊ��
�0�yD�t�1�����ӣ���=6Ό�G@�qM��=_����8���H�v�Z�"{4�w� �)�����V"D��!�Ơ���ͽ�!����l^J��~-�C��UH�|c�[>�~t�<�4�s�W~EN�SK|�j��z�x�8��?J��<�ʩ26&��f����[ty���9�/�֨�N#J�~���~�J��ӣ�Z�=�#A�]���?Zr`�vIz%<@���?�Sdp%Ja�E� o ���U/�2��2o͜H��,H5���*�9��7�����C��h�JO�����d���/	��b���!�Q�a GJ�W�*��s�g�L����l�#Bc�K�
�����Vy���<�Zl���Nr<x��VgZFb���{h���W$���1F��\�3����1[lbGԂ<�<���"s�e6��&��A�F0��N�:^���d'��R�Jg� �E=�KySF��DԞ\��3	+6EmǬ��#�B�m�;���^F�v<�����g��<,�Wj���"��n�F�P� ������W��.�����T�*���!f����ȥ��w���ȇĥR�? b`X���V��ː�����xRc1�U:&�=d9��s���SZ&�u�B���a�����+�ZĤ�^�=��L�S��t��$��vW����j�~�clHDWL`ꮹ�`��������\�N�f�>"�86�Q���t@"���v%���eKa�9�����e� ���G�]m�i��0h�I���5�;�U��Gc�N	�n{�(wǫ�������gn���6P�[�YX-+"%����ˣc�1x@��SW�_:���hDt�ZV�CD��O0�c��O�8N�1�'�Uv�,$
���(�܍;�K�B/4"�k,_��h�֪+=�U]�k�7�,G(�Շ6�<�W� �%4ܤt�Y1<5�0]&���-���:!1�r#�F�;պ���"w����[�>%[�V�r��7�?��͗�^\�=�����/�@L��P��V@4�����$ؽ��@��0�������x����I�A��4�x�A4P�2"ʷe�_���"#5��Ew_��2�f�<(L�|ڋ�dF�mh�/ c��\ؾ8d�z|@xKSb�QG�v��9:��L�����}!�9��I7�����T&Z1���ǧ;-�|���]�T9��z#. �$p�\%�z9���Uù~��	`8s�.�/l��w��Uv,�=���J�M);�@��;sy�����t�y8��e����1/K?>.�u��Q���І��L�Jg0�߽X�s25s_˕�R�6S�/��>{u��Y���f�U�6v�$�ZG���'%�Y&�`�u-h)I�ed����޵2ױl	'('G�5�fn����X�ʟ�����o�;-��{�e�[��`q�~���ޑD�p&�lr�e�?���C���yy�|֏c���)��s�nM���6蹢V��v�@a�tČK-鳧"�{��k-ݣ���B�ڥ[��g�u��h�C���Qj��H.�ZUa�N _�gɏ���U�/��	X8{�Y=���~5׺��aT�s{9�!39c,�Q	ab�b��Te��i��
o[}����x=ڵ�q��Y=�%I��G(�{���q�(mx��
^��#!�[��!����J�GK�h�%��4l9����A6Mj�Z�t~�	(��[jR@��n8;�3���骜��+�o���L�%��kS��Mv�K�A)n�?��;��^7��`��G-4��:���bW�'/�}���ʫ����.Z����U;mR/�D�qÀ31�$-�oI�\쬽}��DJ4JӅ��P飋 �vm�P�B��u}6��ۋ�
�<��%��r�����3=Ѹ�eR��La��6/�O�3w�F��[�nj�X�	�8o����1� ��8���hꕜ�^�P�گ_ڻ�����)���X�f��ZtQM�L
��;��j."]�-�ۧN���P���i�n~O��`n<wEN�o��*ɛ�mR���;�e�&(���2.��E��j)`�g�=,j@�-��a��w(Vч�i(S{�<�"ue"ΎD|�����o�	���ޏޗ�tKz��^���ѻ��M��q��1%���FDmм1��g��o�9�a�	��q9�x����g8��L�csnKt��*≇�a��U��]m�݆�As~뜰�fS��=�����/�^�Ф�Hl�lj}�>��{�+��	#C
fzPU��C�ǖ�h����W������E���g<��U��'���Kn����;��Ђ��bQ�<�'��=�����|��o��3$��[����vœ�f5Ec�I��-O���L��Tp'�*��\F2�Mx���ǻ�"�,�0ŀf�+����)l{ڔ�H��*��s��ێg�UQE��Ys~ƚ#�-�n���[�ka���h�������9<�����!^i��g[im���Sw�j4ɸ|Hؔ�O������/�3��ǿ��v�{q"[a�R���M���\��,`B�❲$��=�7��k5cX��2v�xYb�9�2uׂCm����f��!�2��+:{���އq�z��^����c�� ���Ч�.�<X|��O��$�ƈ��a��]EUVњ�n��2�^��>l#I���^��|zN�5y��E�!��Ic�8�r��/�V_1�H5�:�S'�g�苯D b� �c����JM*}k��S?c�j����v��dp4MT8��U�e���) ol+*b�4�Ⱦ�T~s><$\�e�������rc ��#?z��e;���π�#�[��_��t����5�`9�*���8N�7K��64Za�j��.S~��
�W�|�@�|z�a�Aa�'�R%߱�\b����_fg��R�6E�e\li����J8ȶHU;P�̏*26(,J��u�_���Δ����l�@�� �Q7N?`�`y3�)q���r#��03�E����}`�\'�
���Z#�A��9�����#.ǑrХw�����C~ȣ^�<���~�{��RU'�C��2h�����|�#�U&@F2�ޝz�y�킔/QPm��ؙt����ZotG$G)��x��`��=dT��&�bO��@e��z�_��3:C<�́��N�~�.��W��1�wĪ�/[i������X&,����\5�t�&��ޭ�r/l��l8[g���D�!���rMO�ۈ����I�Ż�n�?5�EV C�T�o�.�w�H���,���#�E� �C�q3z��ᶙ�z�<f��K;�o4�'77u�m�^'�]�b���nZ�e�	+��j[N<\9ѫ�!G�
pF�5�q�p�@ʥu���1��{���ѠI�v�x)1�i��A	�&��I,�gA�
҈~3 ��-a8�;��߻=�ubGo��-$�^�F(U##d�w��;�;�KX���Dx�y�MkVB��P�6�S�8"&s>�'F�7��"�����i��O�Pj<�k������S��l� �Q1Cnn�r�P��G�t0����<1Z;B�S�m3�Y�o���^��+�c�s)m	��k���-��'s%��e��R��%�Mc�]��G����d��@ߋhO��܄$�;y7h��t�����'�B�V �]����'���//u��.�����a"�G�� ՝��XX�:��4*�W�ifz-�+�� �/E}�u۴�iu[�v��Oh�R��=Q4��y�����0ߐqs3C���XW}s�Rr�u�f?&K������~���(��T��n�=��r�ne�B$�����]w��\��0�S�l�Y����0w�b���fx��v����6���ۑA��$X6>��^�� ���{�L�8�UO���?Ӳ@�v�$���T��"ᦦ�UO��E:��~+�R�]t~���1xA���+��N��fʢ]�*)Z��06nZ�!h�G�irH}|���-���B|HjS�T�[�i��K��Z��V�]f�s,-(-�_���2�M��` ;ۂ��h��S��5Z3�:.{[�y�����A�E���g�j�;����Z��v߃<��@�t%i�rJ�������P���t�3�Jx�H*�����VF�Uǫ���<�k�z�F�ב�9�HX�z���0U�|��?h���%�]ڱN%Hv̕�;�������?�� ���b!�.�� Q(�Rۡ����~�U������c��:BV��s��'��"��>zb�Ft�!N�������5��<��Y�b4�]*U*4��`޼�57��yd�εVI��[�MM��M�1zյj�����m?�<Wlx�R��RE�����w�"�<tGc.��������u*ބ�ǯ��9�?n���9}��M5�MKW�4��6Y����M�G��$V��ߧ��mg>�1���I-�?Q�����須��]��g)x�=�[i�~N5wT���k+*�q6rHاA y� mY��%���ޛǝT�{��>��~{)�s�ߞ�5��wz���K��) tp������JL��Y�= ��� �4��!�Wa�1:����8����jBE-Ц=�!�V��㐀�[��#�g�O��U�g��:)��pJ!��:�bV
Nf��Mq�@��|"=��a�54({e�~�#ooi�⌳b�:eg+�~p�P�_��(j�X�q�|e:Q�o�õ����yEy��>�B��`\�C�PTz�ZMlr%w.S�6�Lp�K������ӣ����2��W�6n�KC������ij�5��'�6� `k��<��Ts,��|5V� "����_��2�u��c(2آ�����za3��g�m����d��	WM� ��C�)�:?��7�gd��!_[��!!��dٔ�w�Xճ϶��0 nR�	,c��N̡q�Ǭ���tۢ�^��s���~N8`�jJ�pT�e�����//\�X3���=��<^M��r�����~UL3q�����疃�J@_����\�7v���p�\V2��h�q9\X�s�#�'Y��'�Bt�%k۬�Z�L���u�^n��2�+ j�f�x�Y�ṑq|kN'����ф���A\��U�3&��XkJx� :p�"U�&Wt1�P�?ڧ�|L��0���{pI�@��^�$8W�j�I�8@v-���w�u�ێ�'�Z��_0W�eW:u��]pl^4�/��4w�\��[����1U\g����h��k]�qvݣ�	���A��&�`؉��m9�}TJzl9�5��&�����HƠ,޼iv��f��p/p�Y;&j��
N^�u2�L����֖Y�IN�H#�YW���XJ32T��ے_�&WJO�o���H��O~�-���?f<�%����G0"�Zŵ���s��S���B&�Sg�Dzc�RA֕Y�k�I�^�#�bv8�,w��1����ݚ^�Z�y�Vs�?4)c��JGM8�d�ъ��-��-��]� �����{\9hS�sT^./	@5CxȀ�.[�G�Bs�QvGzds�s�w[�6"��W<���@��N�t��G�v9�Z�d����[���䨽ذ� ��(W%�o��_Ѭ}߈l�kD�q��ǶNn��$~���2���1`?�ݦ(/Ի�%���A��hﯫ7Q�>u�BN���R`��=�]��m>X:�4�(�=A�4ԛ��2��9�(�SC*�fSX��G�7�0�jHK�tt����Ð�� O�x ̓�ܝ.ߚ��N
Wl�W��J��t��1u+Q��r�^�7S��V�/�Ǎ�jH�nQe���+��}��8�}��Y��$b�FU-�0�I�/��r�C�\���m9Ԍ����r3��&�)��m�-cܤ�V؎�U҈I%옍���y�S�_�U� ��wU~{=1�}-�����G0<:�k�m�0� ��)ڜ��5�*d��z�oBEk�o�-�p��DG4��R�,�A������|�f�N#�*_M�rr�(k���|h��7:c���Su�t7������Q3�u11���EK�6s,����&����i�`����k	�Tlw>���C`�u�EJ���R�lY�yZl�t���U�hM iKb���D�p���:��Rd�Of1���;\�'��10t�h�B��PٛxG����~����c{���.#�d%���q)��zH�y+��<NQ���^i�÷B��AP�Է�eq%��mY$�ҩ����*!�Y���4�����q�3=��`�(o@�=Pv;�����g�p�K�4Hf~�j�� �#-X�􉀛�9��(Zq����U���T�j�u�*�IQ���@_��	Nδj��(��u�0 [$"�k +yx��RÿoK�¿n?iyz�2���|b܅V�� 8N[����U�Zõ�`�oʹ`��Kz�2"����=������ޟ����_A\�5ȉ��E=ZOɞ8�b�q��ȧ��������..O�����5���i8��KGn4�t�o�ε���,)J�h4�g��Hӛ�%�����!�)�̞u�O�.�ԓ$o��\q�2���~�QEr�@��m�=w]>�g|�1n�w3�8WP��8�?8�a8��3�J�Ѓ��N1��F�5ذN��*��!���G_[0�܄k];rF���O�~P=�9�N	�P^�yvK[�[D�J�h��d�F��(H�@�%ɘFk�ۚ����!���i)fc��Hoܐ��~�`�R�x�Jf������m��d龆��G͵�xe�pӏ]� ���b�Z �
����d���12�,u�C���"�����
�b���,B�К_?֥��ug��M�"������<�m+��rK�lk�K���tW<_٬X���֯��~��V�`�H�i�d�5��]1!P"7���X�tV~�qln�k�O�9����:H�Җ�f~Am�QG]��xq�UĈ̀_=[�����`_Hz�!��'3�����z� �H�c\Xcp'l&)gl����$�MP�d���~o ��JTVd{	�Y814P����4!B���������$Hz��C}x���}ĀP��T�*��r9�Dws��h7�*}w�:�v���8��ď�e|�!�].aE	c�mv���J\�aXߜ/�П3Vl�u�W��q�9<�j	��^W;�_���U�ȅ�{YG�%X1�� [�tE�b{3���5��A��H��a�RQV�hp3ÞPܬ|�:l/��)ܤ���R�&
�b���o����=ǵ
w��jz�%|A�]Щ
�Mj�{�Dy�U��z�2@�E�x�}Pk~V�h����~B�U㩾�?�v��~ZUv���O�{��0���Hw�T���F^��6j竌�A�s�U�G`Keei�lt��r ��cp�7�sI��O"�q:&���T��]v/��g6�Н/�� -��<&oʧ���c�g�կc����E��܌�;q�'�(�L�x#l�����6�q+P�^J��;�[Lx6��"��,o��WBۣ���0�f�L�P�5 ��rh�����IؚB��E��ݾ�x2�>��GS�|�`����i�2x(�qez�	�0;R��`rM�3 ���!����r��j��(��*�&k�J�m��e�za���������Ȇ ���Z.���T�[<��ٴ�r1�k��2!���t��59���$��!Bv 	��{����h�0�>c�
�M��"ެm�OD=az�#����p%Z��o�&�p��W����*гuz% ~!eF+E�|�x���4	�O��>CXU�Ґ�[�aǟ�s ��$K���*C��4���'�TtS�+��o�7���HD�O|ٯ�1��D�cK;vSM�q#�2$��t���p~}m�)�Q�爐\#?���j�v�����8�Z�=}F��n���p,��z����F��Y�vU�P��x]�F����7�=I�5��n�Ӧ����?烊aIxw ��Y
�9�^�K.�h�����i�OQ$/T�]���L5[�.��+���[����PL�C����s):{�w�pZ��˵�Z���I���~EiS9n�޴BMr�{K
��xxu���,6=�TGE=5��1W�S������h�O4'���D*����Q�Wb���~.��8��SDjc�*�Q�h��VV� ˆ���[��F٤%i�o�8�«s(��
�G���Y1�cs%\q^o�2��wm���?��a���N����g�G���Ę�5��lci�>�W�1$�s���� 2Jv�K�G,
O�ԋ$�$�ir?��hy޺��[�mz�ԶB���L�t���{�G�T�����@7{��@���hۯ�����A�W�H���exء�-�1pL@��;i�#C�8?��'�e{|�֍�f�Il|~����d_Ȋ�%�_��s��6���Ŝ��y���H��38!�]����,��70�^������>�K�ؚT���k�4�̭"r|�ߧ�h�a���+4���nٕ�BH�?>���	��)�)w���ȷz��x�OIؠػQ׋/�1�	��&6☧!���[J���Ք9k��RiFb9��
��82BPgְ/��n�ZP��T��S�ɒ6 �6.>R�1G���?�8��I�j��\w��'���{�~)�Ԧķp�ә�O=b��zeϠf{�r�d�h�pdzF.$�W��gOk?*��Ȼ��K�C�V)�z�U����ɕ�	7�J���B��=�~bђ+]+�Z鱉'�8�� ��K�=p~�r�����ګv;�(E�hC6�)�ʅq�g~��7�&"�i֠�k~m�e{oc��^uݘC�D�~���-��@ؠ�Q��Y*V��M,�ͿXes�!k�9C�Щ��{�[�I?X徠����1���IYA�nmLt-�$��8l��*�j�ݙW��o=��3��E���\*�O�3�]ɚP,lH�&������q]�Цi �M�g/f}w�-���Y�t\\�-QCg���Zz���d���g(����fRD/�O	���N�4@�m��jg)z���Aߋ4����3>����p��k�.��f�a4�őSg6p���a7�������
p���f����?�n���C�(��V$�k�g�����wD�}!똮٘����s��+���y�E6�u�i�_�AZ��6������k���$���S��#+�jJy��]1[����x�C���@�/�l�,]W)��XN]��t7no2h ӔK�~k���=�7/�� wg �#~�U�o{f.�!ezĵn���'�%�1xS�r�-��隲����h��O*Z��N��+�@��Vo#��F|�B|��j��幇���w�RE.1_�G�����0'^���?Ώekyz���d5����l���s��@�O�!�w p_�&O���:�u�D��<�%���=r�u]mw���=�ʞԂ)��ͳ��4�l�_D��4����hH�-c���/�k6����L)֥#[�:�e�~c\��>9�1o�?3���h�#V��ȃ:��/}�����v����;������L�Ӽ}=%��9�01Zi�p\`,�+���8�"ͯ��d�@�B����|t��=՜s�YK�M�&�Y�?�x�%)pTb���b1�@͗�EvF#������C��*?�ţ����{�N�+��fB ��.>a�:��u̍����5˄y�����Z�6s��x�����N]����������#\�M�#���Z�d�Y��o��j���:�Y�~�7��F��:�-@���<���T�=��O�4ģ�R�]���A8�r��G�w�+���ټ�H<K�م���ZIFf��q�q��q���V�������,�;��WP���b�M�	ּ!�����Ҷ�U��/Whݡf�9u�̟��)Z���������_�����So{�����N�r@������#mK�
0#��:v��D�1r�f�/m����T��?����C�bs��[xC)���U�\x�}�/k���� ,�Bcf���)�eŢ
l,����o�e��vm]ől�ȮC<�ߤ�"�.Nb����G>�i��>nڵ�P�	j�����r����2�	���nr�&0$CO@�� ��тKb�y3(l����a!�ԓk�k�n1����!Ի�����}+#�9?�Q���T)��� �n�!�ǵk\gJ��*W�"��s\Λ����(�c��L(�K�����!T�QH����Ѽ�q��R�DP_������1��7/��$��wl����Y������R+��e�Q����/p�h���T�Q��`�Bqp�y�V%�5�P;�b\i��.���H�`7du�>�W�S��yy�:�Y�bWG����X�f'��4�=S5�?�,:v���)l�ꥋ:�"��q��"4�)o�ϵ;i��yQj��<�I���"��Z��(bZ�������_�O�W����}�0_��o;$�{�B����?��_XT�U�?+y�B�{�ޙ|���E�
�i\@�؂H���8�^K�AU]�_pz��?���f�5vcd����^|[��n(���[s9�MjOu���W��Fh0��
���!���5c�Ӈ����Mf�J����S�.���ZK�:?%,u��E �Ss\�j��OȤS,��*�вy��l�S���z������Y�U���~DT�����Y��!"u#OZ1�҅^�2����yU�1w�li��SnGsg��y��o�X��R:���Cx��g����Qm�{^��/t�̥w@$��3�/�D��6i�ȡLw.��N&�<s�]��2�u�V�ѵg�+�k�\��8��'�VcOR��ͽ/A�i �g����A��bY���S�I�Pu3GD9�9�,��6%�8�\�!�'ߜ�^���D�G�4���2�h��a�2-߬��/�ق���[��v���1C�o�=���u��?��$O��z�)��� �gU1x� �3,f�%�v��f��XA�<E�=]���a���D�� 1�)AU�SA^���:�]�wo�_Wts�a%�x�>�;VO9,u�:`�V�8��մ��W!M��|�9d���TjE��[�y��RE}��_<%��P�ށ���8߿��B��r"� �h�����ed����ap��=!?|I�~K��r�21v�t�T�tˉ-��7�]7�{�Ħ��[���*�С�H$�����~@�N�#az`I�~��U�Ԟ�j����/�<��ˇ��h?�"������lX��E��ri�Gt�N�S��b��^\�1��2�r7�Ă;!d=}'ȥ)>!C1�[»_9��v���1wC��l��^vI�( �n[ӳ��X�ߕ��1�k�Y�z�9tmf���i��Z��Ň��e�(�M�]R}�GV�I&<ؘ"��}U�V���B�:��OeĊ�qQ'S��	s��-l	��ee�W�*��F��-λ���a`�w(��=���0�g�N�ȭ�6flS���o"�c�r������ a�m�n5 R���Mi֏"&���Q�s���	�(F�"���w��)q��ihf�0�!�q�ЗF���H��|�$���P¹BE>JcCb"��F�� T͏j[�|98K���������i�I���u"-��įӋ����8�?u��W�J{<�ۃ?GB�0GJ���?�Vr���D�>�����X<�$��F�[w���m$�R��1�kL��s9�;i��T�E��i�x�X�k�=w������Ax#�nf���'QT�l?U'��&��8��	��xP�^�q������ZD�G\�>q3&�廴�K��%3�+�����B�ܔ�?�����C���zd��� �S��wj-h��E�g�SC�|�]xfm��eŇYo���w\������7_6�}>��-^n��*����,5��ͽޅ�;���-UH�M�.2�S�Hu�-��Hj�U�H{�c�N�X�.|�cG���C���]Ko�j�*����BW���i�nR�8Z]��D/���" ,Ϙs�����
	�U|��x��PX���� ��1(Z�b4�ܦ��A�z~��tJH���{[/
�H�F�ps���"ʗR���A��{�!N��yC(�e��@���:`�5
���Ψ�������Be2���`-����ƞ���C}�S��Њ{�bv��z����7�ǞQ,� -�����B�5k�&w���-�^/���=n\���V����^~ﳨ(�%��6�I�#���XƠ�������AJa�3D�5��2>���!����L+�4���@*����c��b;��uĸ�T��c��H��3\��d�C�||���rMF�({�\mi,��7�|��@s��W�[$�	]zV��^�?��`ƾ���3#sLw��/%��%&L��R���h��N��;���BO�E1cS�M|Y06}����v!hg���*��{�OA��
b׵�逸s��C����g�]X�.��$���1���D�S��U�[�\�V�A���FQo�����ـ���W�>��3|+K�����V��*�9D�
���Տ�4T���K�}����pff86�f�b}�$O��y���K'qRR2�rR�.~ZE�RMi%�v��q��(Aڵ^A��a�뀳GY�5d���Y�V���JT��uL4��z@'�⚇��^���t�sׇӭ�~��rrʀ�1.��iۄ���O�E�Yx�?����_�.J_P����\������ݕy�Q��>�ÌR�՞�����K�bq�,�q��lAU�MO�OjZ{}��s�����̢hЅ��u%�u�pĒ�A��ME�T�%�$�A�6�o�$�ȨF��W� �I�s�@�͹bV�"P�T##��y�G؈���X����Ւ�ɠ���r�),�=a3kT�"C�2�?y��i[Ӽ�xgy~�yKf�S�������Pw��2%��)���;���J]����M+`
���f�/����ڗ.�<T��0U+0#-�U*��sc��|g�8��^�.J�wČQ����}K�f��2��e&���Zt�Y"@	eB��\��y�Y�!u�l�?�u��+�o��0�[�f�)K��O�ܟ&��_s,�T���.q	 �{�Bf������Ϋr��>M�ێ�xy�GۢB&��E�Eǫ=���ҼQz< 5��u�����z(oހ�E@�A��_k4�Z$ÛpEv�B���g��F{z�t��sj��LS�!�U�8.�������s�x������;{>�I�AOΐ@R�g��ˀ��ͬk�3����8v�G���k�M���&���`3H���r�!7�S��ƹt��)��;mV�o�0�W+�����8���Sj�H�:��䐓M��Ñ�l�.ƀ�(iHŨ<�,ɩL���,$�<���ߙ�(���(j&�s��*VD��)̔��|��%}}C�U��BtQD7	�]C�h��aX����-AhQ��� �f������\k7�c�I�$�: �x$9���5S_��� �y�p6*ĺh����e\��=F�L�pvLC�j��ޏ�����QB�+x!�  J�?G��ŧ��3�������}����w�V�j0�8Ю�*�	�>v�d�E�с�ҥg!����o@Ǐ���{�!��.�a#6�����Ѱ��̷ҷ�_��5�L`.O�u��ls�	7�q�Ea`7?=6N����O�z���h\x�\�(�Q��Z.�yi h�rY��ty�͢,L��W�]XM�w=Lj5�L:�~�$����Xڕ�u���\7��V�_l��"�9�{��4в���7!�@�/����s-L��H�����h׃���&�O����������f(���$�|� ��\��)�	��I���W��RA��bg�/�����m�DkJlv�OK�_ƻ�������g)��}^w·�ϴ"\��JL�D�eȓ�k@�	������I3��Wc��!����8|�i&r��|����߿Cџc�
H�;���Q�MH�㈔}$3Yj���\�F	�TBs�Huϻ���H���{��47�{%��Hl-~����Ph2�-J�fI�Sk,�+��m�@�М�(�e�k�������Kx��=�b}j�3t������7��	���z��=��gk܆�׼������+�$���s˻2MC��#����%���Y�M��}D��*�����Bخ�(h?���Q" ���s:���~�cg�=d 8�#����x�hfoa�	HG�1��R���=���@�R�~^�6X@��{X�>��4❙��e��]�ī-X�@��qc޹��aU��Wug�̳u�x���v1d���ϩ%���g46�������Ή�`����+׾�:;���]�#2S;�sF��m��ߊO����P��I#癰�DYU��ݿl�&:(��A��(�G�(��}5�qg	Ѽ�+�^l�t�R)�h����O����X���2�)h%�G���/���pn���ռ���ׅL��JC�L*��� �U��f�7!U�I����uM\%�5�o�>[g���)��NX���\�Ʀ����=��!#uf����D�w���o��4��W��Lu���(�^�C�Jp��q�k<�����ΐ�O�F��
�\#B�9=����D��$�������X""�h�R�d�W�K!$r}h�Z�b .�?�>.C�PBq�K&����)�Y��7�8�y»͙��a0�2���3(��j�±4�Lʰ,Hh�$��aPR�
Lm��G�:Xw{�������4Z�1	+�~�MwSd�;�����9��/S�M��u��ysLQ��uI5�E� ֏R�M�B<�w[�"�k��E$���~�%F�g�f?��(�� ���g-t�yK��]�/a��3�奍��fE�d��R�(Ntx%,�M�S����P�P��h�dF'0��N��Im"��g����[�6d�Ӽ5ꢆ��Ko��ۺ %˙C���24@�y�c{����Ţ~GKy x0'� s�i��IW�5�|7��X�so�C�r9����;����M�*'e�H�ݕɘUp���u��� a���gym%��JJ��������_���T��U�6	�0���և�\���J-Ј������"��=�sTgZ��&"�{��ڷ[S���)pf�$� ���HY[�K�@��b#�~x u|A@�J�pN�.�:��gz'^Ν��o�;1���%n*�"�'�D��L��I���	�(�:+��^�;#��M�d�kw;�+]B�r�+0uY�R��ƃ[�u0�6��onX�9�<5��UǻQ���v�#��@���ň�Uᷨ}���ב� U mȕS3(�k�ճ�
���T]��D�n{�:�9ȇmV7{|�լ=��K���-_tA�|!�k��юe��K��D�H��>�zg�J樭)6#�_��4	/�@�i\����J�آ,Vw�?W$?˙<�@��&7�,��2�|�K��%�bj�������VU(ᗥ�g�1����g���H�$F?�	����O{t|�M�� U.F�m���׷�J���@z�s��|�'�|�����{NL/��Є��n�:�!K��;�ڪ��t�?d~�̔ol^'N�;Y'�f]s�UPIa�����V�����5�_��2oC�5�#����H�y��lOE���%Xs�Kyf�n8�i�ܝfQ�C�����:��
�g8P@��c����DRo�sY�s7K%�u���� u�mu���T�=�E2�w��r��x�U�˲�`֢ڮ���|G�~J�����Xu��=�=�ǋ�]J������> ��&��	�y�>�)�	�]��1�IE�]��t����0o�$�S���j%7���V8݋�ƥ�l������!PV��r�>��e�ȈX&tv� S�t{ڧ�8���O����r���-��E��#�f����3�9��:4�F=IE+�BS�P�Jl�d��\@�bx�z͋cI��z���6&)����»���q_�$��x�f�СM�j.�	��9�%JÀ'b�$��?xϨ��8�K۶��A�Ez7O�)d�W���~�ϕs��!�1���˫��+�/'!���e���M�4C��5h�����"�;E�#	Ȭa@jU�ŋ���A��i�s�J��rT2��5���>P}�11�,�s��`�=�#���y���f��s�1�E��!#��_��ck��zd�U�/Ad��7fz�@L�!���:p��Y��'b�������%,�o����"��ҋ1�Z���d������L��z��$6�8���	j<'�@O�
��Xz���L��?
1��zɰn��3r]|I�א\��~�B�p6����t$��fkB-��H6C <�1}�|b�wj҆mt�� �B�^�W�ZQ�3��&jk��z��=�&Z�sw�;���6�<�)�S�1����֍�,ļ]���f��*�*س����g섓R,`��n]�ք4���-q��t�tx
�7����NA /��-�&�P7��Ek�b{E����/��d�Qq&1��<x��.��Y�bn�8�C��&�"0P���`o=��3Gg�=��ՌI;�pH>_�9M�qq�5�(��N��&u�k��v�~U����}�2c����dim_JPr��{8dAt���DZ�<׫��LtAÞ|�2ǒ���5�K��K�o!�e�Q܈�;y=��J���!+ꡫ�Uz!y�㾛�2g���_4� �Ё��2_��tx���P�G�H�����X�Ez��U }֕����z�PA�=���YU�&�
�>�`�QlIF�����P�o8s�vy�?�]���JC%z;eO��\��]e�&�
������P?���T^�y�J��Z_8�~�ݝ_�i��������A^1�i�D�{�|���}��ȓ��o�J��𺡂�S�{{�C�A�],(4�����!�2�
k�xC%����%����0W(Wtx,�1j%F��3����������7e���M��f�R�����R� �}�?�D�;a�ʿ�5���{���������'�^�Z�5���xx:_�	���j��pB�!g�*:����{XR�kQOC@����*;� ���>�����໚dǽ��^T�� �[���Y��X/�E�V��1�1`;�ؠ�kɝ����B�tޔ��9?�J�!P�4���Ұ�~V��2�D'�ZT�����6�!\���2��Ic�@��0��3f���0:.ON�(�s�ps��*׾9�<�^a�~�|9V�~���~��6��Q)����bgm��+�1����`��F�py��$���Z��C�����`N��rɵb�߽Zm�ɻ��� �݈������<�V����렻:��Hl��K��c����������mǷi�	j�z	_'�� !/V�ff��#�s��eQ�'���l�F~�,[M�1������1�(�(�G�f~)Ga��Z�XP]���l/���4 �ȃrTUI��������!g�&��]rs�X�ҌlrA�Μ�L�h�n�U�o���i�"~���Muw��5a�&��QN�h�^����1R�V#�����/���������������˦�N�:P�w7��<�B��+�M��c$�+���M��������Y�­���#ަ�)J���4�H� �d�O�P�V:*3����� �$V���}Ē7S� (��#Y��W�ɽzS�*�s�������`%���k�Tj�!�5��Z*X:0����o+�s�����^��Vh�3�l�&�Ƚ�R^G���=���V�-#޲��~nf�ç�n��<��z�j�L�p)�}�0M�"�$���󆒲�RU�r���r�#`�C��9�{���h;k'���y��.�t�+MS u� ׭e� _0�&��:�$�ߦ���zF�
��uT�XCࡷ�NP.DO�3g�לR�A%�Q��e���K"�RҐ�~ɞ�3�~������i�n5|^��	�3�xI�|��>�&�1��5V���5����YBf��y�>m���c��d����:^�)λ����`�3����8�+}M5�������+b����}N|s�(/�T�w�s���Ȕ��Q3(���:�F�����2���hh���|��&����3����bH�PbWU�D2ヤ�a%�
��6%�;�Ec�^�k��ǡ���G����W�����a���G�t��n�i��73�����v=Kf��'����5 �ti�i3\E�i�Z5���	F��tF�P�a�zI�oS׊�"�$��G�u%P��]�v���>���ӻ
\�����2�R�SB�����o�a��1k�nᑚNs�%{Ct�?��ǌHj��S��I�y�[�Dx(�P|Gc��I (������'6:�v���VG첀��� 7�0I�_��r��~�����l���E�'���� ��˲ܧ����a]�,['ſ~nh�?r�!���_�=[)0({��APZ	�&�����&��in�Yn��$�6�	�`r#���e.����>�)�Z���Kp�[�;D��@9�c.�ZxG���+�uE� �Ib�6'��h�|Q���z_���xQp����#��`�n���_\�@,fu�/j��IE��Ո��Mm�
Sgek��wd+_�X�� ������Y1Tz�Qc�A~R-`�1U'��
��Cy�D��QW��ǟJدhd�3rF-qS~�����6p)���xy�˿��O0I3�� ��)�\
R|e/�ѡ���b� \��������ľM�z��&o)�{WE@� &����P��'n� �-xE�jrNP�(E��t���}j�엧đi��@��?����ǣloz6��1#�ٻ?N#��`w[����"��K�_�we�E��v0西^
����в p�gs��.��@G[uIw�B�AwI�mԞ�5:J>z�;��PK:u���X'��jiR�Iq������I)��f��Q��;��Tמ��i4�mΤ�sEPs��l'B��\ڧ(�ZBKҍ���~�~��cLD��?A���u�yp�[6��Ü���Ԍ�1�{�sV�	�҈?��g��R��[�Τ��Su��.^�j�P��o����_Ҟ�I��'�R��h"�:Fz��j/ϳ�b���zߠ��X�$]�>�ˆ��~�u���y��OM���/_2) iUA����b� v�K��V�>8t.�;�e�XrZ�� ;j���f�U|���t��(�#5bJY�f��������s[��4�`ˮ�^�v�f{���%�G�X!M�� ���΁rG��S��7ᓺ��D?�G���Z�q�*R��#y�Nq�H�.	�oe�si}�A<��g}�(��<� ���X {uUY�s΄���&Sɦ.�����d`b�sW~c�$D�G�R����nN�n[2�	"g=U3�N�$�5*����f��l��D4o� ���(9��I�ɤ�kͨ�|ה���M���Գ��Ԝh�Ȟi�<O�If���mzv�jE�2YbT�+Uu���wC�*��6���9k�`�/���=kS��^�
�-�1|E)E$�O�Q(�A<�*Ydj��ȿ5@�M	�S�fH�N�{7[���?�O���ց�c?�K�\��S�B��V��}D��4g8��1���F0��#z��Ys����ޏk�K���T���[l���W.�D�|w�xk SM��`Z�$bO1#��f �*Ǚ�Z�I�锌�oQ�TQ�Ĝ��#j7�yL��M��Ò�	��:�͙K8�붥����&� 
w�����K�}t���ҥ6$Q���xt�:չ�&U�?\�	s�%c.��}�-{?6c�Yg*�������N���^��V9a��&�˨����"��^t���Q�D�kF�\^\jE�n��Z�����u
���o)��J1G֐Z\`��l�M��H4^�̰��>�v�^�����v i8Ȋ�!�"���?k��Ax>�� {M�vޓ������u �ʗA�t�;�s�wr�s�D�����R@:�CJ�?O����#��<c!$?�EPr"�R��s��}9O���3�St[@��`ةB�ݡ��!ee�W�T}Pm���%�ͦ�����.��	�A
"ɜ�8�v>�`w	b�n6-I�.`n������(v�l�*���k|}A��M��Vު��P����"4%[R.�p �`����>��[N �n�����<���m�8�M���0�ױ�����!Hݑ��<#���j"�
�K��?�8����������2.ˣ�h�����ͼ��3u�>,�,�\Q���`��o������BOBo�̥Tk�R��.n�N�/ef�+�-������"���?���'ly�&
>������H�?P�Չ��_�q�t4HE:k
�6<��v����85�=y�F]��]i	��i��\m�
�i�������1V�rn�d�U�87�i�EeY<�1��۽�����AE�t��^f�������N���U�g
p��4��_�5&�{0�mJ3�0o)ݹ�v�/<������1�c�m��;N�U�#�y}@H��6 ��.9�1}�����+��	�FU]S��y0��{��mS�ַ4 oy��h��O">��������Q��q�=B?N�[G�6N�(p�wɉL7�u�s&�0�)rQ���AY!b��ȒF�A�ۯ�Y�Ep��&���#�Sm����|�q���L�������! j��꿘B�Q,u��BŬd���A��s���<r:�N؀2x��,�U���,y&
�#�#_��]ГIVzیS�ގIZm�蒕�Nù���ʮ����84� �/J���Z�EKi�]�1�V�a7�Gk�w
�h�_�VM�� ��%)�<��� t�${f'�X�:��X!|>�V ϻ��D8E\�QA�M!vK��p�U2��}��c5�Nt�cIc���%j����o��@��az,��}���F9j2W�h�8�~�x!�x�N�wj_���h'B�M�=����
�p��G.1�\N���?���a�QԵ�}H#&��������D�1ݩٺ�i��ğX�������̐�o�oK���C���}5�.��Wj{�Vu���7䌱�"�����w(K���f�+��*�0]Y�t�(O�������>(���Ȗ�V�i�P���!2����ZV���:�� ���U&��q)u��I�G�;L�V��U���0;$2n�j���H��|5p	�zQ[��(:z���.AGN�v�,�E�?�In��Ç��t̷�疿9�u��0��D+b�������:}�M��)�o����SÙ��#�o��T���lFB!�'������Xco���,�/?�Cf��"8V�c�� ���aIx3CB���h0�L�O��]����k�-%�[�+z6�@��e��-�>�c����ȟҌ<��PH�t��j�V��j=qƱ@F}�ѿ��1TmT1Y���0r��-n�I)t@^���dǅ�}���b�Ld�<��^�x2�P:�P���#�&�+xB��f��EU����4�F3OZ�Y��pCu��v�#7�}�p�i|X�υi�9���+n�����A�y�Th�}p����ɐJ��S�x&Ƹ���HH�3F�kA�0ˑ%R��U��J��|�W�M�D;h������K ���������[rIU��1Ι��4�B�4�5�xl%�P\���+��ϋ��`�5R�mN��2���\e���̬�V�y��c������g�^UDs�^-��!<�ԡ��m���������NC�B�U��i������>��yQ���#��2򩘭������o���p��E��6�y(6�RU�͹}����U��cZ�b�VR⶜%��w����ڑ�q���t۳�7��Ϣ΢�.�nI�����4��Ŧc�w�}����	���.�Yn�ۭ��N{}���C>H��yy�� �T�l��M���i$,�eb��㌷���Oj�
���UO[�~Ŭ�Z����>G-�o�������&s�58�O�2�NSjh�~Rܭ$xdUi3�C���2����	�Wzcױ+1�@ĠLL9��z�q�T���;O����p&�wp�?�ؿ�ϣ�c�k�3���aDZ�cnb��l����������e���^-�`��T��x��GKL��K˸�+��׻���tD0��J�����O�wh��R�I~ב��`Y�%�T{�t���ꕾ��<��)�,�[̓��?O��.�(�*�n�Zhj����5x�JI���Z
����,0-D��Jm2
�X
I��/"(���w�_�(V�=�� �+��^�
��y������������`qX?��㗘��@�'M�ʇ^���$t;j��5�-����[6�%���(
�-3� ��-�"���9������#�{E��v�u����ϬLzظg�\%̙d5g6OL�5�E&�KKpZT�]�4���}�`�7���)m�@K�[�9a�2'�!���p��ԾY���<_�Se�5�,Ѯ�lCZϝzjn��ޞ�ϸM�����㭳o^�+F�ܗ:w@�L/�&sz�
C�	�P��i�D	��7�����`�����B'p�ϒ���,yrC�E����p�(6��}���-�l������4ݩ�F��>���N�v�hd�����ͱ�����i����H���O�zmIF�~�l��m�S+�^u��W[�U2A�?$��fC����{�P�_;����cI۝fV�N,�9/PB��
�'x���bEE��o����(:E�[3q*�4f�1���$�?���gv&|���h���h�D��uʠ���ޭ�7���F��~��@m֪
~�H׼b�ސ�D��]��˕ G��Y*���/s!����L��9./��k������׋���5DK�n�(l]�I�-�B�dl\	X����J�����t�|�Ȱ�W���=@���Udب��4'V�ڷ�~V���#W��_>����>�a�+��?�;����B�+CH�Y�Vn�N�f-�mc\�f���gM�&�u��kG!�!���I�M3ģ����{�� ��/�7��<R�utQ�v��f�^�?��p$�V�[	`1�g0!���nn����]�ON��ґ��]�.��&��������wtߐP�3(�F�&FߪhP#�<���1
6����^G9�?��T�Q�����������<�PM 9�Dt��%����b�;)Q��=�^yɈ���7�$+�u�p�Ԝ��6�����~�OI	����Z�Dͦ����l<���%��.�2l�:���Z�s�{�~U*�J4x���_-�<�:���a�
.?�N逌��Ը�٥��\�*Po���
砪?�Y�ҍQ�9��@n��z�Q�(*w�A��so�6h��rR��5} d�,�� �M�P�&��$('��}��*���W�'[��/�`HZ��"��2�?�a����X�����y3��y�ޗ��F�P��[��#Ͳ�y��ݪ}zs��F��}Y1��ȃ�B&v�g��5"����0����9-���A|1\��x�v#E�UT�£�ϴAǺ��΢Xb%Z�i�i�.��tZ����z^": �B�8�ƺ���i4��/Ȱ4��K�H�92��G�3�4�R�_�>T,{K�by4u���#��3����=4!���WR���R����_' �c�T�;6�פN���$�<>6��⸖&_̬2X�,��>�>�V��J�mt)�Ģ5��*li,���y`�/� I`Ai����p�u-��V4@��Ro�x7q���a ㌲5G��W��+.�n�yDx��S[��j'0+1?x3P����_ 03��w�]F=���A��e�_�z��Yw�D�p�wG�rF�m'}O�������8&��FԳ��tݵ]->ik�����e��̂�A���8*@�Ve�W������X;��\�!���/Q� ��;k���S�(�*�sN)�h���q��9(�j@��3�J�U���`��|1$��^8Op�*}�l��"�4䬡.f�aE�.>����)��}��ʠ����O��Ql��� &��ev��{U���sc+��g��6�S�m�pI�b�����e��i��{U`R�ױԛ
|�D���ro�g ���?�O*��g��߹�f;�o}p�8La|�ܚ>(��qH�3y�A�)�w'	��P5'���-��N�C��,G����a��a�_�h�C�wJ�
+7<�|��'�Z����:[Iѓ��T��m�1o'��^�sC����\�KՈo�S@ݾ�/�����hR��V�U���Cvn1w��W���n��<{q���泈��?R�h�w0vp�7���ܕ3e�嘤�۾�W���}��dfK�7}�Ǎ�����0~ĄZ5q�^�|gs\�M�ݽ�����ls�a��I�y1���m۪)l��n1�l���J��)�0Ɓ�5�D�y��=@ �a����|E�ߔ�Z)(6��/�vX�`��f�������k�9Fi
����66a�2#c�"��J�,�� EtQE&B��y�Eko�~.f<�RC�D��PK@Ct	�W�;1�L?4]R��>�๕��e�*���0q���hj�� �e�ap��OQ���(�^�ݕ�H��cF݃ҝ#��ףTC\Y��f�>�W��|����(>͔�kN���}x�|I��a��!���ʗ�����@kJ���:��4��j9�!�QY��&Y��x�8l�$ +�C�}�D��F�̸S�[�����G~b� ��� rH���G�����+V̸�ҞUk�mɮ��*ٍ;C����ԥ(��n�,����;�}g a�(��[FH���͞�,���d�}��K����;>���'��m���o��%Ŭ1�u[����r��^tm��_#��	�T-�ӌ�i�2�L�f��E#@0&�U�Y]�I����n���u8����ߎḈo�F�*�����rN�uN~�̛���I���_1��+m�E�X(ć��������M��-0C��@�@��'3Qy���i)�|����	�O+J��ʏ��wO��4��z�%�n���z�nwΦ�����g���y�����5��Ix�Ǭ��\�>�y�M"��O���sg�Rw�]AX`~6AJ޵>����s��	�@��/���X,��y�RDq3&�����]"P�� �� t\��\u�4��LΥ�AO��c6V�](L��&[Zq��U엛�.,� �}������z]T<��D�/ck�o���)_ g�?����c|�:�;���U~�}
/��er���ĵz���k�s��M砞K'=�'G�f�w��FU�.J��\�8�wf�oI�U�B�
y�]��S�p?Vq��ڒ9X�r�G��2�� �k8^��1��nQŝ��cB�T>]�v��'����	��1n��2k���-̱�T�N��Y���ȊW�HI� �AfR��!�2I*	�+��J�̈́�ɣH��0�G��1wH��qK�������r�_�~V��_�X�8)�Ozh7�y��Y���n��IK�[�<ydY���s~V��w�Ц�e��Ge��R�Y� �+©[�	_�ܨ�����bnG4oof,�>�a}���(�Üh`�o[0Jb�D�	� �b�*�Q���kn�G�B8<$;�ʸVk������F��a��Y��Q��2qD8M��3!m��x$�C��r���j�s[���(귢
,09G��p�l��\3�����Qb�?�l�x���Ki�2�aw�5�o��&lB�N6"�⻤��[QZ����]��}��w�cV��������� ����_�zy�1A��*�C��5hF�G��Ɋp(XY�3`�itS��!����ti[w�@
�$h�g���ԕ���[��h.^=����q��L����CjP;V ��+z��B݅�'�9
K�V���rw4�t����i�&N�B박uYh�Ŭ[�:!����x��U�s��B��:/�e��^�Ȟ�m T�&������0c�I/@^6Gj��c�Z�m�`鋦4A��#�Č�t�aE6��[�=B��?�'$6�3v������K�ț��YvL<{�$ �6PF�<R�%n	���T3
��.��g�XL�[t�gu����In�E�S����.�����@'�]c���fjf�n�}s`nԌ�P�Ģ�A���9������S\�;L4��<�Ɩ\�c����V�b��[c��� �ȷ^�H��]���rr_1��T��/S8p#w����P$ RfN*WX�b�J����#_�k@uה���U�m�{ШAf�0�"��c���j�Ъ?C1 m�c��['o���6�6�=��w����t�ԋ�n�2�H��Y��������������GbT�A�F	��
G�2N8����(e8��C#��_&�	�t'LV;g2� $�Y��=�Jwl��;�n����	x��7��O;�ugn�g>�]"�"g�8��� ��1����v�4���k@p&�G�6)�Z#$%[�=����>2�$��1<�*��w"A�M��פ>o�6��5ά��"��vY\3��aj���i2ĘR��?�ڇ�t\q�p��-q�J^�r�0)Pm'���e�݇�3D��\�/���其nR�L�~�G.^� ������Gcc�-߶{�[r���6�߮V��7̵| �����É���X$�:�
�-����{<%�2�0�:CV� ����0Æ�;���5?8��
�t�ԛ�h �\ƣ5~x�
��R�Kx*Sep��~�Mj��������X�-�/�K��^5"o�S Pv��اu��J_�v�B6k��|�@��&.=�����Ac�>�2�����G��!2��(�������=��@�WG���J��w����W%��d��4T�	5��ހ��$����9IiG"'@ۆ��M%N'#�������S��m,a	%Sh+F�����)$��*��	���/_V���?h��MH"j��u����_[�n�\l�"����-��<C���j�ۛ��������c��?�h�$�	pb��y
��'��A4�2���� �լ�\��`>v%����f�S��T�������y>2)f��L�f�\=��М�}��X:�S�0P�R|����i�B>Pe��~|I��пi�scI=�tA�)Z��_����C�6I�A�l]�f�ۚ����Xۓyا��O��K�	�l�0�f�~���^X$Ay�'����A��0�4)���$d���?ß�d=��h�x��z �N������s�]��H�?��o�� 5/�<*`zт{�Ȯ� 2R@����`��	�a�SR�&k��u'w�$N���d�̀����h��{gڷ�Ⱥr1[�Ņ=� �fB�)ҚG�=�����n���/R� ������?����G�7G���ݷ���'�R ���ivL^F�k��3��@�B���h7�9�4U7u�N�#���_˭�	�4��0�A�\�8?捆dg�R/1.�	D�y�;������tc<Y1D�;��K����̠�]y�������i�{�Ȏ�+,��IUe��E
�{Wo��o��/�z~��US�|�C'MJ@�	@rp�fh�b�Y{񇮝�UR n��t�-�PS��!Ѝ�I�!gi�R���0��?�����oDņL�f�%�;}�]i��z��	�h	����Wت�Q��gi�|��e"�Z}�:�0V��G�@�����[��H�BY��}C�=r����4���	?ru+�a^D	��%>Ewwv�yEd�Z4�� p��X.��Թ)��^L�֪�t�u�Xl�C#U��S3�Y/s,xU�c���N �+7E�z�D������䱙.�h��+��"ܒ��	��/N�f�ڡ.��1�@�ؘ|W���	Y�Y �V�=
-�̅� ��w�0=!�Ԃc7 �"�����C��8�r�"��l�@R��l Ĩ�h. ���V�{������
�^5w�&z�����vG{��3�5 ��G�+,�u��ݚ��eF8�7��o�E� ���.=����-+k'Ym\�v�K2-n�U?�_�t,�"�c�wl\w�8�	��w��ވO�?ga�C�h\tbb�\��yx�>���w܎�)��j�<��Tx���Z)	N��L��lY\�q�͙7vx�y"j���� 1��D�[A���&Q*s�	[�'�(%�SD9x��ڀ�Sޑ7O�?��z�����ګ��fA9P޿b�Jls=�9"1�����0m f/�2���N�utW�T�@���PcFW�-��AV�)oL��7�	���0�L?�]���7�A���ʯ�#���A���)�x����Ց�e��Z=�w��-�ku�� l�ɱ02�(�'�+A�|�o����÷�2:��Ai?{������1�26�k|���{����"X8k�#Wj��^b����I������=Y$6]�<�t�
xN�s~.��؋�-�&H\1��FVɀ�@��6;����j�#J�5�?�Dۨ�
��tG�sl(�Kh	��h�%v���h�V��u��k��9gA�W�	�:�*����dh���CNY=`�0��"�}�fc��y&i�s�e+<�
�я��豬���jt����fuT��W����yU��.P���'�&y��>6�m1'��C0r��+�@��^p��/��'�4k,|�� �h�0(+B����� U�`%�����tpP\��F�z�&���i�d�[����`%a6��k�8ҐH@r��o�Cֲj�P���h۪��y��ʢ�A\s��2;�&_~���GN[�jk����o�`��s@�hA6����M��#�ex\b�|���C~-�^�@��鄭� `��^]KK�=�[q|�H�9�i�͚��VaV�s+߫�O���&�������&��/� �Q|��ު�6�EB�"��"���W�����q}����K,׋��L�dJ՝Y�(/"�PZ�����Ϸ�v
fz.٥����ݣU����e���8��c�A^���)�1��kEG��ɶ �	�����[�+UD��l�eB� ��7e�=�H��ߜ"`��K�R)3�{�����$=z��'��=���>�ca��.꠶&��⧙J��S%�pys�i�����p�^����*y��S���1�%e�M"�0J��h�K}���Bx����|��.R�,��"�W��{r~�o��?�Ƀ�8�	��`�6+�R��!�I.����ba*�����Ps�z�@���AZ�R�{�R[��<J��
{��z�-�5��;c8���w���&B�;��w����ѱ;���겏�w����g�Pp�I�7��t>.aG�2�/�e_�����
-)�H4�-�:�R3N�iqV��3��U�Q^@�a")�r>�/�c�!Y	s��˃|=6"m�&ی�� ��� ���
���$\vs�||ϫ ��j�vg4�cQ�kq6�w���V��"�ěp��mS��Y�o[�\�j�)"o,�fb�4�h�͢�� ����������]�9�q�5���_L����h�)�g~{(�r���4��e��g�k�~쥂*�����GF��Y���H=����@L�G$i��hl�TH9P��	�	R��S��
�-/I%<����v��ȸ<X�\Mg��.���oF�v�t%\���ё}��%?��Gu���yB��!C�V���[NoV�mv/����L,dw�C1V$h);�c$�*E�qa�t�2[�Ųl�`����>h����ޙ���wE	�����S�O��~�nM���9��+:��{������Nav	�Xp1�6bU&t�hq]�>9�g�pQK�}�TkҋC΋��F�7P%���}�D\�Eϴ�Ri0��~R����F<�`�Y�t�
P��ֈ�P�MN�u�x�8!s}M�>@��<��-߅��?�]�����!�I�mh���$M����Uؠ(?�@�q�q��ÙL)�Z�Y����+S�)]K�p�KIyR-����eC���N�^M��G�\��4fcQp���[>�&�Ը=J����b�����
kN���� ���!��c
N#��W� �48�����銔��+�0�|�q����-CV"c�T�3^�WW<����ƾ�q���\4�jT���-����r�!ٟYj��i�H���I�q�5G����2X� ��g<�ˈ#�{Z� �[�ͯ��#[>
T|}�vYo� ���>�b5M
����*�D�,!OHHL�c97�u�3�V*,�~ l�<��;{���pb�R�Շ��:��1%�-0IUV�j��m��B��U��{j �G�b�L�r������ǿh��Tsgm�8U�3����"J��"4/A�.�/,T2��1�Q.�IL.��z0�Z�M��}5i�ͽ�T�Q�F�I�9w�*y&�n��O���K�첋K�N=h���)%�1�e�����=I��H��7�怗{�7s�tŬ�0F��,-����W�y|9�7��������w���BRu��������#(e���"�$��E�g�"�� 2D�#�aKA�È�aC4n�,�)?(v����j���!�DֻR��[��|��C	�-e2����\Q��`eܥfo��N����X��Y� @��_o�e�qg���U#`	���!�s$�-�ck�f�ʯ2R���.�{3>�����k��
"�+�	�^�p���5`̦�U�%��H$5��1|sA��nX������鏥kֻ^�{"	�&\�4Y��կ�p�ﴎ*5%��3�Q�]�o �qc�G��w�d��Գ��G�v�c�nC�ˀ��$�n�����'���I�\M������B���kuED�3�>m�/��_t��[��^��!b�=*�5x��p7�o�Ane��a��:x\?3���W��0��Fz2���R���X�SI�x�6O�� H3���$�b�uyd�
M];���Gf����#��5��
��g�O���!3?;���x�P���բ�/?Ǧ/���u�B�H��PPv+&�++�[w��\�2*��&ȶ�k�I
s��ENi��?0K��\� �be�͞�Y�(
آ��/(�XM&�s����r��^TI���ѷ��)>���(N�~9��KG�˝�F��!~�ա1a�����!�e���m�}"vV��?�"�v�������<�MFU6]%.���e.N`�+VPj
A�U���м�f�.$����ʊYw����W�r���X��`"t��Ŝ���h�OO��!F;6B�S|�6 �\
4�+'�W{^ݞ�0v}�X)�o+���8�B�^�w ~UX�oT�.CZO��O#
p��Ovي2��
�mǿ�$3��y/�hl���O�y|�|��%�?ZD^���Cd�X�FA@����po-����D�����κ[��X��6e� ���녢b�Z�g��y��c��+^�+r��\��u�@���r�#��S�f��f%�K����Ӂe�a��GC/������1�~
c���2�l�;&˓u̬�����"rj�V�-W����M�cVu��+�W� ���G��!P�md8k]�c/�WLP�4~�g�/a��0s���� 7a�Jo�E<!�W~�wgp�h`h�<���{net�Sf;c�=|7`�T~���a�+����x��/�+4O�2d�Cޟ�5��hv��Ͱ�r}9E�@{\|d>ة�ݑ��*�6u��:�ʼz7����&��:����0�뱿Q)I��њ�4*�j���*���ToG ���W=�_���غ6����eJY��8��6�k	k���	~�.�H�	HG�+�[�b1��[�i��a߽���wV��6#0j��V�;�لp���:9�4᧽ۨ��+��G�wI����I�� T�0@���|[����:����Ǧ���BKB	�O2V���Oe�$��X�R2�B���f��Z$1��%l���;�5s;��`ב��Hu�a@v�����Η��@
4ן��o�-��  �&��
p�͍ѵ��Mv����S����5�-^��A}@�e�@+�h�~�	�NūWP�������.Z�艹4%
��p;��H��`�kg�/�űjQI�EX���,��CT#�*���g�=�����N�W�����d��������'T)g�BBo:�KFW)�UK6L&�� ��s���el�A����5s� ��NSAHj��;mt�1�'��=w�OR��ԅ󎯩"�U	��UB��s'�S������R߻vQ��bx��^1{o�	��i�A?����ۨ�r����.�,�]I��5�>���Y�Վd�i�Q���AU���AK���Aמ�����,R�Gt�m��"a@�]�$�ߖ�G;�V�I�ؚ�q���6T@ĥ����n��Yo��[n���>�ǫ�ﳷ��ҳl��Ƿ��z�a�����,4l�:B.�f'b&�����'SI�,�[���8���"�b+2���A$�����'�ա\��4.�Tđ#u��W������܁��g�;,��"myH�)̓�y8r��D�z�9k��U��X���t��K���j\9(B�����8z��=�8�.uK6��1����|֖����"�U��,�����؃^�0��ժge�*��d#�ꓙ���#�GN�{�ԭ �)	ac�� w���l�pl���\�@�C�d�+�����欦@E]�y��_����DB�)b	�CƵ����AeU>ۆ"�c����=.��w�&6��\�k����i�?۟D�
��i%/}�/(S��*��Y�|i���r�R�/)�nIx����p�����̋皁 �p��B4f�����_���hS@�����9"k����h��[�`�U�m{\�G��[di�b#*t�+j��R�1v�j���`�⃧��Ӑ���f,�܉}PO��Y9л��w9�<�eJ�|z��NG>Z	�����X���-��&�� ��� �^?5�"�CM�d�z$�f��U�2:����,����6���%���=��qˑg���&;����j0�wҿ%����@_��AZI�D���8K����)�Y��O"������J`Hj�P�,�(j���� �b�J�7⟆F���ƣ13i�G?�#�o_�oX����82~?��P��:M?GPAyBS�.���f�����4�O�3�Y&޽v|�����dP%r�b�9�d�I�m�Nk�q7X�AV3�=����Cu�i���J��w�кL���ș��7c���Fǚ�E�����:��ն>�!a�D0�:�`��T�ӥ�L�K�[Qd��-~x�J��<)������]6�=�#�-*,�w��[v�A.}Σ�i3�]xb���Ș�d�32�I�����A7Z���N����R���JeT��	�'���T��_�($�C��BN�ii^��|�+���j�uѭ���'�Ua���Fġ����_6m��K��{�F|�G���I�ꑨ�����>�g��S���R,���|7st,�!�&F( rꗄŝ��-7�����pk�:�����pF#�@�K�s>Ϝ��.c�{�ѷ!e4bUj1�6X��>�*/�
�.����I��� i_*^�w�nx��Y,�}��^w��Z9G������}Y�l+��5�Ȯ��J�miX�gD�L��"rɤ�*jz�Mh�[�L蕊�Y^�I��=@��6u�w����y�e�WRgԟ�6�5�V�����N�<y�r�av$�Cֺ�Y�n�٦IfʼVK����S[�l���0���"|`����$�F�Gǜcg��h]*�{A1�JJ�)I6�	��̆�"ꑛ�y}���(�XV���ow� uG���O<B��fz�E�0FtJ#}<>�x?��)M%z>K��k�;;��n.b��ᆶH�!��~S^�����)g��c��_.D#0a�1�A|�Ϋ���'k*����C���}��3��7u!��(��<����P4�	so�%�+����/ײ$\J1���c����pE2�rJ3�;���3�P�����g~�`���ֱ�u�������qv(���d��T
t�̴�C����f��G��A�NH�cS�},�)s��M6J�Y9;�Bsz���^��A��(~�L�^Vm��*z���yؓ�ôt���vL�A\�8S�CS��K�wO j�o���q��Z���wBa"3	G�'�.7�������e��lU휳`����v�J�����"�-lʹ0䄉��},T���#(`G�x����0���d&�]Fx!�8Txi�v	5y_I�s�q�����ܙv��?$ !�C��m�o����������R:���h���Af��_Seh�+���S��"���g����껣b�ΒwCڣ�XU1�~r�I�s5�'Vtt8H��"@R�%U*�j�сV���`�*[?���\�
���Cl#p���V��"x�P��r�%�������j�E &u	��p����[P���#dϸ�/I)�`ŧ���C���t ^*�a�Ӵ%i�hn-#�آ��֭{d�HQ��V/{Bܹ��w����2G,�>������>��);�\�Z�Mi�*C(�A3�'㌯��W=
��3]�O�J�^��0O�0��mX���U��srg>�Go�Dφl�M>#r�xIST`	j����O�|�f�6�?�����TBˆ�j(�<n�)�J�/B�Bzc�{�P_z��iD��D
�A��!�\.j��]�\Im\���^V%]�<��s���y{�4��8�I ��*�0[�0����&}��"�f/��;ȗ�� �q��>�����"E�_}'�PN�Yi�9ڧ�*11j;��U�	5�E��\_D�#�`Q]����g�1�lc�de�6%��?�յ���������Vs�d]шd��*� ����Q����m�>�,A�y	�s�@�9�>�G��l��Yvh��l ��\Er��o+Fł����!�q��T�&��-Fz��,}x�^P86OR��TJ�\O�lb��]J��u��3V����5Q�fĴm"���`iSɉ��}$�8q�2���^s�;>��P\2��b)�GMcq[{��0����	��G{��=�#A�����D����hӵ^�7�����X��j�\��-v���|�F������n����o�<�PӜY���|�_��W)?����<��qW+�Џppk�GR[��|��wq��P�լ��XZ�k>�K_q�p�ǺcV���υ[�Φ��P��ʲ6tɭ��I�J��@�����`Q�8�b���&�b6vY���E�<Wϧ�U�8�U/$�Wo� Y���
˭{?��n�W+�Fہ��� R��}(վsܱT�3�m��	�n>������4���P`-�����h����k�^6�\��}^��|�7;"+ڜ
�<"V�/;^!u��m]�W��`K��+�O� d ��!h�_O��MN�v5�F2��DdI���'����9���g���E�����h0����d������0j+�R=q$O[PF|��V�~��r�-;��L��`�M�*��Z}bfЃ3gE� �dO����
��J�Z9nBdgdL���1��Ȃ�K�y9Q[)�+���3P2�A��`��h����f�F�������̲�F[�sHd%�M#G��{���,���k��'أ�*?G�7�E#9�}7JtxʑU�C����>����3���]a�?�S\��`��_n!4$Λ�z�:>J��1X{ E�>�VvW6c�*(���y��;�w�ɖ�p��id`�>3��:�^�S4��H����&�v��݄��?����*����$�`�+IxҠ�\7`���8醞�w}����k
��X}����l��M�i;���d�cH�����ଧ��,>������<~"d7�"��}x���Q�+��Y��LBO���9P��i�������_�7�bD��hKIU_u�U|����|&�9�̺�-Ն��T��O���sum�ኺ���v��y�q;��U�>!**����?W>�R�-��׳���z�ϙ���
9�J�ޭ�F)�;Y����=�y�.�������n`B�U�~�	۠<�	־.N�r�����"����jMFٹT�@��_b��As�xP�6�ke�3e�A]Ћ��hAKy+e�"���_dY��&��Ƥ����b_��~$���[��v-,!}�K�2S�5�-?�y9�0��%^�ݤ"�Ƌ�-�kk�}.t�^��f�j�q"�*�u��ȕe��R]��Eد(m�9����_�������ζݍ��2�t��4$�r�N��Ux� �8�x��!DP�P�u��Mŀ�gj��9v�qH[PF�f4@g���jC�ڮ��35�<��1:�#?~d�K�}1�ޜ�𭣪�Z�_�0j�a�z$��|��>�Ԥ48��)d�_��e��pd�%G�F�S�:��_���J7#�BV��j��mݞ]���;wL�la'貝��D��6V�2l����0��4�<��O�g�E^Cݖ����������)*z<���(h->c���� 4%������cA4����kC�f���¬��n���&���M����ߌ�45��;���4;�R$�{r�N�<L�v�(�b�w����K=�^Ud�8�u������?���6����p�R���l�ھ�]}(ddrZ�X���n����Z�����):m��q;Ծq�60�_ �di��o��%��7j�PI�_���o�Vg�N�^A��8����}���Eߝ�0蠤�ب��6`3]u,;��0�m���Ȑ��8L1�δ��!ю2���ZK�O�
]5�&M�L�=nl_p�q��i��}�o"rN !�(L��1����
�g�l�~���2;Lz����>!Z��j<;��LKަٌ�9�r�y)�T߹À�<#��OD�)𤔕�"�S]t�CoR׎6,�B��t�ٿ�M�3L���2�+��d�.�7�[���Dv�0Նd�-O����plI8�Eެx�,j��ɩ�J0��&8�r�4T�Wm�WJ!�#�_����.[����SZ���na���ܰ&��"�an
�%>����ĕ���A�*���h�`⽻Ζ�x���fjo��{�HyB�r�ϲ��8n���*m'6��w2��;�vŅ�$�A�#Ikqesլ���o���z���At�p���Z��~G�_���������H�	��w���(������<�"��-��#��a�f��ڱҽ�7�`_L1�k��d#�u�F���k)� f�5��E��v
������/ރO�o��d{��+T�|Kdd���\�9��G`S%�Z���bw�F��~�Z(��oA移+/8�٫4[� l����{Go]$�ϐd�D�P|����]�|� 8R\��D_����D'Ge��#w��T�� s�NQ��͵�����I �&B|�C��/�0��캔қ�e�Ɔ���?O���e�6{y/��@�w�or���HL=Z��X��7������C[n�R³n?4��6�H_߮�=#�P�����F�R��1J|=��36��5%���ȍ�`�'�cmR��'8�1|������br?V���n�J�R���~H�UO����0��5��̸�����ւK�JU:l�(Y�������	~;����[�����>�h�TX�7斓l۞B �*�Eh�r� u������E�C�4؀`��6Q�P��̓���kp}U��[
��k�����a�����̜��=��s̷ewA��{Ό���,�U~-���{L���T<i�A�Bx��ul��'0 Hz�M4�;V�9��6	(�
-�H�����	5�r���A��F���`�i=4G"ǃ��w^�$P���!��kZ>"��I���J!R���ވ���h���.j���5v�Tƽ�[�B�6�?&|aE��=+�!W*�ȭs��������{=�,��o��4)x
����]���|ܢ��7�w��A���E����!ݾ��~����M��xha?D�ou�L��p0*���	��s|
;\4y�T��L���isM�ߔ�mK�+�լ��s<�n�U�U��宙�!��d�d��)����m��'%�민���T���Z���;�ܷ��5�pӸ%�b7��9��.T&/7�Rq�ώ�Ȝ��c�a�"8���� g9bڲ��>�Z�STh-��tni�.X�fr��@��!HYCS����w3c��:H�B�K������A�^��8��AQ��
���f
��Q7*L���_w��a�bkř�Ѣ�����������(��JV�8OQ����|D�}S�5;��3.��HQ���ٜ�"�<�;�2(td�.���p_�{�*�e=�c������x�h�q���3l^+o�Lը�fN�y0�5��+�:iI��Rv�ٝ��D���C�&=F�Jb	c�-U�
N�o�e�����_���w����Ȇ��j/��ip	s�%=�O|1@�y0M�;$wy�c ������h�P·@L��ӡv�#Ŷ�窭-DLzһL	,��%���24L�ѥ;�C�?���o3�eRۅy���0ɢJu��f�+~�!g�U��D�#�,��vV��%O�#��6���?5�2Ȗ�;ʆ�-�ԏ�4٢Z�wr��|#�����a��pK6�K��p�����?��
6�+���}
�G��Q�ӭ�:��yb��6$,�����,�"W��Tv�۹�����iv�㺑����i\�����M���O�=RJ\j��f��X�����g�<���NZ���E�~��~y(L+L"#���2.i�����J���)��-�^�Q�VB��;����xȫ�$���j��R��<�������:����<��L<-�ň�@O�P��ӥuV�]�V��@QK�h:p1&�yuuєɎ�ݱe^:�{I�8[#o�Jd��o�������DJ������9�ߋ�-���(�uc���M�d���=�^b3v���'��C�q]�c��
"����fO�T��}�눐�MW�L�|�3G����t�,�Y�`�B���jA}�>�"�ou��nE�\���6��(��fM�()�������ͪw!AK�v��C�q �O�.���ip�(����$�܆d�#��w0�/ۀ�#��t�b\�8H�X.���1�f������^J�+,˘� ?��-+ �((�u��G�&-q�QnE���~lO��;���0\�4���8ݣ���&h��P��؞b���W�o�M+�_���D�[j�2��)�m:����k��k��zGN1�~2Q��γC�0$r]8LqM2�:sK
���5`��jP�@�ðvL:%���J;�U%7o��%X�/�A��Tx"�bnz��c�
����z��~�t#my�HC���X�|T��O�$6�˾�T��g��;�� ��&�\��LLq�cd^}ҤR����t�* ��H,�ح�Ż*�!������q�ފ��Gљ�f�["�s ��|��ͦk?�{�%��g�#c��P�)Ch{���w�s@��/�e�em	����s�܆�BUZ�pD-]z�	�l�n+��UU�3c[�<�<�`!�SG-^O"����j�^��h
Y� .`H�M0����9wgs$y|7J~ 4�����}����7V�-�gN�����>%�� �m�ն�X�b]�Y���_j%�+V��MyN�[�l[��_���c�	9$��r*GF3#Ԃ/��Rm^�/ �~)��X��� �E�:�G"�L|J�m���͹a.�`/a��B�|�E�:����������Zf{G0�c`��{��jV0©���k�(�n�J�M�a��!��T�=ɋ�q��5j�z��V��a��ӵR�ߘ���-;=JWta,���
��J��)*��M����|��Q���g}�W�Y|�"�������̗YE�:W���n�*J��/#��K�Vevq����
�kFd���~����Yϼ2 ���N�B�����ҁƝ��W&��fJs1ut|fȣ}y5���M�N�[s3cg?�8u��z��D�x�:뷑���(K��e�F�z����<�Y@�1A(��x$.p���'��??B��WGul���=}�JQ��dx)nDd�f�B\qy�9��RՃ��g�}	HA*�����h�:��5���ǝҨ~��gi3m�^�h&q<��7�3����N��7Y��~�ކ̙c'.
.�zJ��+4���.�H�Q�kiO(�19 *�h�~8�b���1�D/F��j-����a��q
%����=�o~��~�ٹе���J������#����$.xY
��q�E=���p  H�Ǒ�����ʡ�����W������$e����������02��v��*��GY�pb&�*y:���G������Bv�m��Wrϟ���b�p�d�#����BSh�`=!���2�O�|�����ON��RwUV�>"*ѱ`��Ydf��+��gыV�+�3\��Ƴy�������樍?1���b{8�tz����O6OI�x�R��Vk�ö�S�sdaQt��Dat~I�%��K��@ͼH�&�Y�3�������ژ[������ƚ]g��kEZ��O*܇�;N��B�4��ї�H"��6�F�Y2J�!M�?�G��J��4e<U�������A�={7�&߻6�ټ䤬L�z�t����(Y�{k�ŀ�پ�t�*��
�è��*�L*�h��7� ;�cw��(�&[�c�\��9e�uЂx�ma e4U+������Ϛ�����q��i�^������#���]�[!�����jRE2ŇFl{)��S��c��Ϊ8$�;�KMOF��06`t�����|[�eiT��;��H�g��|����f��J���r� ���$La>3j����㗫�Pa��ȱ�b��
;3��(?Hrwh�Q�]B�]c�f͵~�M��j|w�Ȱ�N���CY"�J��hA\�j�>J߶fᕲ���2��吼�a��c@Kh\�O��c��Y�tЃ�����(�rR�:���G�h����t��8�*�[��?��M���C?Ek�
���5��-��l3��V����%����
�r��v��t*�����'Ɋ�k�v<z���F��k����h������&%Uq���%�Į��@��I��痸'v���g���[�و��f�4�h���,�"l��ǋK�=�.h��	������#���p<[�g�j�r�b��ֶջ��8#\D���MD��.�_��8��Y\�A0p��)��E��[��$�H�+z9{^˫�є?c�	┍-b9�&~�i�9��s�%�.�a�W��A�V��i�]�*�'0�������[���j��<��ϣ�G^�_��Z��E���h�^��ۡ]��#����6�g���m3*HY�
���+k��lJĒ|;���b��T��x>�����N:�d�����b�ԭN}����ȫl�,�f���q��RL���+Ô\���%.�4�6�7I��r"
� '@����g�n��?��D�pWY2fī	�jot'F�����$|�vDM2R�D)g-�N�۸���	�z�!p�2���eƝ�@� .���
���E�Җ��n���
�#P�>(#����+b�ϛ��"�IlI��v{��#��jӆm>���-\��K�v���ژ�>u����ܖoY�ݩw�My#�_6�����JC�y&�*���}�����Ƅ�5���R>ɱ9��t{��r��2�G߱Ro�<��?�������>�kȊ�����|�K�z�+����h��Y���rCI5����-M����;T� D�����A+ܩ*uO�S�rbU�� |�.��
�W���]>3���P�y�YF�UZZV��������h�p}�#�U��_4bt�n�������Q�)�+��֬w��j�"�)9b���RA�oJ�O�fp�?3.��m���QH9Pĺ�;���H�|GI[�N�-@���ϑ�%�Cof�����S�w����-6l(n�%�]�M�����cG������,�cDt����c$e>�d~��Q,�q�奅��yB%��d���4꩏�J^��������ߎ���/WX����h2mY���P��{�9�k��I�C�âT��7���2�#u�3���%GEժ��ǍCy6B��i�J%��Q4�s�h��D:�D�`��E�P/�ʌ�O�U:�"r$��O��5 \��'.�C�m�{!����2��l�NL�%%|<��8J�m�0Ԗ1U�(;/��Ps��$f|�(F%~Te���Jy���U%�k�.^��ć@;��L�)���.�\����M~���-+��P��@�yg�_((Ru/����#߲�����?�W�2�8�IOO�_2��	8���C�f�ЅV�����޺�K�h���m���͂!���Ba��;6~:�Ϝ�jɿfs������A���#��wZ����>֎��W��-z]�z�8�f���1N�Ûr�����OM��ن��fYbo��1~�7s�Φ>�vQ���i����@W�<a�|.7�e�[����p��ԏ@�p�H�B���p-��|��h;�0l��������6"�ilv*�7:(P.鞦O����ߖ};�Ğ�W�7fFAx�[w��[8T���}^�)X���0�]nNKi2GN[��q�nA��ט�R��T�|�$-�x��6�zU�od;��{��G	��o��I�NB��U���A�s��m��0c��!	��̈́�l���i�A�6��!V��>i��&�{x��'etu��%�i�����zj��C�CY��{elO��t��eh�d�p�6ӥ�,)^�h���'�0|�J�
~�4��*�;.��d���� ֲ��]�ϱ�C���H#f9��'�/; %�U������tX�`&K��:-+�LĿvɫfIb�Os�̸Z_�'6=H�'������C��&��sB�\�S��t6\ISߔb\�e�a���F�ߜ�*}Dq!�}=Ǫ2�'v*��o�|��H�+�͝�RZ�T�����`-�I����'Ωg{�b�0V$�wZ�p3��	�����]"Cs�@�N�o�T��g6�����(��lW��������?Ū=j?��&P��%kmF�� I�%���8w5)f
z%��5u��PB'wěj�����@%h=a>m�1��^,��%Z�@8ٜ"�sh7��ГmU"n����d�� )��_�\7�A�iSL��[O������3I���xf���4�ʸ��.�>���J���;�g#�Tԛ��?}���Y��i�0y��Kw4�ی��@��S"؀�g70� ?��0\j�P���uf�2V���:�F��R��	�3�qS���!3m���[�S���=.p�P7Qq�͕m_�(e�ٳ��C?hy����E~]������>|��U8�����4R�nq���󵥄��r�x�̊��_x�EHtA��+T�קc�4�֗'f��t7�^��9t��I�Wi!UAi�-<�O�ôk{")�
g���@�L&O^�u��~��j�'t��������*3��ͬ�,�=3��+!�I;=3��;����nM�;��E6���2iw���Z;��,S����Qg>�X�s�X�k�ɿ<s��Z@M�I.�����:h��C��`�g�*Z1�����]�~s��@���Hm�B6�f�����au�O�heK������1go[�V�\SSq� -���;�T<�Č=Y���{%���%pd�ؤ>�H|f�T��2��GT|����. ��0����>��۲�DT���P���rO�wq�lm�O�߬�#�����p�'�B�$G��#���x��_�˔<ާoOaг�GX(�sT�-�
�9���%X�7_�xD�d�q���/�_��볋�*�]�Ոf�`��{!듙&uE�A��`�jR����=�¥P)FȏZ����_r���}T�q�o-( ۿݱʦm��.�]�
Igk��Lp{�S�����|�ӢzK��w�8W��3��	"��C�_BL�Pᇵk��A�|c���o���e�ϪA�=��IJ�@�q�Vۤ�+I�R�R#�0�E6=�K|4��!����j���l���n�����:�K`��9E6h}�6���6l{����l��ǐ]qh�`_Ϳ�̥�c����wb��w�������n�������ݡ_�#�I�]p�
P��������L|�)�^�%�id��ήG���7|;�����PK��T���Z��dΥ"2:�����/��z�0��oL4Ll��4|8}T�Q�D�j0T����x2�`����2��#dO@�wC�f5�����]����00���+���.a��=i��w�V`h�zP��'��[pWp��O ]��5�n�?���J��\�>���z�=��7v�9�Z��ZF�X5#���T�&�Y�	�RY[�nk�DH�$Q�� ?�}O�?\j��:b3�����]([yV���~�,��<�<n��b�����Մ�7$��\ܑ0�OQ���4Fd���h������ш��S^N�kOz.�4b���ȸb����� �lc��Q_Ne�ʎ�`�)�6���j�a�)4�5�,�P�G:�d9��|��r�����fU�7pxOg/��� �lM1n����]��2�dz�;�[Ĝ��J����>�V>@����J�g��A���^ ���<�SҶp'*CHZm��^h��棙5B�%����<�n`�cbb�8���?���V�ԇ�F��V%�o�D܌ ��M�U�Q�S�c0�7U��3v��&~1�_s˨E���D��ǻ�gG���nȜ�~�X��7�[�rÿ�{Ot�x�ˌRx�h�gG4{!4c�Yq�!��{�T��3l4$�`Mo�)�M������;o��0�I���)�e�LeD@C��0�N�aA����xr�Jb�T��WS�Ͷ�I=
=Y�槔����F/�A��/�A-��7L�A@���m�{�-W��}�˛��r�_�"P�.�7>_ʏ�*���C�������n�	�P �`N�1��K��uV/�*FwƷ�Sk�[���#��`v,x݌5�J�7���:���z����jE��9C��&���(�ɄqH�$��8k$K>s_>,ߪ�WH�=�����XyaҤ.^
���?���{��7�U9�T�-|(ީ�9�ZO�B4	�+�Ͼ�&��R0��ƴmN��w�b�������V)c�i�eJ��7����C\�M{��j�ܕ4<p�p���zcf.�j�?�M�Z`�������ؔa�,�]O��|IZ�'���12X�^Pr�,������k6(���QS�,�P���M�o��3c��,��tCl[���P�5B߶�u�sO��3���!�T��|�h"9�C�����t@ѹ7h߳⚃��FG������=���K_���TE�`%�����~��Xy2|	z�&Ke�L���\��b�{�[],o��dR��ǹ6@��,{M�[������]�
jE�#V�Y��:)z���N���d��w~�'���:
�*������VgOB������9 ⇓U1�n����I��;,��p�/!�V��p��p_}��Ij��eY��l��r���Y���|��oQ|@�������!7W޲Fm1�	8gۢF0�1�w���{�ȩ?s%���� �A)��I�C��G�����4���Gʁ�?�8kK���b`���r���\�^���C�m�M��]�b�@63l�:�J�*eܲX./�BPd�����btu��PV�����ݰ8%+2Ȥ��9w�ƃdL95�$P@����.�Z���v�tt��l%���
-ߊy�yRt!�l ��$У7-�m���h�l�gQxq9��Z�E��YL�uD��9���V�'�-H��&�>iV��,��W�-�F�x��;_x��`�[���V���8BWe[�6�߇U���PM�,{�3r�x�o�Y��{�?��(|��(�>�3?j���7`������01V���.TN5)��0����"�W
|� mqV��2v�Dk�CīI3X�O{�-e!'k����RDz�!��ѡ�C�_`3���V��l�[������N,y��q�w���0�J�,b;�Vͧ8�3J0}g��+Y�Q�?���v}�9��5u{Ik��;��m��a��+B��ܮ �-������!>=m�0)��C'ց��\ރ���5�`��� Ҟ���)�n�~nI-~�k�Bz f��`21�������+4&�[� I��T�;m߭2�p.65c|{٧�^�VD�b���a!���(t�l'd%�+Σ�v�#.�ܤJ<۫���Œ��$��%�`�Kb��XńdI~i؏��7p,gcR�
u,R[Io�~�����颅 xZ�ٔ�>ka���ݔ�2��L���(���fsq)���w���X�j	<GT U�mٍ��/
���Y���e�Gc�m��W�vV��q.ߥ��u�����>6����8;���՛��+7ڡ.|��Ec��z�,�b�[�t�:H��K;<����=�0��j�8O���������vg?Х�u�}vM��A��-,�� �4�=�e�����rV���:-��h|��(y=QpK5�K`�m�.�OVt�{�L֦�[�+�ۮ����+SƯ����������P��hև_	�S�c>o��B^\�ĞQk��b�m6�¡��jʞ]b�<��b�� ��/�[�w�����	@\T���(�^�ޟJ0{Q�bbE��%���n_�mBZFOά*�Rv��K;������ڏ|%���B>����E�����Ǔz��,��b���oV��������J�{�t2h�.�5K��,�ۮ�����6������/�Y��%�h����7��������Oc�8)�:�pƙR��b��c}��-�B� �W�Oi�I�W�)�ҫ�W�h��M�[7)VDF��_����J�D9�.h��\�C���|is�H܉��� )$$Ybx����OQ�U��)�ofA��kZL�4YS�чq-ũ�(��7�Yy�B�$�����_d76Q.d4Tݍ$��qBI.�蟭��W�=�>Բ������#�<�aT^��;���$�EA�ƀ/M��7��w�	N�-I��=�<&<�ٗ9w�8��5O��Cv�d(tԑ��8i��B]]?�a�7�X���yMT�q���h�!=��y�9>���M9�~a���5��]p�+l�
�:����,���K6.c�Jd1�Bt�i1kS���l4;�G;�����l�De��F?\�F��/6��Oxв6��h�a6�~�XV䁐g<r6<�Mާ��_�3������Z���,d����.2����p^�b���֍�/ܞ�4	"��S�Fء�? ��	2����_���1��Y�� _�|��*='�s���8�5a��55��i���,���%2/u��<����[�ޖ��N�b�ʷ��2�,�L���U��ѵ�͌��l��܍�(0xu?J��iVe�Mn�}�����<�H=����ߚ=dO '�.��FO�ɒ|�H9D�=�`ʉ���XW�*�F�#�7�j�����	XT$V�r
��k�L 5�,�A��4}eu�H�
�D���3=��t�}�M��+�?E��';Y�\��^ه��5;���$a8Os�.��qSQTm ɚ�O$ns���a��RU^ i 6
��5���"�O�L�
�p5��C�����l��X�p��-vL�U��i�^�C�tr�8>�@E���k+��Q�:��W#7�A|RwN̶�� �8�ݶLm���w7U�?)Z����_��I��� Ɩe��ɝ�eJ�FoN
1�G"oi&�jO;�9�7KF��@�^���ʬ&�Y�.�1�ظ������k�Y�( šO��*�9U`$6g��:�x���J�ue�a��8�'�2b [�e��guSʗ�UĖq$���)Q�Q�����FD�����(FH �aG�S�z"N���S�5~z���0�	*����rF�G�+M�Eag'�#	 ����-u�'�@rw�`��b�����1�eg�c��˓~\Oly�i��1W���;�R�J`���e���Y��[�u���<b>[�����X�0��薈���L7�����Vwh�hW�ɪ{3��)�.MU�A9�$@U ���ć�����C�@&����{���sJ��Mh��C�2����kaq��k�Vf�hV�Hh)�H|�"�Mt�����/9Gߵ��z�n7/�6�\:�b$D��ڶ`˒�\_:Ղ�Ѩ��
>�������?\L��-��Qӑܾ�k{'�H������l@.�	��	�W*��;-`3����!O��>���J��O�q�6�\��
�y�<�L�7f^d��Mr���ߏi"Om�:.�E��<�����$��Y�����F��������p���:�,0�������w( y*����#僓~�����*K0A�KQ��h.���ƄRn�! �_��$c����*C��Pᐐ�b��ŷǩF��C�p�l)JSOζ""�L�D�**/J�	��I�9&��ԑ�o�m���MU�)�)N�f����CL�&ni2B߅��W�lr����[��r����:v�!$�9U-�
`�q��-��T]�t�[#	���� ��iB�f�Qϙ�@]�&j��Vs����Ń&Ϣ.�N߃�g�9�d>��,�k��e#��kj`5�Y��0�ѓ�W�m,���2݈}��U}@
׸�`�,_kׂ.��4s���?�/�y�$�������j;��ee�7Y9 ,��!��ޢ*��Pz�Հ,vZ�-����^�����}���7/����-r�����f$=Tus�Q�>"��4�|�⏵�=c�_(a�V��-��C[h%�#3J��m��	�(�&%(�"N�ӥZK,B�G��O
����ѷ#�4$3�nxE)���7��/Z����4,��J�2�x�	�u�RQ�C�9V˕�v����
����E*c͚�i�x~��yp��:V�-el�r�Pq�⩏z�C�c�� �w�NЕ6�K���4��֜�iZ�����p	�Ik�ӄ�R�zv79�v�fow��r�6F�0�\�RQ�p>�[�`�����E�r������d�X�YB����'������3��w�������^��O;z���Āfdژ�A�����4/Q�h@=<g>�x��K@�8:�y!�G�Ǌ�/`����g{�ǭ�Vc��~�I���8xv۰�н�c�RƩ�@)�~\\���*��o��r�_8����FuU���ܑt����U�s ��$z潍�
�Y�(������Tm����$��z�vefm]�u�Tr�kS���#r�d�]�Ob����S���~I�v��1�A����z�Deך�2�j;XbH��z��l%��ۿ^U�)���Ԁ4�����y���8����w���8�^��������{5N�I_ۊ���L���/�,�HA8q.C���$j�a�e팖=\�ᴘ�!`��w��[�c%�}H�d�[���c��(O�ƅ�(� �#��7qoD��mnS�y�#԰ ��?�4^�z'H i�JM�A�����@�J��;t��o���| ��M�8,�����M�/|����Iy䏏�F$<
���FO��U'��;f�ę���hmC3�f�O�W�%<je'Cn�l�:o5�X��G��������:1zy�#@�0���������~غ�M�og���p<�h
�&��.ڃ-[���jIcu����R+uQ�\n�X�'n/�zY�;���D��e��8.�~�'���%*����l-i$_zd����A4|%H����m�f��&;yF��R��A�&�^e�CE�,H|�(�u��w����
�+��Cҁ³Y�珬Uq8h�P�SN�S���W�1;պ���&�Tu�0G��H�{tZ�85�i��!��7d����ml���}tߙ3���yy�I�r��CK�\>�׺eOk ��Zd���ze��< �F��d\{�����}A
��J2΀����'���T��E�K�!�]�͗�xw̭L'�%y^W`d#�܊����FҢ�(m<�v�E�*,�)��;15�W枷h�/<�lh��"��8�͐�b
��ͽ۱p�J�JH[���+ dէ��*#)�Ab7PN���(&ο��$�Sax�{���6����HC��}�)%Zg�\H��FMz8ߞ~�&�.Q`J<� �F�/��[���h�(����.��� �ޡ�VԄ��7���{m/���}$h��oY�M�����K4찍wPR���6q���37�?{�Rm�����{l�q�&P��;a5!o��y)���咗 ������}م�z�^�Ő�dpIe��A&y~q���b�5Rn#�,�"A�ԕ��"p�@z��8y.����緮�|?��F��[C���{'��.L�?L>��}�y���2k� q���㘛�Ĩ�v�*�1�������M��a��$~/H-�vxP��6�m֐	p|	l����V�ٓ�j��ZS%�$�S�g���C�K}�o��#�e���;�N���C���+���W���AU�="�߆��$���0�$��p-'Ϩ$��*�ͨ�h��z >(iy=v"� ^Tq�������v�}�A��ӝπ�Eťn�O�n¶u&Z+5'�CL��LGz2�+U�%�_��ה�M���(HM�Yp���҂0������;ͧu����+(RK�Qa�K�BG�˓ŧ�3UQ�7 �΃�˗��а� 0:��UH@B����"���D����p!�5�y�ʫ��f܉jn���o'�q���M� �k
���ӺL�[Y��Y民r��QhqMC57= ��O�
ք����͡Q�� /dl1"��!{_��*²�J���R��(��+�$��b����4TM�{�=��u��&�O8��>�1
Y�q���_�N�rn�՘�yY+ݢ�G�D���{��53�%���A��e�������yӐ,��Ǜ���tuWt�S�>�VQ��t�����`�`ަ��{M7�}�Y���΢{��Uפ���S�Wс%]����f#|�>H�' 5�괼lS�T� ER����e�����&�d���U�'�p�^z$��qS�A����O�E�B�r�]�O�,�"w���s�[�',��s��5O���·/�����u^߸B0:Uy��.�Uk-/T�+��ɕƷS*tK����l��"#r&�Aa���رsb|���CI=�ډ-X��n�2w7Ae۩ɮ��S"���+��J�	<t��h�i�L�j'�����ǝ�y��k@#��������X��r�5��lE����)�I�"?G��OWHX�Ŭ8�@Ʌ��5��p���Bcm(��_i�ƛ?��E���X:<���Zp�\��s�k��w�F��]M���t��dF�V���x6&�G޶��ڳQӃ�zLq2S޽�����W�Q�5ݳ�-H�(h�O�?��W]�;� (/h��^N\B� ��j�hm�ܛ�m O+l�,��f�1�ʡ��r�O}���y.���6�)y�r���������/�1F��\U�k�e@�w/E;x�AW��ߎ�:^� o�Q0u��ܶ�dW̳���=�C�1_��w�[��ᆑ0�C�����{kꚅ`<�s���ڏE2]6��V�`�k�-S �x2��܅���k��)�ЉH�(+%�*$�0�t�:^!Q씣�1���0��=2�H��:�����cfv�1%��Hڲ���:!��k,AG�)�!�v�ON�R�3˱�id	��Ӟ+����!�n&�1�]q��M-w��gÓ֕4VH;�w-j
:��zc��37v��즶��DZ�"�l�Ӿ�F�p;��4P�t��;��Pɇ�:�������l��oc_�3I4m"�]'vne⇨�*����X���6�����VM���	���̾dX��"���������U���*KK�y���OQ.�{�@ �F?t��v��t�����S��+��s�l�VM�����6����0�^�������q�,�Lx����N\�|&�!�m��к&o��FK�����նXn��,�n���1f(�l�tW3¼�5����Ԭ�>ڏ��!
x�<�OR�zM�v�hf��Olk��g�i�Σ�اi=���=ݰ�{���
��F�)}���U!�&q�d��/ �u�5l�{�\�MBݎ�
aj&�~�_�{����j@���hϊw��H����~��ۥ��������q�@g�TE�=������*��N�H��-�s�v�L�5Z����x����`�$�S9�o}ְ뻷\�Yyx��/��j�z���6�4���=6~������"�ن�Q� 2Yfv׮L2)y�\ZZPUg��h�
E�_A�|�Z��l��ؼ_ȝ"���IJVr�>m�֣�k�X=��R����"���&���Q�^S�B����j��W���C~	��u6�Y�Dj�5qO�SQ��v&�-�kޓdn�O��
%*���W���&���|{0;fsM]�5�"����]ܥ�M�����#Z[��S�?�������������ؖ,���Њ��2[��uv'��δū�>��>^����6ﯩr��.7UWC��X����v�8��]�0���v���)Z�x�X��/L�T�G�|�GpGH�������?2=Mد/^+�'n��o��YT�y-{�	�kd��E!k	Xh��/��dp_(D�/�����;�ѴV�0��P�s��0㬋��O��~�
�v�I�t��
D�[��� ֿ�����֊
	1�� ��T��>����\%�{�j�_���88/y��L�Wv��
0n6#�#P9aZS^�k�I��BH*|�[	 ��%��S�Vޡ������գ�8]�Q�C��~���bXgo�q�&KN>��Pv��&��DQU{l*�"�vf�s��}{�6�i"dM�#�uid:�*&���ތ���^ӆ���c1a��pE��������::ߑ���VY.R�o9��k<*�6{�<+��n�L;p��ߥ
>*��rŉ�=�+���L9'}� ��p� �d:��M���&y�x��5X)�ƅ�p�ݡ"����?�D�Ҝ|{��*��z3���<�o��ً�d#6�H�T���o �}�O{ /�6��e����|��IZ�:"�z��uN�n~�y����8���%��*g��4lTn�P�H�F-��o
l_l*-��*��cڳ�	��C=��_+�8�I��Ӿ,�6�p��RQ]�?���h�����5�L@}֞n54.""�ڏ5�*��4��Oq�22��q���{n�kw�7Y�K���(�1-/<�dzD�h_�J�i��L��|Wk#�'�����?ޅ��x[�b	��g�b���U&�:Q��B� �w���6U��e�,b@)+�����s�_dg�AD`�/Bs�N�y\t�	���;�u�g3�ɍ�b�y�6���+9�_k�>�9�;��DX@�����]~���F
-�%�|��Τ���Q��_G��G����{SB��C�� 죂t�DaU�����<��*6AZvN#7m��gu�s�}�_�.ո+�R-�P�/eJ�fK�]��ΘGvF����a�����p;��9�y��/&Gy�􏋆��m���ZOg���w�C&d��zh#�:E_���-�@���ռ�f<�S�a�Us�8�t6��q�`#�(@���\h��R��4��#��X�[G��8��ʕ�WdO\F\J^�%�.x$o�a��^�fψ��W�2C	"��mgO�č�0��\�/5��^h
�B��X{ī|�M���
%~n���U5��;EU�X{�Ucߎ�|=�������-�u�L��l�~Z��Br����u'���Ɇ��	�ɘM�*��HUh�Ca�|d�����E��� �W�~��0�ө6�*�cL�(v�;����� �b��, ��j��(=h�5O��w�N���S��+�V�x�"	� ��Ei�cd�ܙ�  ��.�ihg{�������kvR�z�n1��c�U'��P���X�����}�*z��dӺ�Z5���5��أVt*ᑟ�|{+��(]M�C9jxK�x~YY<�6ם�t��o6��w�VD�[���)�l%ͮ떫b��� ��9o�L �){C�G-�{�0a pv@`BQ��L_��Kҥ�#�Ib�8d��^:�4���SOd��"Nz�I'�y#�cYVI�W���Eῳc���A<-a��,��hx����ta,+��柜�"�t����3>�J�ܐ����q�d����qqtr�s�E:�U�i=�z�P) 所>;�z�W)@m'�{�w�ƭxv�������!=R�\n[����Z�	b�`�b�N&����bM�����B~@t��cwE��4rz�y�ll��S���93����$�>�;Z����"%>���=L�3 ��r0�O� S�������<��B�
��D+\Q�&��a��Ǐ߈��4����?9�
3��h���k_�xFE���ad�����ʌ�G{Wn��xK������p0����-�"z���-���*�4p�P�fE�����-F��ϥ�B����xlC�,��Iyx&~��
��.qT�%̗��TA��O0���ٶ:�s�YB�F3&�[�xMߤL�fԻ�	�u��+l��f�;+Ŀt�/�����l�D?ia�
+�����?d���q��v�g�uì܅t���~'u�L�>��w[��=����7�R����C��;_�P���C�d�G��+A&S���vVX��u�o��3��A���xu��+���_�r�"ܙŉ1f�$1iݓ�ȕ�1R(�211W~�' ���a����b��J��cw�Ĳ�\��A����배��s���5�̐WC���6q�W;��*�����zUaf��t+�1��p��&;k:��ӊ9��:��Ѽc�wBX`mMz�g��3Z>v�XwS.o�_$3˪�j�	m%�Ά���!���VF����ǬrQA|�ک��C=r��jo�X��l��k���4e#o.x��z�=�v'��GP1J	�~�X�t#�y=	�����^�Dz�J�l`BԿY���7w�z4 Ċ{;Ӿ��Sk��*�:*�nOqȍ!���̋?KKcb0�W<M�p=������"�sv��i0T�yK�YE��򑐅��ne8�RT�R������Zl<OK)^M�k����3	6%T!vk��(F��{k��$��H���b� ,ɪ0��,}[D��95�l\�?������#k-aBt����L���fH�/1K�����v<�Cf�]ܱ�Ͳ�W}S��Q��Dos>�k'd'����B�IZ����3�{��3�d.���=ufX���o���Q�v����Fc>`ꑿo��2�ӏX�|f�!���"U	ư��+Y��c��ti{q�r�.�aB�o'P�0
L=���t�;g�!���u���;�v����E:��{Ƹ���MwnҼ	޼97ǧ]�v��!g�Cݟ�8WS4G8Y��_�d�a��6?��zG�A}�D�.�l���tFL�Y%����f�}ǫ��`-4��
���%��7��>�D]��:\|T_I���	躃��0�wr"jg\#^��.��</�M4�	�i[�e����8����a��VRP*�Q�f�;��\w��E���ߦ��-"��	���S���NX�@%�2�؜p���L�R��F|ܜ@&�e�����Rb��0�w��\�� ��)�^�u5o�0}.��Ѿ(}Rz �Fn�WDH^ǲ���c���	��q)���Vy�wB���L�E1l10��v�N�v��L��Z��c�f��z���p�Fq�%��b	�p�p
�����Y��%���f���xL�h�Y|Fש'υ�'jK�$4����ep��H��;�?�i�����.����f,,:q}�����5�s�I�Ky�xI�Ds����;���W�n����𲲹Q�h�(�N���Xۣ�$* ����Ht�@ȡ�
��zB��/;��[�ذ�C}��Ϟ[�:�:��P�O����9���ű�����Q����x��������^�k���rhtҚ
�r��|�A#�3!�7��'��7c~��+�5�c�A]�='��Vݪ���i������+>BWs�6�)�>�@�@cH�qY-�T�3� ����@��M���J9t�ߌ��^�e�{��ُ���U9�XJb����8pm�\��9��=�k���nS��d���y|�/�߭��p���^�"�[*PN�H�A*!&ޢ�� ��\QT�2E��p4λ|�g�S>v]���.T�o>�>]���T�b~�-��*�9T��Ԗj8�0�~�����!��S�����5t����­���$<Xy�!t�踸���E&Z[C�[|e#LV%�_J��*1�?�H go"u/����)(k�	�Ef�/�]�˛�Ȍ��a���	@p��HN�Q���k!���/�7��~{������-�<�&m�A�-�}��Mr�4���8�KB7�����2�.�O
��X�䳏�Kt��˱7�s�4O��n��@�+�^R�10[��Wm����u��\��9���jw� 7�Ϳ��i������跶u�b�3�1?��n*�)�wi�t8����w���&LS��x! �1��o��R�v7��hk�w��PEC�sҪ>L�tv�.�6۬��RVnF�k8Ƴ��m�PLIT�cDőq�N�!u��V4�YZ��,��m.�6�I7�_rM��Ϡy�없���m���r7�3��4tY[�����X�ua�`D*=�U�*g@$�R�^���u����5i���:���T�(�9��;3�.ͬ�s���@@�et	�B1�+u$�z*��X('��p�[�&���0SD�j!ס��ޢ5��������c
�t�r��}�BY��iQ�������Yn>s�3�%$\��w�'�>Uf�:�S)�$?%�խ{,aK��P�@� ��E	���<�}�F�)��5�>R٩�	�ϟ�R�^J�> ��,���PT���ٛ3��=�v��3�팡d��fF����0�	W(^G�)�򀑗H��Meg�KUm�שt�)͚GK��R��A�0g�."��~�x�iu䛉X��Nټǡ�7'�)&�fV��
�]*l�[�j�ٓ��G0{�2���`ȕ�)�\�$I��bύ��_�c�q@b'S�8D���`d������g�������'�"��ǈ��|r%���b|%�U���^���{+>��,�&�&����ڑ6a�N�//�D_���g�X��E�{ �j��a�A����m}wO�c���O�;+ǆs�Pp�6�h�*+�g߯�έ�V7�uM��<^��R�x/YI	T;��3)|ީ��Rc<L��h\ڭ�B�)�p�t��Y|�z�L-��ϟ�5�=�>�W7(	=˼�P�D�V%�5�h	]U���k��J������ܜ��%"aT_�Ȗ�����T���>o�iq�N�܂�^jO�C��������=Ej��6���d�!)�UgL^_n������d`Q�Bbc!A݇ �;�b�Ԩ6�=��oz����1�+1���_1�O݉��p&ޢ�i�o����8^�M���A�	/o��C����J��vq��3΀�Bv斑�d��L������4w�~_`�8>ުz�R��@b-q��n�#�f�A�3��!'V@�w���=7�pN>�2���&EJ,�I���`4	�PI�{p��������
2�~(��+:Ja�dGf�9��ؤ�
*�>��%|�_����ͨ�-��qdץd����@H�}��}%�,���kA�)��ڶ�E�M ]�@;��\�F��^�|D�٢��وw�9���t[�0\��LP�GZ'�N3y�v���`��X�Xsmc��}�*g,2��2��eS�ޤ�#�?�}l'��@OV4:p=}]��,r����I�9�������I����W�Ky�dY~`��)�t+��6)����D�JUC�E�+S�=��Ⱦ� ����^a�� H~@�k��q�:PH���+�e���XF
�Z?�]B�E�파t~��M�G��_��1���pS��3m:��G�6��s���7��6�*}�b�-���H9�V����?��$)���Xe��pX����޹����7��C^Z��!����rK?�
������~�*���}	�)��L�����ΊR9e�z
��,Y�ipX(�
<DHS��h�o�M4�pڇwJ4����qc�����9C9h�,�n%W�J0�Arp ���)���d�D�=�O�B��po�~.H���� �6:�J1�s^bU�7_X�W(�	ՍQl�A$�-qz;l���HG��шb��7�a.���m�U�8�����Pf$t٩E�K�Q�#>P���f���b���VE59��9u�}�Ե3��:	6�݊u�I�,�~�,�,��f����hi��fᓀ�M�!�0c��H�f�v{qh�A����S�W�����F��oX����Z�P1��E���Ri�f��%�>=J,����=qR[zc�l�F/�РV���U�qK�myr��=
ݝ��5�<3�Zs��8&�B�}D9���%�����ͪq�ѵu/�ԓ��D�1�)��Ghy݊V�� �Y����R��6�y���8���S2����N���vb��4J ¯�χ��`G�⨴�ގ�B}_���rqy�C�pE�nN��Yԛ3߷�k4���d���UM�^��.�7�B�UX�ݒ���;��tQ�a*�י|�Χ|Er�;%��=����?�����A�{���+�[�/��&M��������Ѳ�1
D:`]�4ր��^���r볺����_w�A��|h�[����<D�(��]A����'��ۀG���
&zo��}�������G��!��DXB+:\�H�7̽pd�?��O&����6Ĕ1mMH�O��B	[�O�1;ӦCV�U��k3��ذ� ~���[�t_>),Z�q�F�̖���7e����D-��Œ��V��w�i��C����J9oF�%I��p*R�����1�l�NN.���I�cy�4��$_h����M�C?wi��u�V"X���d�����n+����qU)�x)������ Um�;�se�H�e��oE5�!/T�_ĎM�H~'��gaet#۠�%�_��!R=0�@��[�/�8�Y�H�$��o��I��MV����B)<�tF^i���,�mꉱ�^�8u�Hg�>Y�%y�40��թEkYBD����sGx�s]�~NEم3_�	6w�ߠ(E��ܫ��^>]aQ�D*�?�� �\�>6�g'�.A���;8fz7�Ni��X��z|���p=�������W�V�K�#iL�{u,��7-s"��̯6�0z$9cr^���=u`"o_T7؃;���#
Ŧ.�w�\����WhfKԩ�9��n�"EJ�خ��C��uR�a �Ie`�Fp��o��ۋ��Q���mn�������%"3��%}�����JZ��w��d�VS�Ff8r��;�8�CZ$ �����z�x:��l�zo�qL�0���rH���jfF�R�҄��jζ��I����.wzA��roc�v�7��K[��=7'��P�'�R����S�}�>43$��i�> gd�%6!���8���a~邀�L
�`��� ;9-�ب),]�i�1�L%�¤�ً{q�����*�T��}��2�V(�،V�u\O�+s��u<������BQ'��!���H�O8@���,
H�t]�l�6���p�����U�b�9PIڒ��'iT��aΆ�����9.�����J�YywW�����:ni'{�f�f�>���p�	(�n�azZie�^����$�U2%�Z���)M,�E�~J�a�>�U���3m�I&u���	��b��ٶ�q�h��[/�oִ"�qҏ���~2���QTy
1q$0�<&5�Ē4#'q@��xH1rջ"V��HIἃ\��+��1]�/�� �r`�t[�%�ۢ���|-�.q����>�}���5� b�t�mq��J)��Z^�s|�F�@síi�?�1�C��š27��~ҧ�g_�,���T�H|�l0�hm &�*��~��V{�`�����~��N���/,7��E���`	�@0�}���S8GI1#�(��I0a3��,�x����\��vs2�^#d�"�s����K|9�z�Z���X���!d�o���D�!EeԖ�;JR�g��B�P.��i_c����E�s՟>T�7��d��V
�O~3n�9X���_����f��e?o���y!( ��r>�,��>����Gb��&/ ��6$�*9���Zg�`��]^T�>.P�Q"fO�W*7S~8`v5�,�"ăi�'�2.p&�-��*��?�#*S
\ǠJ*�>�ݕ��1�[t���4 ���-��4�!"s�M�*�\��Z���uC&k�!���gn%��{�|@ ��1��r�9��B�˩#��=�|ݭcrGZ]��zb��j+W�Z��Q�Y"����x�y���d�C�w���D�~S2��b�z�cp�yMz��C�����||�!���H�c�|�� ��5�~����e��L����E�������)�G:qï��(�2R�VA{������5��[|�
�*ʈK,�[��O�֭���7&ݙ 5ͼ�ְ-dv ���~�P�*70m�Tc��Q� t	l���P����f �N�z�<%[��u
fq��s}���t��ȇ-���?V�6� -H�w�ڭz�'�֡`*zsC�CHgnEg����$�렾�`| �.ą������B��*��������<'2����=�`m;����Ϳ�3;��LF�Q
�7��֘�=�K��DH>Cb�V_��A��N��'��V�"� �pu'0�Q(G�.�D�w�%>#-̳��� 	K�����9yY�U�<��D���Év��j�
a��izv��	��/���!�o��h!)v["@���H5C���������8���X>���!����{<�_�4�-����s*��S&U�EA,)���2��h�^\������R��4$8�s8VͲ3J7
�Mi���X�E��w��ɒI�јeH=�,�D���Z�W��cȭ�9��<�u���V���%�B��SŞ��S�C�,?����qF-��2�@<�ڕ��8仧�fET�����HX#���w��nx@0�n�Ana�3
�r!LgȓG�u�_ZC=�*�걉����n6�����j��n�m�$qz˸-���j$����c嬷��LF�p���'
�o�c�,���
���_���#���)���NS(K�4rtf�(ށ�Ha���K�Qw�f�pF��d�vY��X��470���4�ɀ"@%he�yTv�ïY����_���}б4#��(N�wU랠����#֥Z��T��-N�	:�m�e�\�m����}&%�~�d��#yx.����
��\�x匕2��L�-T�b�7��I���Z�O搲8��S�CM�+ub>�p ƞ�"v��(}1 _�>>1����\[�c#ő�k�3G��'�=��[Mɖu���(�V�T蹩r�
*:I&#;xr�t`s�ϛ�F�E����A��9e��U���6�����r���!��ZI�:ڋ`�fh*��p+,t/��K�O䁔h1ŊA��>m������/������o@V՚2�WP�h2�����Ag�����~���U���_���0��9��N�d�6H���,;��~��&�&*p���)ο��QRs}�:��C��.�7"�i�K����ō�R�a���5f33[�o�/�87��qD6_�,-K�u�����͑Z�fT� !� ��I���R^��=����R>�7�">|�E��a�{�.�<w6�PA����&��D�ꍘ���
�Anep�j"_)�2~��RW:[:6�! ��E����!E&.�J���r�=&�^=��$!�ù���N�� 4��b�)����h�5��H+������~��Uf+�s8Bc��#d�%пT��Б�ԑH����_¯ϫ��qsj���]��;�k�[�lify�nZ��\���z ��H�Q�]�v/��Epr���qK��b)/�*�n���/��CxP���M}R�D��t�@�}_�g6�Q�Z��'�·�8w��-�����5v�w��g[��@<惸�jE'V�����b�W�2� E���f����#�4�N�'K�G7�'�����W�W血��7=\;������,�#���$5h��z�c����ur��jA��y��
�͑:~���b$.pƺ
� �(��7��
r�I6�<I��Cɟ�A���j�@�:�<�
��Q�|��1�Gʖ���R3xV����ף���
a ���Z�I^�E�N��pP)�|�aBO�G�.�������r���!ٸ�m�r�l�_��8�t�z̳��d��.�R�[�%S�a���6A%�X#yd�z��A-���l�>������&y8��[�?�������*�tm�˽q��
ڮV��N�O{M��1���2k�zj� �Z��Ud)�8��e���8��c�� ���f�"��cW*[~w���Mʵ�c��J,���C�Y�Z`�ԩQJ|w���Vl4��	��A��E�Q��br�{>r:��ɓ�>�!?�eq[�ѷg�%E� #B3�	�|H1	�J	>�V���b���d �1��Jń�kQ��	��D@E/jOf��AW�Wa,��)]؄ˊo]�?���j��\!�h�*y�w�����P���c���A���g	��A?Z�>
��-߈�7���D��p�`��L,�Ƴ��|}T��)|f
�L�5�`1+H��Eǭ�4��h�vȊ�q~!\�(M��lJ�����{�j�6���KP�bwy��5�%\�e��M�ߠ~�8�I,���?Լ�,���[��ad7@�
�*��ߚ���oo4�����\���acm�U4�����-4�WI(�tma��#��HGE�;��-m����d[�zM	�9/� �WƢ#I�� �l�~"nI�\�P��b[LE�	�u�`��9���}����8�β�!��%S���:mo��x��z �r�� +���3[Kx����Ļ�;-�l����Aх3����ؕ�鷐�3?��{B��3��Fф�#2��?��Ă��}n4��|A�^�I����bh ׻���.H/�J=Ȕ9�ald
_C��m#�/���,*�F���w�i�ƿ �B����={0��:�6)s޹#|�u?�|^�:�f7�^�*W�֌�3���̐ͳ���,�0����Վ���cZvn[/������tu+�x��	繵Ю�[���>z���)���&�7&���DT�"��׆Ti��)����f����%�WɣH�?�;�˘�w��0qEǧY'�"[�NΜY�t��(7 b�k;k*+���AK6��~�]_����K��N����}���O�T����=�r��E��4�]<Χ5�q`P���W$�禼��a�~�i�br�pUzօ��x����{K ��逸��՝>t�̋�m�p�z���Z��dv�4L�_/��m;�����;� ,��)�n6 ȉ�!�;r >4�'���N2�I�"{�3n{����+v# G��nlE%`UG�����4Sj󠘀�x<��MxX�´�ՈW�(O�����G�O`���G:]ˍ���)��� �+�V$BSgM2��7�xp�#��[��v[��U��U�1�s�ڎ���(��iw��>�\��n��[�B����9]p���vgBZ'M�W���DCC��d�C�a����������[,y!c� p?Ll�jmkܷ�$[��u��̐�r�o8�����0�\AYUg��ش�"�+���v7��L.�S#��I����{KJ	��s�FIo�(�� �Kf��g�7-��T����p��k��闱�DF2�Ɔ�Ӳ��D�)հ�E���7��ʯ ������ؖ�F��e%����n%4�NQȜ��v��6֧���,%���ا[sT�a�{�3@������F5U��N�|�Ɲ���H�޺�O`�x�9�^<�������������� |�qSZ�f<�����q�a�7nftĢ����C�K�vIPg�6���1xU�q)KG��,�
�2��lz��$��=r$^&(	�@��� _T�9�%���������l2�<����o���!V��ǝ��Lq�[�w�IOzL�f��˔�Ν���sq��9��)����o]�����Y��;�{���c|�[�l��ӚK�	����a��2�g�M]�t�������z���`��g���!��w+B��w�׺�����?�}CjqL��Y2DJ�E���8-/[�g![���aE��s�L��3M#x��H*y)G��(�Gܖ(�9��!����K��<YF�8^^u�p,.�u������	_�@VU|-�#�L-.�qS�-Qp��)�~-2\;�vQ��t��+Ѱ>�d?��q�=�l�4�����9�;R1��U>�8��Ƀ��$��nzV�Ր���ϻ3t�1z|��7,Q�U��V�c��o�e: �#���)��%�����R�:��"U���A�������Yh�`�ƴ�c������H��;i�k��,�Y�1�*����[�VTr��;r���|�E��>�lnx]rR��&=���*�lV�*�ċ���JZkZ�	Lן���;����tTi��_I}{�&AIF�M$
^����p�z3ۖ�v/��ߑ<X���c�����"ÞHb�Zk��wf l��؏�)��߲�W╼Ks�H _�yK������%�N�P�Y�ߢ�c��p����8��5M��=�"h����ӷ}+s���;K=J�+P�����K޳P!U��2�S�/*L�*�O��gF����{ɴ�bi���@�A�����Y��'������$O��aǹK�Taq4�s�� .@���vE��N�v+~��D��P>�4��R�]?lx{!�����f����PE�=�ΉAB�����/+�j��E0۶�,�(h�8�[<y�Tr�������u�^ '�ho�x�5�=.��jD�����dW��&H3�ZH����=�>������_r"��K�@��������/�ǧ8͙�7Þ�7ˢs�m�O�I���^!�ݺ�(/�RSGz��GP���m4��s"�������L����Le�e|T��9$֢�@=�>R���G���#-8x�gX&�-�	��;ޱ���d*�"��;��*`F��\ :�Ax�dbE@�����s�F�Y�y������ �+qd��ǋdߘ��<w��z	m�,=$��
��=ƿ�v�	��CR���n\Cx�:W�;�5�����*��p2����	����(�zn�
i
�w�R�Gz<�����5p��vf���'�n�:O��]WPp@ ���v��h�p�3tȄh��OW�ό_M�����P�Z��q�mZNM���w���W�Dr��TQω�^ �k�6�+T��$�V-�EE����V�Z��rLjI��yG���#֏B�',�����)�u_�e��@�I"g��%�	��Wh;I����o#�)Q�Y]B��aMJdMK�ןL���w�3�0i{��U�����z�k��DEn����5=)�A�Z�D<y�ar'-��n.��/wf"sd��	��d{+U�D+���
@��p7��ଆ~Ό��lr.�}�NY`�}{�rBe�go�S�Ȼ1]8�>(�D�w:!F�u�:��,(���I�(}��Z������ �Dr��"=�Z6h)Y!Õ�kB���*/7O	���8�����}p�E�U�&�1E�l �e�ꉓg�=dZw�Q�=�{�7�m[�����t�?�5_l����V[�iU)�s���ٴ��\V��=�f�^��X���+����������k�7��`�.�l���C��b����'!/ �|����i�б5����kK�d+���au}2l��� �N㰕:�4���U~�@��.�}�<d0(�Ķ^Xu�g���2o���	u*�w�0ϣ�ah r���"�<8��� ����Ҧ4��G��W�$-ͤ"��3�:b����0>f`#7��"�F��q����CI����Z�k�vy�(0���%K2��EM��s���"���0JQR;o@)���2�d�Z	0?p �b�U$n���l�?�þX��,F��H�Û��$(�߀��478g�s(o��Z�����fgǄ�i�ɽ��x2Ք�/���`ޫ�ϲ̘�nd��q*�M���#R���ܙ�>��V`>xL�J�Ѯ��@�~���˹bN�}3'$��"�?��'*]�MP��ZIO��$tM���dΩ$"ߞ��̕i0[ta֒c�\��]������c���f��8�r�L��{�o���K<x�G�,E�o f�c^��T5�]�,�]�o��?OdN����9�[�f��83��'�%�J?a#�!7�ޝ_S��?=�VW3C��d�S�z*���0>�^�U���o��JA���~�V?yen�t��6OR¿?���2��P���&�����*s�ʦ ���J�B$lᅋ�T�H��Ēz�Ru��v�akg�JԢ�o�����#�)�� �7+�_}�,�!�E��Rݲj��o����c���5�<m�̛ƛz�e�sA�9w+k�쬄vk&�\��������YUG��x(=!��$oWU�Rz��^*���F�I�2E���!pʰ-�Եn�(�4�A���\4�N����%л��Fs@`�dQ/i�����A�YJ�W��_�T�Z�'��"�N<��~�@_�R�gO�9?�j� ~�,8і���>���Z�;����p�R�zОlm�ҿ�,��Y�u/���~*��]6ȱH�ɧ�x��VB���2�/�������'��4,�7��ܴ+��H�M����&�4\W�����B�	�2-r���&�8\�wk�<	HU8$Em�t���ʴ *-}��.GƸ~�b��5�1�j�c��]9�|�iCF#y�4��k���*`����/��!=�E\s���X��r4�#�b�� �?�:�\��m��3�e��B��.|qN���ð���_�b=�U���ݸ����w
���/.���<s�&���{����M�n��}�Pun9%�Ϡt��g.�Պ�y͢0�b�Y}�3E���lz�+�'QKl	8���ܹ�����8N�8WS߱=x�� �%�	X�Le�[�W>Wό�dj�PŨAJjY�n�~�\�`2g/����<b�e�#{�)����t����b/,"���4	B\f
��4+�#�	�_~	�E[f�EeL^gҏ Z%��Մ5���83�v���P�
��,\��T����d�j�|�6���*cr�z�J�V��c2�ӵ%�R��g����C�w	�șW�O=#sZ�_�8Qx�|��s��_�w��	}��b8��&H�I�r۸��P�K�����1��:]�S��z���0���H�����<_p��3������^�����$<JW��+%��L?���.!���
w�{$A��rήр������Մ�~S��KBh�m�����IK���%��yDϛ�闯�/�9qA�ho�Z�DB���r�"�����¸�pwg�}j�O�I�|�"�=�Z�e��e�NbQ�L�\��b	���*�׮�+-�)!()|�������v���0C�h���p+�;�0�_ֵ���៶q�!!�q��Bsj�1�9rG��[��+�͍���+�zV`���D�R��TC����/�b=T6���j��-��ed�z�u�X!� ��6��+m�Yȧ�JYXPXE�x��/�g5������:0( �Pk2�ɧ�Sܗ�(�f���pU�����eSh�E3CO!�̔�����GQ^n��jA�k��ɻ��%' �t4�?�����:R�H��ѓWIw�V���{/���$8u7�S\�	b,]D�Z��"ꏐ�r]��e����I��'��#��&�DMAh����S�oN����̦����|{��a^}���76{��cl!΅�,+��Y�V ���I����%���f#*��"tn��7|��{M2�2 �����] p+D�_pj{s�i�+����E�
�&�"1����,~� Dbߧ�Ǔ��Ը��~-�(�u@O@7&��A&R�I� �>[x�V�Zz/ �cSd����"��x��ﴳ�T��_~�vE�֒3�S�t�P.�����tp�I�&\�e�"�a�7��g�0`�6��������kƕ��7��	l1��6��-Lsv+�06��s u�h����f
�ľ�C� �.ɰ�V�,��7@� _��y!���� �f�R��JG�<q)�,%�~J`� ��f�X���Ľ�����-Aݣ�I.��y�GR��q�e�+�����V.'�f��^y���o�n/6s�Lo.�DfN��X���v�V��ъe%��N��0����~�|���_�����r���:����e3Ϯ��o����l0|�Äj�KM���e{WE��ӺH%���Cd,��������&؊��p\�������&4q�4-@o&1Id@^_��]b��������J�I�IH�8�*�{���%7��_@RG���za9��>�<Ô[޽��D^U��ƥ�����ՅI���L1��v��)u�kNr��jv�xd)w�p��|S}�n��Iq��$��:��|]6d/Q�ڸ8#�����I75x7=(�E�g�� ������˳�����f"'-��sɝ�\�b��w&�L��1�,/8A�ź.$b�B��F��.�EXE�e���Q:���Z��~n!aZ�[�sr���)G���)��e�H�W�
3�T7�+,�ۜaT9E�ϥ�]�hT���h�y��@��cy�;s�U���Y-����/�,�`�7$��K��Ы{��_���+
�f����s=�1V��m���ߚ�V�	+Dgx���/���~���J�M=8π۹̓Z��w�����飜����?SK;`aFqczUd��V�N�݃�{%�(�G����8��xG����G`֠2���l{%3Ӂak�`��t��o������8�?B%Խ�1dR�#2�9|���/}ba�u��d���`M�ʪ �d�#��X�����f[k�� Ѥ�bbr{M�t!#Q>2be���k�s䘭�:$����wi\_�0o��ڸ��� \��՚���u���$�
�S����,��^e/m�0���c
y�%�riZ�mþ�����ɸqI�!S�HF�0*�#�	�����p����	�B& V�v��?�</��>N�<���o��j�hM\e0z�r~����	d�,�4��T�Ec��լ)��� 7��.}*G���Л����S� K�@��PQ m��9sب���T���ny�R�4{H�ͦ�eʸ�8��?�^��N��'$o	yclV��ӡ�0��/�)㷅7̡ �U�ח|J5��'�|p��T����0���G%�]�U��~O^�����(��D/�5���A���Q�1J�q{&�Ul��n���[Q���8v�.}Qs���V��O������$p�s�;\���FrЄ��������:��gYnR7u���^7��e�2�b%,dｩwZ!S{�$j"��ъ�d-y���n_�� }��<��hI����������v���D�v\���;
|Z��C+���$)��¥��[�#@�6��[�wQ<!ؑ���Z2��'��_���L��&N�90�b��<d�O��ٙ�hz���J��l��*��+,����a�Җ,����w��]����G���8
��w�މ��o�����
�08��/r�2��Ə�4����1v�����O&v`��(�	� ����6�R2�va1y�]��*(b�^ ix�����X�nq?M���_�W�U�j���tr�4[�>)�!�1��ˀ�?��
Ej��6�
'5m��AY�pw��+6$!V]3{����%X�;@��'�"���� {)�Ta�4�U�Ƅ�U QH�6����Jw
�.��p�)U&���*wX�������#JH��y-�N[H�h�1����kb%���nEU�e�B�`�t�C�{d}�#�mrCR��M`�j�u��r����ٓ�[��;�ݳ�b �}���~�ޠ���%��LL2�63v:6���F�}g��s>'l�UѤr�L9�?����bTu�Q��ҽe����U�:�����P����]��v�87�h\��6�q5��,�.j�O�x/6GPΓ����#$��`�*\Y'�U��T��3A\{��,�@҇+����PN7k����5��6�JbQ!�zI����"c}3�����Y�� E�%���O��Pʹ���d��yzaN�E�Q∸w��
 �!U[�UR"�6�YܵR
�hw;�L	ٖܺ5����u����n�|[Zh*��]ڸeQ�ڟ�J s�<����lQ�_��5�^Zeځ���I�;ٸ@���=q��6y�*a�"��퐰��xf�E��~�"������_��ĩFh��`jP�*�a�Gl,Z��%��
R4 /��RG���lg�D4��+���D�6���G��k�>�7��\B���D.��۔*��q��װii�&n�0�"�g�?��(r)����s3��5+�8sX�v*���M�7b2��&Mvb5�!k����J>x�&�PX��w�ڀj���DA!Z)����a�9�Hs�R��n�\��ū3��<�v?�(r\j�@!�<��D(�N��FB��ݩ(B��n�6W�x.�����hKc����u�ذ�&dG3�#��)�j���[zi�����@�[%D-�}t:&���G�X	By����ܦ��kq�m���Π�8/�����ސ��Z����vr��^F��J �&B/�аE02�����ėҠ]��5r�=�6K�p��ڿQ��@��G��UMVv��)�k���" a�Z���K]�\�1�x3�f�,=t&eX@ �^�]切P8V��iG��YYX�"$aձ)��(�8j5�}�vXo^����(��s������<q^w��\���6���gՠƑ�,�>$�ި3�Sdb�L\]4H�\�r�5�N.dA���5f����oI��ᲶU0~<���� �� ��3K�!J��19ㆆ��1`���k��-�^'9�<����!x�v1�)ے�C,I��/��Y�=lO��6�l��S��3���NU>�ܷ�&T��kOI �|��7�'�<�T��W�`4(G�5���+V.ȤO�"�<��lPԧ��H����I�Z��n��ʴ@����Ƶ:��P�|cv9���~���q3wnY	r3e���F���>�ʵ�Q�3,��ҍ��� �_@YX$7�	s��ǋ�o�}c 2�wY�EK��sG*��~����4Ҫ2�+mb�+��z�.l�+��@f��IK8�ߴ����9�v��լ|>~[�^���_�l�(�)qg�C�<��9��@]l���˼c�m�5���9ڒU2)�����֤��d;ˈ.E(&J��0�ѕ�b���L�[�A���d�	��R��[H���h[�S���V6�R)��yC�l�l���{����U��Yh)t�p������w�(�̨@�� 4���Y�Tf����� #
�����y��1��
\Zu�۔�r¿&M_&5���ŉȋ�4�����x*�e���c�*�k�c��炝xz�-F��t����V�j�5s�h����O!���,t�(�aU�ǂ	�x�Bx�ߜ�W��+ݖ5bdE&�^� �Sn!:C�.j�'
�AJ:V���f}u׵�"�C��A���Oߓ��a�}�o� �ia��Sl��6�O*�x����sH��4�i/��9�L
9�e���S������|Ք��_O��t,ܣ���1�2$V[��1p"uP��{ʹiGm���Ĕ���i7�>E���p倕�;Qo���z�#��B��-g=-������V�6c���,i�Pd0���c2�E��� �>���$����2�h�4j�$�}������b�I��1��#���v��.y�Zi*��qe�.8i}���4&�5mo[Q	�d�'GVk�!/JD=f�&��`h	�y ���-F��)���s�sH�q	�=�bJ7y�q���6%�\����vM� -]�z��tF�Z2�խ�m>?����W�[Q{{NA�)��I�����uqӉ�P��K褍���O��c�����j�8�u��!�FJӰ�C.�&�#��JA��6Q��A��f2�`xG� �C!�I	8W��w�޴p�F�.����#z����yGs�+��B�?��Y��F��*T'�ZK���+KK�`�.A$������B#�*�3��2��ve�{���c�ؖ��$6���h�/
�z���<	/��`<]6����:�>a�x�x!F9�+��λЌvrDu��s7���gMN��i���2��:�`!7����@4Ԧ�%<�_�,X�äK1A���D���dt��������Zdxh �--�Nd��S�h�t!��t=��%9�D�X�V�f2�6�	b�2�v؜eA�V������Fm泳��Ʈi�����ܜ� Z�y"�,R:3�S�����K�IB��Ê�-XX���&wӵm��0�g�.Ψr�luں�gZݤ0��Q���Q��o6sG	���2���Qr�x�N71}_��yJ��'�D��A�ח�x�^"*�4$��܋A�$����I���s	�䥗�k˙{�e�>&�V'%���EY}>p��|�(��c��vwB"�<͐���8�&�.�!����.<���7�ǅ%[�<1�<��"cdQ1�`m�u�T��O���܋<	 �su�.���@�%Үtja���R��l�Ū��Af�PC��b� �B��8WB�M8:L4wq6Mw�Q�u�J*��۸�p.3�ʋ�I3�C=��R�aLEw~>,�1��օ�?�ɷ��?&xG^�H,.��4	}R� �ћE<��-�`���+��^�9���L�&Dѿ���t�t������;�M�K`5����έ㈚�R?�3���L����F�ߠ�+b����z���G�^�jA��?�*����?�,�Ѥ��b��aZ����L�U��r�	.1�2�//z�/��&�r����:�^��A�����N���&}I"�4�8�o�#:օfhJcKJH�Px&w��&�=c]�CF�*���@��id�$��Ԣ�`��WJ�(����~���� �"���}JSm��QM�d��S �ˉpk'H\�B���Si�`��,!ٗ+����6$���m��"}��8$�%�]��Ԫu ��S0�B�/@Vh���1lP耝� � #<��mp��w,�ر-�!^���e@@8
u"��ln
�R$O�:k=��$���?K�S��o�	��J��M�H��x�"�m�;�C�&��f�U��/���ӳ�t�Է���K�,�s��Y�#�:RS�m����J�e8j7��Q5'B���$p���a�@���� �vי����3�ރO���[,��"[: �V#Ry�0h ��Eo�!O!�3�0���D���Nk&3b@���B�A�^
m��ox��j�~����Q��]$�N�~/Qg�ԫއw�����5���N���AΪѩ�'+w�a���r�]o]�E�Gp}fȡ5����)lTax�����K@�Yb��o![��N��lV��g(&r��RpP��4c��_L��L�3���MI@�D���MB�bD�S�[��w�	�z�>OާT� �L[�ʠik�N[��DIc~\Ⱦ����I.f���F�����y|�<)4!䙅^�������X�_����/�;����$$��!�~���G��r�{��fo<G70u�<��h����������?G�B$	��K����%�6��L�~����4�����./r����V�N �6�o`�3D��D-�F�k�u˯���|fm\Z󭾆bt&;n�+:���	���IP�H/2s�섒���x�������+��=��ǳ��(� ��~7��ϭ�E�
����K-�4w38�\����cL>L�h�j!C��� k[��]'^"|l~���i���)�aK��Me�=��
������l��3��E;�ޗ���1���-�?\�!��y�w���d���m�S����W�aՆ�<
 ��6�_��g�Օ��}��Ks�I�6���7���[�'��M���zR��9�rǸP�Mb6�Ѵ�r�p��W� #���wY06K�m���Ա���PK�|[~6H�|�7x��s܃_3��&�'X9�T(MZ^�?���`���+���*}.fN���������"�ﮞ�+x7Rm��À�r[g�<u�^�L_HЗ1����{rK�\6�bRr���]���M�m�V�Tb��&�Sܧz����RG^I������bU������8��W/�c�x��H�KP����#=�нs�crS��m>�=���{jW��y�P��(�ۻ�!��u�I�g�]�XG$@��{�k��O�g�U��\M]���f�ڵ�\h�,,*o�2a)���xgl�ܻI��X�܅�����T���}�r��r9��@�!�-b����	C�:��E�K\#w��m
�"xl��(����y�����Z��V�#!)���-�� �Ƒ]!�\�-#\ƪJR`�Qrdۘ�k����8 j���ŷ�xH�pt0]9������~�A2�g��r��E�t���&ܚΓ��$��4+�d�P��B�����?�2D��r���P�{w?"�O��_.�ڝ�&�-[��ܥ�ޜ������I����B0�۲��K�k[˙�D���I
�����B�p��Br�$0��f�.�|���s��3��mfiH��u&u����Z5Y.����17�[��E+���*ho�v�sD��j�٫�<�vQY�,B������{����L�����c`�U�����D̚�A���+��~���MI����B�	���דּ*�.���@@� �r�T�*Z ��Rk�8Ǎ�
h6a ��,WLN:6(9��Ǝ7E�(�ntt�fM��#ф��h�i�Weӓ^��_��z�;��@���Tk��u�#���.Ő��mAX���WGMV/f�YA�v��(Ž�W~�`�g�<;Y��2�C̔���+'d���O�3V� 0M\+��t�kD�sm]Pe����� QXb�a�X���'�d�
�������~5�9����&���Xv๪���P	#8̈́x`X���h�ͥ�:O�#��{濽&FL��O��}�y��_�|Iw�ĴYÐךC/c�G����}��h��w��z����7#nӨE�yT�d��J��L�����OVq^v �?}r153��.���	��:�1�g���|�X'�h����gM���'69�%�)��؟����yF��1i�)��V���<�ӕ<�����s�e��G:��izE����[���t�<6.�oH .N"<����p�OLV��MA#<���	����b���oQ�N:��0wr���Z_�S	�-�,�Q�����p��̢&�v,K��&=�����LN#��q����l��.��;a�4�|�=�(' NG¦�^�D�hهq�~�F�;�pv�texm "�h��ǀ��3"y��.8�X��ؿ3T�f�nx�&N�ʿk�E��6 Uc��S�M����􎌜$#ӟX����pk֔M=��|�n
��)n,�%Dg�,8�'�����@��Z��-Ϡ3�oL�����Q��Ԭ)16����������*D�z��-G�
��u\��tT���~��BO�:2	�D���#��s��L�:�=�������Z�$!n�Q�)���F����7*C�&$N�K�D?Ko.>���栝Z+�(�Bg�j��ͨCj6M�: f��!�����"� �8�0��79Ę�Vp�%ey"�}��D��wg2}�*�,��qm��I��?��2��*�6��Y���!�jYǊ�YL�����d1���9"��>\t��� _�������o�{��^��Pd�=�gև��\����Fc1�-�7�d����%��%�m�{JAx�s�18q�[B���z�wh�+�~���Y�{��l|n~��v1%ފ�8�2J��`W��<]��� ������`!S̨R�xG��˥S��⁧��s������u�����/���,�e3��Z�4�׹�6�m�z��3d%z��rAR���������\ds�� D.fT���񰫄P3}��[��8WF�Y"�_�Ɨ�I���F^�!8ڶU�0��m�W�#�X~4���B�/i�.#=ԍ*��=A��s ��)�;]�����H�v���,��$l�J��N ����j��j�e�E=��.�������H����aa����jн�r�e5��Iq`XG�<u�]���@�'��d�$2�f����h�"Ýy(���4#�U��ѿ}@�>�d�� OCw;�?v3�V��L�̈́f��dB��_�g���K�X�=���
���Gmzy���~�.�L`��y�9/ �a�aD�z�j���M�W���A��LՇ
�~��$WRۏ�=�"}��T����ɝL:��.��٘���-����uZ4ӫ�o:R�q����ԽZ�2� }��$XiѺh<0�7D\�cs�/����t���������P3o��
J}3���`i��YR6�BW���Nr���N�؛�q�X�-�i)Β���~Q���:�#n�$�Y����n��9{���$�J�8�H����e��h =��b"�]�߫s�Z�*�s�1ogX�6	~�UZo?�K&v�2��O�� H��Yo��,5��-x����K��}V<�́;t����aQ
�&
m, ���ڹ�G��I�vw��]��s�W��W�gk�Yo8�u@E+腧���eQ'Rᩨ.`��F�����ߝ��N0&�l'_e�+"�{3}�!\�g*>)��0�4����4���u[M	{����-��Dn�sH��{B�Е��#UY�j�3���f5������epJ��
;����N�-LO����sJ��ס���֠ǩ�<ʻQ�,�QC���R��1^�?ͤ>�Y�$��,,�W��]ߛ¢j�z܆oj5�7���Nܮ�L�%��5�5#ʢ���j�]�4�w�ɭ P��I�)Ѐ�����$+L�z����u��|��ֈVV&t�ʓ8���)r�H��DE�rG�Y����6i6���I�ε����W4�:h_�D��&��FM\_:�`�������!Z`"�jћ�]��l�Z��v�ߣ8۵��O���c;�t]���P�R���x:�3��#BO,���!���j��Y���.�H	Q9���ܶB+p�6&�[��d��ی��+!�۫|�]j>q(Y�_Ԯ�<���7{ϳ��R�6��D��ŷ+X]v�6�H��FTIx��5F7f��Nٟ=۩ܓ7����^I��D����]1�iLT9�2Xwg�����ůK@�����re̝��?���\_�s���&�g�5�_&p^�F�-��B;�}���	��� ���y�~zH̻\T�2�$,������xp�
�#h¼aW>�AF!�dL����F�}�D fcụqX�E�SER��\u��"�{�n#H�ǣw��m1ފRE`�E�w�	�ޠ�n��.]Q��� �U�S�# fI줴�;B�������u��Vd�z�F�̳�)+ d��*����?��`8c���2(
��7�SNu������G�,MYm\�Ndm5����&,�m�=�-;U�#s�6�dKyzrrG��E�Eϼѯʍ�a:0��7g�f�O���F3�̾?�t�`H�f�.� �#"���K��-�-2��#�W��c���x�9_"*���J£os�%=I�d�������G2	�G������1�i����߽,���o1��벨TtH�)�ہ9�0�A/CԷw�L�s�ꡟ͠t�Y�<���n�>�?/��o
����2����ˁ���_�7˵Qrck���R���<��`d���^nt���z踫[�9&��s+����	t�`d���p"K��v���	F�
�W��J<��^H��"Ӌ9��f��4���[)�I	7����y��N_�'~B,�u#�8�~zS�v�`��W�D�,����?�?sF�Z]SGD���_u��/�[dc�.��1�#�4kNJ"�QW��D��78?E��'��|���i���S�C���\
	B�s�����x��A;��'��^7(�������@<�`��"�h���0�TwzbkwD>�kd�MD"d���f+��J�������I�䟍�^]4�цC�+���~,����~��JS�W��i�Ii+�kǫI?ss���"��u��� Q��H�,��ʽ�Hz�&a
��jH�xކ��.~'���}�'Nl�O�[<����U��/�7����e�NQK>��=��&^�����q���+#`�s���DaJ����4\(t���E��EdpD9ь��3(ih�q���.�Dm�bev��"t~�ut�]G���Vt6s�Z(�^��iVb�6�8�t�M������.ղ=�U�v	Ua�DU�	��KH��c��Vs��Ry�U��P��a�(���'�ɏ�,��r�/Z	fxl �d��yv�8�_� �N������y���  ȝ�k~���&�.�;"1�q1�R�s�K=3 l�mu{g3m�Ɍvo��-���H+���tA]�����1f�,���0�l���0�4P��MU
qO�:�����}jz�kߚ�EI�M9WQo�Z\��DS��$N��2��v�H�4J! ��H��+�T��v����5F�Y�2��]��~[��$�|�l+�׏c��%��x���~���Vzr���9�Z��V��d8�G\L�r�,yvlaޏE�{a��܊Ǟ_
 �w0��z�4��=�����:����|�s2��k�ʾ{Rb+������|*�K�e�h�l�Qm[���5�}�=O�Lg`{κW�w�S�3O�~)���_���ηp�y��<�Թ��?v�Ց_�e�u/h_��!��Y�1���֦�G?�zIv���/*�A���$��<@��K�$�@+L�S���u�&�u�d�=rn8|h�z��6�7����(�D��?r�KHpqOwCn�����$Kf��t�|^K�D]���I�ˤ��}�ilX�KB���16#���v���e�'������D��� ib���!v�̈�;��Xe����T���\vv�6�E=3��|l���M/��9!$\�	՟~?��$��J���p�4�{2�<�oE��T�,+�!�&+
��IQ㖔�KIk�S�����f���)���5��l�s�04�I�x���{�Uw��ۥp��9�yD^\���l!�sK��}��s��Eԫ��G��s;y*�cd.p��Of5����[�Rn�����HE���M�Zt�HD�Q�H�Hh��5O��]&I]� ��"��4�σ��
R�D���(,��!�Y�<��U@�k�M�F#����Aڣ�5D�'�}��[��U����9[��N���J8�]v���ғUh��z�fL��y��W��K��/��$`���D,;=f~wZ���E�8"ԗ�%yo�RCf��G�:��e/�����UU�%��<A�*}��ʽ�o�ӵ~����j*Vr�kv0�`x��	�8�{��2�BD���w��O��2����Pv��� (��dRm�)M�����b�;�����"�B�b��m�3��LN�4~�M8��/�!��sЄUvMnP(�4��1~WXm��«s#EG7�f����.�,��$o�t���5�����QB1�OJ��d�J��řy���oJ�7��7�)㺕�ZE��l�j��5�W[3����y�����<����j ͔�P���� �R�Q#U��$Y�7��jFc##���hyt�MWx
+��<�'���]N�������Ǣ;\��O		�a1������>�V����2:5;7�@�H�L��������e6���__+[�����GǛ$�fݕ0%��}Ӧ�O�r��A$pCG�da�:���[��rnޙ�ʏ\<��nMs�$���K�K�a �Z��I���)��S�=�z7��k9R���#�T5��OϮ�T��r�?
@(���T^3uBs�E!���l$��� ��څ��R{�2�6h��|-������c���Q��v��[/>#�PT�!�{Q���"D��w�SC�u�O�RD(ɸ_��~��!Y�
9������'Q���]�����͹�7���keg��+S� ��������i~��*���(`V@�V�X���w#Gb���NB�SD�@�?"�E�co�\���͸pr�]u�7x�UQ�0H�h� a[W���H�����G�I�h}C���#��,�U�[��I����JP@���G�!�cc�����y��l%��u�>����mD��DO�N�ԅ��>�h�@;���LyQ_굨2��:�"�o�a�|�b�e���c3���0N��[TŬx�Gj���U^�ֿ=�N���Bc�����K�SzgL�lL]�:s�<G�O/��M���W���UD���+s��N"�?���q������Xj�����yA^��WD�rv5�jow��Sb�lY��ڹt{оl�� �b��mIzWKo[!ǪC��:k��7�`U2��q� *k�����v��(�����c���`�<̲ށ���d]�=�Т�N/@T�`q�#�ȹz��2j�B��5�~��.�n��f|�'�����@�<,UG��E���O�2�l8Z3R�q��[Y��p) ���͡��_*f<�xXO=��$���%r*O�m���t�B�����`R#��@���E�0t��>���Ż��2�ӜŖ��݃���=+*����)�S�*L
7!V@xK$C,P��
+�~�.ts�$��m6&�{)gq�+P�ky��n2g��;�=Z}J��g����\x��r���Z�lT.U#�f�C����)�
yn���j�	����T*Jk���5�Z�6M�Hh8��Coɿ�~��-2]��}��5�Rs)9�2����9;r��"��a4\N\�)�a6Db��N:�1@�X��+�����ٙX�o%��:�/��)�ťl���pېc�LvW��s�Z�^�J	p� 3{te���� �"��O���_�a�x�HW�a��~��g�����r�>j�3"� �}Gɔ��j�Hs*��0=��P�wD��ԯ[�(�������ֆ���l����iPc�̥}Xg7fA�k���$e��\ h�Y
F�����?�J��w�#�O���~�l��IA��>�6����|.���E��C�].Բ}O]�"���8��ʶJ���h�>�\uު�q��n2�6�^��f�Js��G�q��k"Y�qQ���
�bh��9[��(�F0�b��7*W���_&o���]�����$�m��	��x��;�{��B��D��Q�uT��s�U��Z����A��� �o#��0�ZD��\T�I��
�EDB�*�_�L���w?W�i�aI{2m�D�P�.��>�6NU�N?�U$j@M��_<�!���V�R�O�}-ȡ{$Pdj�d|ZipY��y:PO�E'�>|�rt�����A��Y�H3B�!o�`*�Ta����K�~�BC��ŹC��P���&V�^���pX����H��$uGD��hC>y�J��2�U�J���V��[��k�l��w�1�	�q�Rۓ�S2
,*zW����~J鞼�ʝ��Б�d�gɄ���sŊ1t]	�-.���:9�4�ȵ��ƌM��M�%��R�{&k�z�9��	�E@��m�K��P��Α_�%aFi>�e�:dg�
�3:�j�aW`�|ڰ���2��ֳU��G���i�����P�w��H�޿�YzR�Z�/�C���N|��"�_1�dD �&��𫡱F8g7��FǪ�w����}�Z�$6�Nc݅�^��:&c�tI�{��%~i��ج���7�R��*t�2FX�?z�5�u��iV�����\��L%w��K +.�[��擽Zub�o�M ��{p��&��"9��X��UW�&I�>97�)�\M�}��	�j�h�q��ueBL�c���2k�|q�X{��5<�	�� ^��HV�W��ws�(R"ߋ�(7�!���Fh�C�.w� -i���v�O��AI�B�����Z���D2���f��������z��H���%����h)�)����� �E���N#'��M�Ώ����Q��S�E9@�	a�s˯�j��j���<�I*OMl�(Y�����=NFI9p᫺DJ�Ć��v�Gj��G�����k�˦�ŗ���%�䌘S��_Z� M�E�"�6�@���h��-�g	��R���f�&�.�OXƁ��1�2���!vB
9�S��u�<3�2c
���߽����@�~�Q�|�W�n����	��=>j�p�8�y�ȸ�R]���K ���z���	�[�OI���_a�<	�f�|�M��ו-,mk32V"�7�^��"�iZ���{�������n+-B}�ڙ��Lu��a���m[�fZ��S�����7�k��qэgm����+C��ߵ5�p�y?���d|�a���y����ȑD ޮ� �6h��g��!���{�.�o ��}SJFhzHz(P��Ǆ���h(M�y�:u�7z�@ף��
�	�psl #�AvJ�y�����|3�!My�v�$��e�� 9>�p����>/������Yun"��[Db΀�R�ĥ��cFük��n�~;�i�Y=�E���M�췓,}�0x�kR0� k�na�����{��������
6=���y)�g����R?(Yۿ�V�S\�&{��0XE�SN��eX��\��RO��j��h�[~��S�Ḳ���Ԡlh3*=��+A�5��O4���P�Ath�� pZ�n�m�;��X=|w�	���N���%�zX6�!�G�7v'mv�Mf���9x.�8闸��e|Ie4P0�� u��˺ȟ���8%=��d���ۂ4��7!>��ueO����B^W� �Y����P(���=�*���Y[�(TI>�mTJ���6+ڱ�1S��q�>sg)A(A?�G���C��׸W}eN�l���ah�kn��z��8��~;d��}�84�P�9�h4]Gf�[h9�XY��R��\��*��"����9�Pc,$�"��LP}���y��y��Spx�f�NY�*�Q���S�r��Fo�GL[I�`�y�zW�X|Sum�^V{�Z�q
]��Yg�x?%6s��Ҙ��.��C��\��O��BE9sT)��O�.�C4���p��K{�m�%��ʺ�@�&͋q�9�H��Z!�����N6:���쩍��<�G���y\�g�qmK�m��j���n7{Q���i$Ш�m��y$���q���i�OU9L�±�ao����|_��F�^?�v��ɂJ�����A�h�b����-b��g1���f���iT#�2��}�fԬ�Ã��� ���&�#�`=@R�>6��d��	@����-�.X�xcqo�ՌD��
Xu�.l����ڦ�.��O>zr�T��ó� ܰx���p�QV��dqf�6�>]�#�쐹s<$+K=qdQ\�jz�J�nv)�2V��'���Oo�q�L��� wk���$��h`P�~�@3�dw�;YnG׆��G��	��8[o3�ڛV��U�z>���'��uV�YV";�<��Qad��D�I��/���[�6����n�:����[I�5g�#-��+AߵE��9�!۔��$7#�!��/����,�^bi���t�W:ȝ������sޝ"��w�ӨXKz�|�!�ᠥ�.�A�g�'�O�K $�/=֕T+W�"`��UuuR�{��L*�]�t�KK���US�$��?,3�s�:rqqm�)�SE�X��y��(4G�v�S���YH�T��(w��Z��DW&�I�
S'{m�օ��\0�ܸ�EIL\�_)R��뒝\Em�y�X�j�Fnht�x!��ɂ>+�C�f��-Xh�d�P��㳯Z�	5�	��Yb�B?a�z�w�&0������I���)^8Q��� l�g���)�g�f�w�+���ۓD`VYUu_@n�wX?�z�`-=w{
Yy3�fbm�c���vӆ4�������Ez�vv��]�c��.�@[n[���>r箙0��dsA�����0S#N7�42F_㩕'��N�,v��o���2�a3u���Z������Si��q�9��+nM�C$4�JLI$=!��׌m�B)��BIn�z"_�nl$��	S���Dc���n.Z
�'s^<���BɆv�+zy���*Ԍ pw˧�@_.ɨˌw�3�>���a���!�J���NOgp�rUZAn~%�����:�y���u�^
7'K8,ਛ��1�l�N�W
��r ��l��&cb�}4�0��_�ĵ��������E ��;��~���`3���Ř��D_W� �QJ���t��/�޷$}4���u��~�R��� 㫞�{`&��F�#���`>���_�a:,�B�e�XyW:K�WppЄ��9��	���s�9�,X|�L@C��XD��� �Yb��08��u;���v@�F�,]^= ���p�k��#kl��d[� ��=�� ��)G6��@�I��$Y��w�T���Z�P	��]/+$)�A�q(�/}�x�^9�X�'\.!�J���Z����vt�,s����Sb�oV�轶��G{Px�l�0 D~���P�=;[��?_�T���F��Jh��Y#�;eIT��$S�����c�����b��`'�řւĢ��:j�X��X��oK��o���*�iީ�Q#�T�0��ǈ�tF�V���V�@���,9� sr���o��tn�,+����#� �0��(�=�3��Į��k�lȷ�M�qwҢ��=���ҼSO?<��ݹ\��|AorI2�T0�ݮ�w�l����(-'��&���e�E�#��J�,��A���2�ճ�(�1�����ʧ��Y��uL�]�%��h2�r�LC{�>A&9 o�{e���D��JPO��P�-����78Pa�|�A�� ?d����ѽq���;��*�Jշ42�t�
;��h}0��H��Y�kl���L3��֧v��0=.�2|���yz7��Z����~:ا/�&�D"������.���V����
Ir94��R?�\�S���4�r�G�	��$7|
6������T+L�]nU�#�JA����W��d�b�n��D�DEE}��6.YZ��T�ǌӲ�K�oɩ������4P>��L��EQa#/d1�� )d3L�NK�*�����^ױN��dE�Zl�v=a�Y�~���/R��F��Dr]g���>7٪��9<���ƂXXx,:9F|���@gO�J"����ۢw��쨰�c�D�DZ%9�`�G���|<0���8���j8�`�؏'��5s�L�iC�t8*��]Iq�_T�JWá�:=W�����~Q�s�7�<��B�,�bE��p3nh���D�:A3m�ke�nw2�J;�	.\�	���^H�gdUჄ��ڠ�{��[�L������3
2���Dt��]"��O���jCb�Y���P}}iR>��ɘ�x*&�<(��w��:+��)���RjC#��恝���Y��9����<�M_��b������u~��0
p�� �X<�-��ٚA4P�6��,��K�~��!���$����j�LF�6.�b����9�V�I�k�?.(�v�l�9p�B5>V�M��>8DO�ϻ$$��q�5/�)��DfY�X�$&�/�����؜A����sZb61�Ff�����,m��DhíM�݌����zQnP���Jmt��v�jq�`�d��퐙
�4۩�k���]��A�h%U.�*S�3�̅��FF���⿦�x�n�4�Ǥ�/���09I=$�-���ot4Nh�Z!�%�	�䄧s�V�9pb�s�(OT/�^
�ѪzH�hY�{)#Ҝ&f��r�E�E�>Ň�fqM0�a�/��۶j4\�]��yb�| �wX�?W��r$.���z_�/ե��>��VT���-\��+��)� �szx���C�Om6�<F����,d�8>�$u�]�)�R0�d�ǯ�70�5Þ
�_N���ٗY���p�Our��,8˒V)A
螯p'�g��ܺ�]31j�ń�&��;�Rl8�:8��a:��)�_;#����N�9��f��A)�
a��y�޻���i�'�2���['@xE�[�� b/���j�M��!K�Fc�g�M##��17�W���c��fD�xc�
�ѧ&7ƽt�ϛЬn��fċ�{���"��Hg@�,&�{�z7$S$��Te�j�C~^�Eu�Od����02������G��e��uZ�-m2�}����3`"�@f���d�e�nf��Έ�#�$^/R�^�O3˟���' �tέu�	��.g	�4�)�5c|U���~����mh2u�8��\P��W��h��_�D��rJ��C�ʕ����q���i�*��nְ�
1�}E�|��B�Þ�
!S����cC��L+p�Pqq�g4@V�����T/p���9Iϴ������\�u`d��W�6$�n.��4�V|s��+2��o�\e|�7�G�ų��;x�J\�$� o(���#�G�!P��B�N��C- �|<[�J�Z���<�ҡn%���Ҽ���-�:�=[)�~�Ѧ�c���S��}��~�H2�Xs�����ʠ�"��0]�OrG&ٚ#�[��\��Gݪ)�����[y��$�����>Es7�9�:Ñ:�$��r�N�f*ff7<b�΃L!
���A�N�����G$h��a�,A3��6Xf�,����fC]�n){7�[�Ҏ ��	0��L��d��Cj$��R���KXMl�
���
�"%m���y�u�Z����p�Ȓ�43}O�T$�x��+E�c/��\�>��H�i+�P�$��S=i[���臠vWr�Z��T��� ����y��rNC����{���γ�\����%�k�������pfO��̒wSq����0�K�}y� a��g�C������Tr�%�0/�bd�ztT/X�Q�X#�|�>%^�G��J)�ME�p���x��=*k��U��ö��S��}0��p�%���8͂����=-;�ݾrt%��E��QP���ٞch�Y���K��<(oT��,�����J2�A��`?�ņ�h�ܑթde���Y��LW��q@6��	�/l.?���!L�p"ە�у��
�/�g�|)~�+L?�W�G��eQ���p4Ix�L��ݘ[ݪ��ң�Q+˧�
�`ԃ>�4N���ZK���������i�۬o��r������ϯ�qr������r�[k  g���Y�sf���W�>U����Mc��^f�ͻZ#{+�1>��T����7m��;��Zֲɍ���#��Jʲ��Y��8f��S���9	h;4�e��C�Vl�*N$� �� ��s�w�_N�	��'ԷI��FTk*�g�sP�1r�q�x��^M�:"д��l�<��I� _%����V�cFS	Uo�����&܊�avlv�W��?I�f7>,�A���_�p��NQ��C��xa$d�C�XJ���A��&�įB%``a���=jH�y�n
<J��a��A=��y��H0Ľ��j{%d�3�e����Q���h�4u� xH������5��H8rF��&�-TԺ�Ϸ��k�cM��y����"g�X�xN��L0P�(�ɣD��������w��`��-�����kOM�c^�O�jQԇs���;Ӗ6�9�@y�(��99m4v�[��F~|���i��,�T��9�Y�;ҴX��.���6m*�%��:u2�KN�h�泯r�$�8��˗��<Z��(��>.xӔ����k׻�!�D���˓@�%v��F��f�"2Ǘ��sc�A��`�����b��F	�zS[�l�*#���W9C�YA|1񅖝�/+�+�e���N{�p6����3�1�W�f]���곥t�Ҍ��J'F��@�8tT��_��Tw�g�8~j��v6��U��lo�1|��k��Τ_������˘f��LY���κZ��A�976��Y��G��:%��q���.��'w���� =��kQ}�jjB�3����'�P?5����H�����0�'<=£����Fa���gΐ�fi������ޱ��H���%�`�d|��	������R�����t\����xU ^�����Ј����ʼ8��M�MY�azwFi-b'?��$sk[L�3h��a�2�WgP}�e+2�8���_��jMBTQ�'m٣<��ԢOp��k]�=#�&�.�.��|�#�X�Suـ46F݌	
4٧� 5�G�y��i@�tn��y�)�GO*�}UaƘ`��&�EЇ���t��&f�t5�<���zi���\��N1_a{~	\����(�p�*;9F�����1���f"ǡ'������<���?#��p�����}n�:��г���OSZ�"	�;>e��D�~�#��D���ر� �ʛXᤏ�On�9��\M�}L�C��J,���?�񽃘�J�͍�����>�������w�?՞�po�q��p��4��cߤ5�p����']�K����Q:�6�޹���A޾1Y���V�P]�iB�21J6i��}*��~K�B��z�z<>t����`o�krzfT�w��MN|��P�<�&��[
��- ��M�p�ׯ3��}�A���ꇷ�**"[�K�h>"�O�Pk|�K�_�,�Z����'�N�퓡y�����i��BW��9Ґ�#���I�;:�9Ex��5~�æ���3z�$d?��(��`mia!mSδ��q�L��CC��Y��l����U���έ��+��x��N�=��~@�K�X9Kh����e�����q>�2%��9�/����������L�������O�W���7{{�p�S���Du��w^��SSW�mey~��az�tx������9",:(7j4����>���R�ZXA�N�vlx�����V��Ĉz&�5q?#X�����nS���ô����48���[�� ү���'jS�=C��A��N�<h�љ^z�Ŝ�z'Z�-G�H�8U��p�	ܢJ�
���%��i@���4�2�|>���qx���b#7�Յн�ԑ�o=F��i�}��&O@������py�HP�0���@�UX�#�'fЕ����L��.���ϲ��܊�\K��kn��	.�
��!�N����.����<�)^|�0<�Ⱥ�ױ���ln	-����V��"�H�FYq+�}��a�0%Y�jJ��U��C�A�tA�t5��}7��b[Q���	��@�N�����l�Ģ��wթ4j���x�pU}C�꣸��ŋ6���_z��$כ;�Q��/&E
�d���? c+���ȫ·��6�ƮkC�K�_9~����!���@]�i����]����V3=D�����h��#��/J�q�k��`��f>��	�e��̮lBO����y�ogԆd��0/���u+�u�@�j$&B'�>"����a��r�2���E��kyB�eJdi�xvO��u}�Y�'��+�/}ׅ���:%w1
it�rD��B�Ž�U�!�������i��ޤ,����UZ#�DuS�ߜ�S�	D2O	��'����F�����~z(�=Q�����w�=v7�%=�X
�Ju�E�a+@�'2;lT��������������9�C���3R�K[X��.}1����0����wǷ� Ʋ���^ &��͚��K�d�!ґi�1��IgX�J͂)�ڹ��RG`�s��P���D
}5T��=�dN��菧qmN�^w�u3/:5O�3�;�B�rc�Ok�/�Ku�ʵ������K���NFpF��-;��!/��tղv�6}��{}D}\#��_uL0���Vlu)��RN��\��
Ui��j
�<���*���Z8��i�J{�*{B֓dt5j:zf�2�A,�g��(خ��K����t�*"�)�[���u���z�O$�۶_#�vPj⎩� I��y���/��O]=��{�o.���k��W%IF�idy���Z�G��F*'U�S���'DY��HzX=��z��7��5�+�UI��d���������n81VS����]u��I�ؔ'1�\a�B-��1���⁡$�������5wM���վ�&Ӗ�b�F�B�����0������?k��F~[���̀�����x�����yX��.�B1)?_�q���z��B�������X�D/�~����>X���4��8ͽh���y�����&g}��6k����+f��*�2_�XL��8�
zHG�chȢ~���%��ݙ1f���i�	F���7�JO�ǎ���|�M��mhm��N��᫜�3�z�)օo:=�(���)B�P�R?�w�њy��!���f�r3~���6��T��`v-F�� �T/�t2�e����Ú��ܚ	]Rl�r��"�q�#���
������Iim�3��w.>���#@2&&��{	�#�\�7�k�sc�Y���6�,a�	����B���j������o�'N�<݅�[����s/F����g+! C���8<N�.tE�g�}�*������bܾ��_wf?�4�P���� d�I(rsҊ:O{��,Vf�m�1�5�r3o`f>��ip���sna�"|��._��)H�%XA���zJ[�̕��#��Ҹ��9!�UV�9��噦�i�"Oz��OHˊ�Z���NS�;Oj��e�F�,N���
Nb[�F��֫�L��F>�x����Xd�J]�8�\ިk��j�*Vz�����R<{WL{�ZF9��u�ɢ
��"��B]�]��8Ǔ6�r�����3��5�B�qoN�	�}DN�ĘZ�u>�=�&�S��.�T�3�s�Ty���/zmI�˸�hi@� ��0�AR�ql��?-w��o\�o��Ac��wm�!bθ4(3���M	��4�3ť�5�m-T�^� ����̉C	҂�|p��$J���q�Β�
?�a\��6�g2��(6$sH'�| �9t�'f+a�MH����S�e��@��gk�C ����K�����e��jewh2��~�c �.�>�l��|p�nZ�����֟Sf�|u܀��Cb�ߍ��I�nQ1���C�n���*�[��f%�l	i׎.9V*���%K�����I�J��*G�6J��5.*2^?�-ֳ(ڒH�B�/h�.��#Q �8��q��ԦoaO�c�~=nA�0ؙѳ��.5p�,��7�D���OD����9b���ՠ�-���@ԙw'-�ܯ�Ϟ�����S�46�Z#�"9��à�8���V��2�3�Lj�m��`�m{J>�v���d�O;T#�y���5�"ZԿ��]�%O���f���}�qC�v3<��p����F븖�\�l �-)�ᆿ��
�ܭ���̕"��.i?�GRD���&�E����g�r�>�����m}��
����ȏЕ��Y���LiX��8�m'�� ʙ��,K k?�|S����V�o�t*�W�R͒�8Dn�����M!�!wUv�8%��2?@Yڻ����o���jD"��a�-T=nk��?��@CǇ����"$;(�!��\��^D�KK����5Ζ���N��*�m���Ғa��[�O����J��9�ۋQmϲ��H��Wr>E�W���$�o�G#�/�6LŔd�7���D�m�炻��~�Ӭv� -����^�Ϧ�W�\�G���o�WV:'A ~����6<m��� Zc?�gc�JԖu"p���|���$p�un��̬f���)-�h7���e��/��83C�Ep[�H���0Z&IVlo��� ����2;@��`)]�;\k��e$x4R�.��s����Q��@�G�'���a.�����X��ЋH�a�틩1@�!�Zk� ����{d.\�aAV�`3aT(3v���~&�0���3'��uM�5[���B{(^�r%�5E�Z�����h����]�0U�A�2��Q���#|���h�~\�1Ex>m�m���?�����hG�����y�8|���X4��tl��3P�Ɵ�����a��m.F��I�����Fi�t�� ��A-ۮ�2b
ђ���7�}rD�Z�-���
<ͺD�X�Co�8Ĉ�.-Z�'�����' ��"��)�iY$ҧ��x�B��#�N{�%)NƓ������SND|k�n%er)Wr����or!���T@�K݃����ʞy�d�'N�/V�@g��;����$Ԧ �#CKrab��%�����`[r+���>ܮB�����.T8�{$dl�.iC��ǩ=��}����Mb>�Y�dG.���(��v�+�ı��G�[+��kf�)�y֕Vt��]�滽q�x8���`-/��;��$3�K���"Ù��4�$Z���Xs*���?���I�7@�qV�&�����H�$��R�����lQ�KrB&[��Jg��IW
9���nKs�ˁ`I�~��8�S���l4�������b��䍕�c�U}�ԋ	���E4�%zi���}�����@>Ck̔���rm���k>b��,~Oi��M�o���cy1�gG��g�E�(>-G���˓�P� �nP��X��G+��s�A,�p��4�D��UU-"�jt*� *V��љ�N�^0��c��%���/L��C�M����oB��J�@E�� �m�T0�&ԥ�ip,y��I��u7�~?�=MJ/�jý��-�pߤ�=��HL/�{������7��(1mN������a�;7�Tt��a�joƸ݁�!�dA�\��o�z��?zG�p��� �i6����K�B\?'SIK���P��wf�+f��yLS� ZP���kT��T� F)-�=���_ɾ���w�>1,M�m���z��������B�B~&�:#�cM+G��?�������@��1-�t���aYć�=�������ό�����R�ʤ��e^C���6�"���aEDF:��%�}�p��X��ȜAly�I��3`9����n=�2vjr�m��Ƴ֬y�b[���)M�ؗe"��Փ�#^��^�����%��K��6�Tp�Z�Fʄ�4u��i��Kc�������FB��-�S��ݤ���	Hta�'Y7L��U�r�^��S�b�G`����sEѕ'�TK0^��9�$ƌ�����?5fB7�co8у '>�}c�"��QTnv�w�����](UZ�7��&���1ZR����A�{Q��5���vג9��q�Ux2)aZӂ/ ��{,z�@ۨ
����X��$�;J��"
=
2���1���P����\���X��2�nV��\��X�jxFfl��O0�]��hH(�T�<2}j�nQ�u��Y�F�v��
��� �r�n�h�U;�v�go�q�|��z�p4y����@�p�8#,D�������p�ꮙK���=�>���RNu����>�
tW�^�N����I=wz���BU5ODܰ�IOV�a	���UgD�;67S�#�5k*eK��(%�� GǶb��mFL�A��G�#Z���V*kr%Mh��$� �>T4��D���w.��O��x����:7=��=i�k�i�f-c>+;n?�v8��V�=�=��B��Y0�<�GCSF���A��5��"ܶo�W�@۲'���칖h������*[6�1�AGm�Y$ݳBb� ��h���Ќ�~�uk�"W���Hʒ0���z��Ns���,_�3wG���Kc��BS ���p3MU�*-�pɜ�-1�ې�E3�Șz�W��]�K��/@���T�
E��{��2�dL;ӕ�^�ܠ^���gA�Q�¯���f`��	o���V��}+�ɡ>�U~��M�&:��.fփ�F�l�Q������}F�o<A�RRW��5&q�.�����CE�N�I��y���tb�Q{������<��C$�&���p,q�������<���q����}8�=��Q0� �D�\ɶ	!�1�$}�OSQ?��J���85=���C��T�=��b�|����XE9�QH�C����=m_*Q�u��{)�*s�C��%��^[��{`I8?c����9�,��:78䕆R�;�Y��"=�{W��� t��{⟚\Y���q��ƨ�G�~�I��"'G�p�{|Ւ��i��{��F��7g�� �uV���JBa���4��čy]uvx��I8vd6�gч:���2}�L��e6HdJ@��Q�!ARD�1�d���`����D�
�3�#��m���<1="�e]�r^�뜻zD�
VK���=m�;�2�A[�έ(3���陖\�Z�3�-���b��>rM��9}�rz3�]��`ߜ��;7]�N����Q�>����<�-�4f˪ZO�F4nr2N�ˮ�~f�����Zi8�-�P�[�P�V^���ʯm�7��&��� ۜ�+ �w9\\_<k�.��^���x{-c���v�پn�������PZBM�f"
�?$�@���6���0H?zD���˖*EF��Mb?qJ��(ȥ��ޓr��9�a������b��n��X�1��0kI��9�%��_W*�7.�&ݾ�W�,�\����qa
���CCr�y�}�>�UL��Q�g ��.���<1pY���M'����8�F �K��\%J:E�h���]߸��s��!�Y�B��_W�-����5'�M $��i�>�Q��!���Q+������$��쓸��XQ���wU����ҁN��I���+�������U��N�?���r�� ��SP>Fg3<%����_���}�(�ggH3J#.B�Y�HJ��P�PP91�?I�t<�To<�T�l��k:W݀���Y��) �+��z�옔�/>�n���"�dә�Sw$��A=�=�@[rL˰Q�D.�?�ę^9�=�e�+��M�Q��� �8��/�6 i1H(���Pv�S'��\��{�0�sY�Tt���)f$i�>/�]�7d���и�����a1���]Y�i��-���s_ƬS$��)]�B?���fs�B�o��1��|t �P��K�Cjg<�ŧG��s�K�d��ڒ� gW��b�켏!
Ť[㜤q�]�����8� ��n��Lr��} yԊ�q�Ǒ�qM����+����k?�95l�/n"p�~�]�ji���!���'=�<>��Л��ho6ω�2�j���W+J�����ٿ������%|!� J���	o����j���fh�%U��[ N&8��k�^�
Df�y��M�e�=G/T@::F�Xw9OCg=O���R�������υ�j:m��kt�Tm�_�A: �8:��Z��H�Q�ŵ�5:���GK�]_j�'���t���a�j��=첀�cW�pQSm�9x	a�jN��胠3@�1��'�f-�D���ke�]�n�ٿB���פ��한;���/�+B7�z埈ߚ�9�;�
ؿW>1u3-2����C�� �S���C�b.y��B���F�S~sC��0\�q,�b�ٚ�:s�}�q����V,	�4Ai� 1���ꜜ���,t&P����U uWaI�EK҂��2C�9帄\q�t��ʌ�C��\g.��D'Nń�m|G�Hʞ�8G�߯�W��̖�h����Et�����3�1���C����tl�,x�̜�V��0��~�^�d�>0��ұbD�{���>�19h�����~�K�K������a��]����`u���ž�yi�uJ�ߑ��7u�|�FE? ���7�mj�3�ᑝXҒ$;�L�w騬a�&�Kf�Xf˝�r�kK��5����^����b�����<�!�+�^��&�c6�+��%C�Q[����>Jσãҙz7��o�~��N/8@P(��ZŬ#��'���B��E��<Xr�H�<��U1gc�<H,8w`ҁeoH(�%
9ϑA��E?��d���9Xv�Gq-��nHv�q�n�C�.��M���O��>��m@��l/Ű^���M�\LMA�)��Jf���&a�;��y���X�3\!�Su����Q�8	j.m+ZQ=��.++�}����D�E����'�߾���F[����_$�����U ���?a7�e�Ҵs�(���s2'h�uw�D^�:�)A��U{6��e�.�	�<��=3b�k'�G��M����$z0b����ʬo$�[�6���/:3T�E6<�o��VoA�7�[V�
�2 _�_��ZP߬@ l��$�aP%���Np
{9��VV.�TD��M���<�]�6��v�fqg�����W�-7�C���w(��k4C����&)����k�p�X�i�Gh�,c�x�q�����Fʔн ����\5�zr�AԔX�.��s8!�g!3Lg��Qf��I��@
#]�L����a�&/r/ᨙ���y�-NgZrbo&%���^q#�LW�ol+M�X�э��G�N�A��?FN��^g\�f���A��
������7ڣ�x�7?*O����*4ڽR6�-"t ��N;<a�W���nsq$f:��?~��>�<R��2̤��O���9�C����A�z�!KBIY�D@>ϟ��tb��-o�*���F(*��~�:O�,	�OQ�M�acge/�^��BMH���+ؿ�C��TH� ���7j�=Mlj4���k��gw4v��Ꮂ�@j%�>��Q���980Yv��zV�
��`���\;���<�z�_K\^;�"^ߗc�� �B��6�N�N��� EŢg�g�tݔ�X���G�]�U����Ox���q��u�G�+�k�?@�fz��s�ݐy)� c��O��H7�dP���Bq��:?�<��J=#�E��P�,4���ٽ�]ߏ��_J��A���?����9-�o��<��tBY̵f�;�#s�k��2x%�C����	z$j_�E�S�K�*1;J	�wї�K>
R��Vp��H�������1�B�B$��{g�ԇ���&����iQvSF>>��j��������ڐ�'�k������`=�fU����υ}A{;�6��������|��w��
O@�"���?�UE�I�����Q��PP/ܬ+��,�qN�yTL�|���jI�j���Pݻ�����-�k��-:��s�W���w�<�qqL��O�B�<tm1���$D�,.v]o�M�����s\Y�I�J�&�*�y��k����P?"o�i���F'Sޘ�Vt&;�����>�i�4o�*g�j��	�84�3��#����Pb�c�7�3�����iL���G�ZiZiӌ���a/7��w\�eaQ��~O��Jv����e\U�G���Hh�S�z�����T����G�S��B�-�'����^rۺ�<�2pZ���s��~�h��Y]7g/+:�8,��a�z��b�v�^?mA|c�d���1����c�����1?�,uAS"�n��fO��h�^�AO�cMTX��9pNY��� ���MI�'<�n�[��~ZC��J�u���t9H�Z��=��9�1Q��H	��C;cQ������=�0��hU��G��|Zկ�bK�.m�SM>ᆲ�1^�¶d7��~�[�Ɩc�ɗH�IZr����{tWBR�/����#�_J�N�<K;��Tt����.d?��﫺W���ύ6:���?L28\}��Ջ~�~�m�0���{
�{S����œ�l|�R��Yӯ���[v�j�U��"ch�L�}
͉��������u`����2m'F��s����6.Ϟ�[Yh�Ş�}QZ�{��5���4=W��8���8����
4���Y�3GC��9��r&�{�7��<{@��8�q*��F�H�!*J�D��Z� �;6U6ɭ����X�0�v���������W|6���I۽��r�'x;��!8;�����Zي�bg�[�J*����䀧���;��l|�Gэ����Or�A UE�,)A��p� �Ѽ#�0�Q�)�n.���h?�#W�Zw���S#�
D!I
�t�9�k��+�L��@y��ީ6xR�d���Zz�+�b��Hf�p�Y�N+�H6���#I{X��3!i�uȎy���VO������B�}�����"��Q *.7V&�>��Q®$/��$���}�V]x��V���LB��;�����Q	n!J��anܙFNAű1�9�?��I���4��J�a���3�����z|Z�ǮWK6L����=��oò�ă���b)���Yn�����nXF�9q�Kyf��8�Ǒ��k�B��_b(%�РXWA��w��d�6�J:4$�,i��僳�=m��W_j����*��N3Sp�U{Ň�_��E	<��^�J��C�`��{3y�t�ۓ�[��D bŪ�3��;S����ޣ*o���B"��`�.ß��`��r?r�)��R��Aۛ�}:�J`��&�@�t��ib�<���z�3Fy'	��"������m`3��.Q�^r��t��Z3�sݢ���s�&L�ϧ�UF,^�����n:��T���@Њ�b�[맠�ဪ]���\2��.���7�
�Ըm�n�]3�y�[���u#U*�ٷ歛�kSz��=8��0��0x��M�|KB�-$�ϸx�WO�p�hzO��x��O��$3|�,>�h������,�����ذ�b�L�c4�i�K������D[�m{�Nf��SOru[_#npQ��/	�|ٙ*k7����-~1�;����g��k��1�Wt����n�2A��;}���wWJ��61�">�:�M7e��Z|,�@~��ң��S��^�:(0�C�	�}yBC��k]��-;s! ook{@ �?�yc��:H��V�r�K�w<�$�G9'0֛.��zٞ��P�<jQX�;g0Gz��BFi7�m=G标�/��,?��!�ؐ��v��Ӡ�6G����V!h_4Z.��rO��>"2{`u�$�l�W�kЕ���<�"�(�wM$=�����ݭƊ�@��+������%��4�=U��c`���T?NO�~YxP�s�9w���SO���k$5>u{����;�i��&��b�����J!�Fe��EBӪ�����,}g��ac�=��^�5��J0���)(Gf4`O=���.o'��[�<)���Z�`f� kØ�G�*v����<�2�m�P�/���I������ЁeQ��In�[�p�]��<��e<#"��������*Út�����8u)><��'3J"^_�9t����Kw⁒~���&C�{�2�R�ѵ�.�!2�P��	h�f�B����nYָٽ=~nH��C�̃���A��+�x���	��)I���t�q:7H��f�S/NB�Q����B�ջ��nд8(^s03�e���I�w��!��Ha�V����W��=û@9���_&2�0�־�S͡ɑ	�!p��7��F�C����� ���Ҳ��J�
-��?x�u%���C�|a������/�J�Eczo�q����3�����{inK����Y\���߀�ľd6�g]5W�cM<5�R���N܉|6*�J�,RN�-���Ԩ�0������yF*��ly����m��Ǹ�J}ڧw�M;G�r�E44	ry��*�u��#��Nzc�W�*�*A�A��lf�d"�Lr�I�`�h����"���V�������~rev~xԸ�,Dmd�;����=��?ٰo$�2d0��H�e#�b�n��ɍ7l�M�Na��j��Z>��_�+v�c��P�Ql9Y)�B$��%��FT<���_)�����R��V�l��&���<�߮���6QK�%݇N��I���gQh��� ;-G���pIE�딪�i�k
��~���,p���-I��ށ��zh�c�����m>��]FnZx�Kܗ�!~m��K����H"{SM�[����*�W;m����I��i���*L��U8���/c��0[������L�% ��vٰ�]��]���m�GG�q��l^��;(%��1F��-;�3IQ������	q���5+��:u�����ϫ��T�� ���g ���\���=������x�4�2}�z�u;�|�՟�1�NL�.�E�O]8�!��8�H���K[�[ B�z�h	Q��Y�yE�L�H�/��B"7מx{1�O�r����?����L_�I?��G�Cr3��}	����Q>v$w�%�Q[ILU����E�*��p��sM�e?�{K|И.%B�	U�v���&c1�Q�߈�$b��ت�������M�?�o�cqo��u�c�g`�W�Ȱ�G�f�h���F�Z �E9&{�4n�g�Z�w��\8}�~�d�sMn�!��v��P��o"W����3���%�����Bv}�c��*��a6�a׌O���
\n.��hP:bz�	��K<g��ƹy7K�#�.R����"Ӯym\�y^Q�*��;l���v��5a��>�[Ԉ�x��Io�+WU�T��h���#o��,~��M-[���Ѝ���E�2�$�z���hY�z�Z�U����o���_�)GJ�����N�'�-l�j����ݬJ��Y�*� */mmぇ�SpHHT����Ȭ�4>��=��:;��՗��YĨ�.i0������EH�ٹ圠	�_��Ym�ro1���Bh�*��h�
_�]���A
A� ��c&~���e�(�;-����}pTt�<؄���i������^��a#ݿ�i_�x���b�q?��[�^��kW��il��M����YAt*r�燓q7<|�i%Ahrqסl'nvT�ɣPd2R�<.��M"RP��{®s�䈬��"���/Ջ�X����1�%�pC�t�Jdf�h�a!L�Z�'����9؜�Y�Y+��ܺ�o�����7ql�5��f�eiS��9����z{�7=��韴x�s�(��=Mg�B�������N YU���R�u�;'� ��f�WY�'r͞V/B�N�񕗸L��m���=4|��Y^�N2"��Ɋ�����ߍ��ob®ӟ��:k���Z�g�-#ʅp	�ד���o"���Q��:?.b}-�suҗ�BѢ'����-C7.R�]�� ˀ��pV���u������=�X����8�\��@����[���A�&�^�\4���!��  `BMMZ�K����oN?��G09����zn�OA߭�i��l��r;�ؑ���F��*������Y�YK����M�TU���ў�T��;q��`a;s���h�iȂ���%uL��W�&&�v�VC�[�a`G2���xQ�[��'P~n��Q	t�(�<��M���X:�09t�0m���iu�Z��6A�8��b��]b�����7i��Ӫ���+'��A�ua�H���ya���K��&���-?�	pf�I�ٺ�A���T��0�N�2k����-�:�F��v�/Vh���X�����s�<����ӓ?�`��@��ƈ��Uh��}$��AME��X4���,���/ϒĀ�	@U|��lf�1��*s(�o
�ʨϺ��f�N�����nv��̂����+k8�z��o��9���Ȟ���EE�^:�l�ϩ%9��Su��->w�%;s��j��[��Z��i_�-}��&��Qh�ܔ<���x��RjȖ��(5E��~���$i�;TP�z.U Qal�ܖ]���&p��]��zOL$^������ o\3`�^CXu_e)��Zei����̴?#qY�����&u�3A峐w�h[�~U{�F�O� ��0%ɡ㛚�Č�U�����&�Q������/�z''$��	�H�U��5�>K>Зo�W���`9�S�s�D�-�r�I[��Wۺ|�I��4���L��Z��,����\J�/G��U�wx$T`Ԉ�B&���d�-I�F��B*E�i�3{��">��Ph�\�ze� g0��%�w��L�'� �^��<�e�rk�??*x���@�M��ϔ<��+���
�ɲrT��5�P��@��l���"�f�P��T5#��@�S {w4�����i���|V��n
yy���N�$�\P]tFK-��d.oLʂ������K���'�f�W����;��\���w�&9R��eێ+�f����kp�w����F��$3ᩨ^�ۥesH�aW!R���� 6uߠ�����e�v��\>ZJ�������H��#ŵ3�~&�T���6E� AFA��z<�Y@~(���8$(��7�Uu7� ���׾Cy��@�ر�r& \?w7���F���k��x�O*���NRl|���W�żǓ�0Ə�C����t�\��]NA�q�#�B�zLEĎϑ
�%�5q��E��-D�T���4�; #N5̎8p=)2�/��a��H�1���6󗌿X������-����:�;�b��W��a�˾"��SO۽��c&׻~����$5ۚM}���π?��߳�����^H�#��RqW��У-���(��y��%̫���CE�9�>+e�_ ���=� �]m�g� ��Bה��pa:�=�T����Hx���@H��`帀7��ۅ3��,�h�o}�,��uܪ�����1ý�0�-B�]��<�QC�7#��v�'o�բ�n�)�����o+ֶP��]�<���B�K��9�{�W����o���x�%+��[8�\$��=@�����g%��1�%�k���aЬ��=����U�{-2����m��$�.`��q3��A��-Q�"�n-�p��|�,!��,�&}f{׈�*kP:Ϡ�� ��@"�=U����EK�M�'�饛=��ܜ�E%(=�����&h�M-�j���E[.H,�w�7���������@|��8��Q>x|����Q;�;��j<�7�OB'��ӆu�B�UG��;aǘ�'�P0*�D��\�*`�KI*��}�Ģ�ӺjS(���,$�,�ɥ޲��MR�J{��b����Γv���^G]2�0�u���Bw�Z�M���a�d��b�fז�\��5n�_1���MA�z��+� zsn�5��wx�{4]��*ȑ�խ��U�ҿd?����D������.1z4��yԭ�5� 9SSB��O9�5Q$�������)٬i0OH���TR��$_�ޥ�<��~�e��)�l���o�g:��YQ�$G�`oH��i����K]��*Yo����mh��A���u�����[|睴��<a(=�u��P�̰�ᄡV7��,��n�9_?�dd��:8\��� �"àZZT�-�"��������������͕�o�d�ez����嘎����tи�E)�e��J����}`����R��s�MOє�ֈv��4O�eA]�Ʈ{K�o̰��<!E"��f��	u����W�L^{��@܅Lέ`��&t{��~����1���=��TR���i~J�^F�O7Gn��2�����ZLǗ��X�|a��<���L$��k�V�%O�VntEyB<k�B��������ay%���M�P� :FЗ�fJM|���<�C�?6�;���]�9:�j ?����9���3�\ɰ��ŷ�vs�h� Q������*@ox�g���;�q.!���{�=
��ǩ��\�o�����Xcʑ&քx��AHG���	��5yT���~���r;����!FE�K��{���������KV�:ÛN_���(�2�؜��*RU:�U���˸%���b��q�r<cN["�=��������� ���Ōp���_����=�+�)Ⱥ�Z��K�����ky��$W�ڶyɝ�_�8c�+S�0��J��1t��'D�C�u����J��jde��}��$�f]�:8��&��r;����-�)����2 �wK�C]*�Z�o ��2����,t	}X,񼛻	r�\�c!H��v#��\�n���C��Z��"�!_�5��ۨ�� NDc&Y���z��}0�)�%�q���f�5�j}�\$z�j�?g����9L����F*��`�ns:z�m2���Tw�ϐ��L�2����#�!�*�ӄ'!�"Q��S2��������Wn!P����k�yd#'b�]E�XљR�6����(�5@�Q�+y��[�,�Dk�TF��K*���S�����I��(�Ɏg�?lD�[�H�6��%�\q4�D�0���hŖ�,p�V�d T��0ʵ2��o��a�"���!&��g�&"3�zҩh�$��og�|�vB��f�a�+VO)�Ɨ�*�� �תC
 Ȯ�N�M�#�k0���:�+�Q���.��|֦���bzB�D��ւ=)���RO?�[�#���6�ը�] ���K/��R�b-������w
��&<h�ey}�Z��}�l�c��W�{�z�zJ��a�ϵ�Sp��B���V)cbt�΢_�(��N�����؁�X�?�Y~��>|�^O���׭k� ��<p�x�(�%��u���>�㞩��_�f��g����I�.8�D�E�6�4,��;u���(z�UY	]|94�i���>��Ή�LS���)��M�S�M�[�+,ǖ��в��І�"^®��ak[��x��K7�dn������xd&	8��/se\������5�	��蘒 ���Z7�8z]鉲�����`k�B���s�8X�`*Iz[W2������6e/��{2͏Z"�C��/�_]%0�]��R�ي�7FF��]u�R�u��72�X�P���g4x vҨ&��"T�E��Z��D��@��%���a�W^�L�~(����%�lc�T!{���0��s+��Ss����%.f%)�l'��5'�y/�P̍�ķ*��)������9��m_���
d��yG���}��#�$��:x|�j�6U�Z<zItǧ�I	GY<���ެ�����d$Z5@va�K4���E��Fd�T")�C�Up�xc{q�z��io5�����3.�o�n5�����}"Tv����� �O�ˣ�-
�#�`�gVޫ|S���N�V;�I�s!c<ᄼ���s��(I�?��������Ę��
�\�d��{m�]�6$�>�*�0,��K���<AWF�J�{Qr��ZT �x��!���JEF>����^K��Ƨ�pa"[�^-�v6=]yD]����U��"�W��`Y=�p
J����y�fDY�-ř�K�$�"��r��/P�4�7��
��(~`�L,� c���x�E-4)�Em	�C��s�4�o�m�r��z���y���qua1��`Ƨ�74/T�΢ ��{q�<�Y_1��~��iWM���Jb�O;���i$��I�5��Jn	O����Q����J����U��v*h?fw_g�{e��qf�C�͌��w7ta�Y� ?���H0�ź��v�]%��]ӻى����Ⱦ���e<�Du�[��I������f�nt��ZA�*˻�w�Z����o��e�
 uw�u�	OAM���!����}qЕ�|�P��*-_������8���A���*��&͏!�Н��~�'��h��ίg����3|�p4>��� G�`��5�'zˤ��=��rh<�$6a�ٚ%��
�(��ܼ�TF��w���3�x�&[r�xޔo~��uӄ$w����z\ n�L!�ͺ�^M����m��a��;e�}�����[+`�I�G�����A5v=�;��Y�#���Ƕ�5Мz��$k]ȡu�*Zmn�-<��U�'TW�w:���4�"lZ��-�}<Pd�!�R�B���H�0Z�l�'C���o�,�?1$)�>Tt? �{��b�=�� ��-JT�'�P���b���3]O��{�d�
pSBl���� &����
��tbi�.pzv$w+��#fy>�tw	�Q���k�䫫&��YR4�� XR����C�,�ZF��g�K˲W*�Q�s�o	Y�,��R&� �%R��oG$g?�'.G ��"խ����`Trζ�IO��R�,������x S <>I�	�W��Ĥ�8����FK�ݾ�����.��5�����f�فз�-V�˽m�DH�eުx���$P����#�]FKOE.���G�[
Rf@gjB5vZ��j����Xc��?)�{�e�'���`o!9Ph���"���K�h�濋@��=�Yg�V�r '��t!c{�� h(�#ZZ ޟC���Pц��\@h[�לn|�{w#D+Y��+G�d�U�*�B���U���aY�t�M&lfy\�G���~
6z1~�,՝פ�f�����^�Q�`FRK��6�N2U�Z���\�8h!:#�y���+F�b���Ϫ)��K�%R�l�4�<�R��U�$H���a>��j��<`&S����&"���=:W�T�GGB����Np
ƌ6�g���t�:<�W~�O�Y�́�C��'��ЂV�2'�����UPh�8��&���G$]���I���Ғxf6�
���&���߁��e�!�M�7���IK�j�̛(9>�����L�iݘV��+B^���+|N��:��8���g�� �2���`�9���k��۝\�NtJV4t�O�3��%�f�w)AO⯎}�!w&������.JIph������$�֬1}@.����~b��a�)Q0PLc �=��R��u���O&>�eZ�h�	V\�ŗ��1R��ɰ!��Ɠ��uD���I;�)H�@�R�~o���QE��$�&���w���v�ݖZc�E��+޳�:�.�Ɖ�6��!�T�b�c��$.K(9��c���=����_|Z�|&"���dJ�.�}[q����6�a�$������,M�z���xX=F����	�߿����KޘS0Ν@֑/ �?S����D�o��| �l�G-�y>��#���,�\P��1�h��&�d�o���r�+����Տ��+����e=�����-�7^��Tރ�=�C�74���9���O�+I#�:qHU��V�SĜ<ݓ"[݂%���Bd�R��R+e"S�8$�w���U�Ǜ��`k�7�a��I
�'O�:<�se���}�_�5�����@�mz�;�f5��P�_�󕒺�sCw;Y�vM^<�)�|bm��`��p���}��',F���zѫn.�E0L-�Hp܇�N�f��m �����>����?�/��������轌ڐ�%��Csh���>���=E�8����Ъ��_�["�W��Ć��8�K��ab��v΍�M���D_c������+���t�Q�{�)!7���0
�a�<�����{�e�]�Ak�u�3��HE�oH��S�a������Op'�b�9/�I>M��t�'PE�]�l��C-���yz$�Wǘ����:ͬSh��s /ia��w��C�z����P���io��ĺ���}+�� �F�A?|��J�EiUچkZ��)<u��N#�k�O�8��i����M\@ɯ�10�f٠�\d������"#�+��op��|�+)F��a�,�MOҳ�
�U�Kx�Fj8ނ��WB�2T:Z{`���U	�Au}�F,�����So�d�!{}ਨ�M��s�V�ց��(ȃs�6r��.�?2���Jg
�q���Õi�bU��:E=r1B�t�JQ��B�:S���+��Yӎ��pIۤ4���C��%��)���V�t��{(�;��/>���M��%��J�>#���Z��o8@�FwWT4X�G׃0}�߂Բ����[���K��n���u
u��X��r���
��<���<�M��F��q2p}_e#�;2�Z��ߨU��_HA��?�k��?�P| ��[�ve�Ed&Ue��sE��;ci���r�\���X!dI*u���Rٖ�o����O?�n�����d~Bh�����,������m�la�A�q���w���AzfFW���^���!ie�\Īk���'����;�7X���9M�W�_��~=�5}k4��ŏ���;�m��+��g��-x��O�A�j���	#Gh3;���6��K���ȯ���oOx�^>|�Y�S�� bjF��
�<iɤ��ˌ��I+]e ���W�gJ.����0}RQ8m��Iʵ�)�f:�$yiTѺu�0�}��#�tE����j���A@��0�� �����PU��|OTYA�0������#��������ԄfI(�s3���\f���T-�!�P��(ߓ�V������ɀ�~F��-��W:mr��BsH���o�Y��G&/���3�����AH\�������8A��_��7.����C�r&C�,Y�D��{rEbRq@��0�n-Rz�����͝O�H���ETg��~HD��Q�AI�m�/9ʤ���ewЍ=ʈ���y|��[���Y�Xܦ	5Og��S="�)i�$�U�N�.���8zÑn���@�!�������`��!���|{я���� �~��-�ȱ/�}��h��!��p8�t�GR3!l'����.]H�Vs��gXX�����ş��Z☴�H>>���-�C����ً!��?H>Y�aF�a�A��%S�������i�Y�x$x�/��M�����e�� wV
4�$bˑ/�C���Q���i�{6�Rq(�T<�J�o+��շ%&������Dځ1�%~�\��}��<����x?�P�i8�r����&�8�8���
�j��b����;��eZ���m#�~���!s�}���Fa�!�xȡD��U^y����:NgD�eL0'��/x�J)s#�����j�-���P�l��p��Jɹ���%��.%�d�r��ؙ����^�0Υ�!��4��Tu[���$�p?(�P5��9�����,{�jl����<�Z%��al�梹|x�OYP{��8NⓏ�I��CUX K! �=p��hИ���@2�� �˃<�r-�_�U���(�g�V�����S���ѭ������٪Eo��3��u� �g�()$��;��f���H0*&�������VS�<7�Tu�������u�.��ʖ0o����G���Md�*~��0�%� {@%�M���@�����AEɘ��B�|a�z󌉽j�ڲ gK�R:�,�W�[�u~��*�i�^n�;!}A���O�Cn��oX����Y눟:�u�c�0 ��腚����!Z��F�����Wb1eыBc�[]�������tH"v�����&�q�a�l��?�!�j�>ܜ.
�;Ԗ"6H
�fmF���:rfVaf�:(�7�	�c�.����`ׂ�`�Y��k"kb��t��"���� ��@��p���9Q�O�| -��9Jǡ���n���_�~;�.9c����f�l�e4�aX�,���լ>�6�h�h��lثc@�Y~���^U�zQ��&����Y�J�r���pK~zI��e�bw(���B�ޭSDNn���ʤ/	��j-�+勾����p�j���" �Z�ƐA�m#�v�ź�E��]"˝�&T]�;⑧����T�"�^�Y��2s�b'�����$X��^�fq��D�BI���ehO��mb^����\��A�dq'jឨ.����;�J�<���H����8N��	}���¿K*���D�5�"�[��.�&�/�֗���,/�eWW�'Es-:����C���&�Io��;?KX���%'	���5��a'��i��i��N��_�����-�:�=�yT�J[
�(���J��;�?�q�A�������T�3Vv�h����ݗ��]D=#��F�֠�p�N�tW�"s�q�|�@�A(�wƚJ�N�;%m���H�C�E�]W5�Src&6�0��b(�ϼ�k�:�� ����V^d�wU�a� � ��1��c���ڍ*�K:������ɶ����]y��t�~�� �/�v�<#�Ƣ��C^=��څF���� �s��#)!{�AG�y�����U������z�������u�!���� >
9��((������I�!�6ށq6D'��P,Oj�2��k#푢����[NH渞�@o
�,��_6���X�ۜ�E鯳��Ś�%T�&�"�u��3���	�?X��l����� `����8��!�<攧�]}���V\gM����nwD<!��!hQY|��E��p @�@+F{�z8�]����-�M(2���)d� �TnH����L.��Q�;���'5=�ٟ��2Q^�v>�����.ϓ
����=1)f�w/%�6��L�;b� �j��4�P��B�^���3�:�'�[��r2�d�;��]�#i��zr�
�$�Q�y�9\�#��u<��l{�����gֻz����.iw���5��*���:2�|�<NQ���ф��1�y�� ��a�&wLeMHVE4z��4�su��\���O���P�F��j�C���6ȶ�\Mg�)��J,��T�ջ���b$�	�z�z�Q�)p9�G�7̷ڿ�s<��'R�����o>����)?aL뾷�$8W�V�W'��E˻�X	��f��L1�\�s�S��f5;�uķaW`�*���O<�]��[�a��	�o�����,�~������)T�]/��?qq����=�F��!�c9�C�I�=TfZSͿÖ�8n��p8<�Z�����@�e&򣚂ɼ�D�/	�a���n�*/�@��]�'��*�R)!��cz;Z�hdNF��JfٟD�O]V��]�aG��P3ǹ��dʕ�24:�7��xuJr�Q����� �o{�3�]��M�i��gZę�6T�oH��h'����vR{�Ű�L���i�4��Q��5��5q�a��P�8�簏���$?�>[��Շ"���YQ*�Ѱ�c[U�����9cN��Z�vhf���>�9��u�o�<�#�4!���°���ۨ�\�PW�.���%;����t�!_��(�yb)��d�}=5�C��D5ЧS��,�0���zH�c/��uY
f� �w$�y�F#�ju��rr�o6d�ՓGƠ�Ů�ZW-�D�j��OhnbD�c��Z�T�$�GiT�:�m��o��, 2趟v�TL���N?���VY?9K)��o�������`T|��4}�,��uc3
�!�¸Z<�N��Q���ڪ	���S��s5x2m�sЪ����lr��N�łP�(fp��� �E��,�X羂�㦉!D��g��K�N�U�5�\I�C:���O%��1��ಾ'�
��Z�Ť9,*�A;7=�x�S`�f&y��OC
IT.���G~��!/o͛K �����C���7�(�I+F]v��s;�� qY���À�NaG^I9u9"-���h�[�0Y{�HQ0a�a�{"9�v��QkH�vMIB���j��Z|9���Y�;9 i���B�V���S*(!��2O�M��V��M����Hnf5iy��zQ���R=[��2�m/�eJ����+�2"}7��_�&��s5�k atɁ�6D����"�d�d_�R�G�Q�K��l�a���\<|��S��2����=��[;"��+f�E�G8Z�a���i��T���aJϋ��dCn6�/?a/��,?�GiS�>x�m���%�)Hd:�	�n�SZO�����%r�
~?��5�Wd����.�%j�8�.Xr�U�������員'*�Px�q��#&@&�`(״p����'ˇN	�W��C�*Bz���'E Ş<`�j�H��՞�R��|t��/	^��F��g�M]�E��rQ�.�i{�\;\Fǿ��v��X�)��M����Ұƺ�Ӭ:+���f])����`�����(#!ƆdQ
�p�D�從�	}�v��}��F�5��599	�&)�-�|�R��b�&��)Q1��M*�7R���ԙ��[0����x�#V���P���bF�AqΞ8m��v�5��k�ڳ~뾴�4��1Ϯ\P�Bs�X�Y����e�/"�{�*�a"��tRru�@��HZ�(!�OjC�	7|R���(�1��ҫr��jV�뀴h�5'52)EO��Je�ݵ"4=�jw��q�BW�����|��R�<w�5Y\@5��U�b
4Y>�s5�yU�k"�[~!��9ɩ�P�E�Bg�~�a]i)��2
��}U�N��'+jV	6������[)5�� ��8�D��r�<^���&����T�����f�H�e�2,e��Y���L�,��k���ٿ�b{��l��W% ���C&�l�orؖ�7 �j���
�L�'i��B�?cU<6���B�#�Bp �� �wsH��yA�(�ՓC�Η���iPlt%����$��wI8�	LL�eƐ�W4�2�AUE
�d�e�s����ty�o�H������>�ʕDә�m�x��%�Y`Vج�%�]P���HN2Tb���#('�1N��!�����b���%�L����#�~0�#��H�����{��u�i���x��bR�;:�a��R.8�E�X��/
���{o����G&��c��R���>Q�(�<[a�_յҌDh���<V%Em��Zp
�>��~rs�p�^*�=���T��lR�W�ո◳[���4�Ge�+ �t+f�H����灌O�����*��t��J����W��
�հ-�3W��P��u�{"␷~I���W�{�(;3^!`��޾���I����:qT����_������t��b��x[ն��?a���˧��,v>���z������4��T�~�@�h���ɨ:\���ޯ�>hj;�!c{zꨛ�������ݱ�)tS�%��o}��j�8�v��L.f�V��l��K���*#nc�����Rw�����&ܠ��~a��o���{�T�l�6�C��U��[Y�WDJ��Q��}��N���ZV2�;Uܺ��L)�4��߉ovezEes���`m9욥S���]SS�G��^ZX�iY������^B�\%��~�c�7u?�sJ-D�zoys/�N�/�6�i�Y{(�}j���,��D�g���f�ۻQʶ�H�m��*����3x������_v��H�҄���4��,�k)`z>�iw��wx?��.�p}
/���L�ӑ�N���_��� ��!�e�h�_RV>���
N�޳�Z}�� �:F
2��A�w|�����3Ʋi�F�
��n 3�Cr��G��1���XQrt4���!ۚ�����4.�gvm{��̽�G�j*��QDK�3M��{MM���4��S(�ܒ��R�o�q9N�#<�zqp?��5
u�DjR�:η7B�4b��q#��d}�a�JNWa�p��:�@��7�76��/%^@�}'�v��B6K�߾O
��+�S����M8&oε���j�e�5�� -���s�Nﯨ4�U뚔� ��B�j��^l!/|�:g����#��Aei�� ��-�M	�������� jZy��J,��8qQ��`�mo��Tc���Xſ��X��g��Ϧ�]h�t�o��p�4��N�Ti�EEɔN5S r�����p�sڙl�`�v鶒���|�6�χNH;���ŶHS�
��c�ײ�9\S�4�Wv���NJk��%���i0}��I3}@{bxR�+���Z��"vN�|#�='���Le0�%*�uV�[�`d���� �H�o���l�ֳ`Z�S!F�T�Q�®�����&~Ss�T�l�qm��*� ��A]�
��Tm`�J�/:uqҸ4�Dz�r��lu�/����T�+�yԮB���$Y%�1I'3zώ�GCnA7�/^�$&��^�˄�kHo.�O������iS���X��<�pѼ߰K�\��]B�"�Ã�eIg���W�Sq��;�ٓ�@M֟�G�i*Zj�y����u�ɇ��>pʐ�s~��e�n�&[�<$7�i�{+�"2ÉT0���� �<%l<WZ.��h����t�ϹǸ�Zte8�m��-|)\�K�X��v�}��`Aϐr�@"���~[V��Sz�����m�l�zጱ�7є����s�Ѓ��e�bҶ�6�F�����ŀ��6�;4�2\��a���#�pe�ک��|��'�Y*�k�螑�90�d�J����Y* �H�O��sӏ�N'����1��=�C���饁2~`i��>@���J���DӼ[|� ׮�+�EEפ��w5����U:Ģ���:AכR�L�c!_h��Θt�������< ����o\����)���i��n<h�:c�j�t�,vmE���i^9��7��%w��)r ��9X��̓��hq�'ޮ�0�w:�6�'�%��87��޲4d$qm���<A{zIj��l2�]�K��P��d/�Rhz7Y',��ACm�O��qݧ��ÿ$~���\Xh��R.w��).M���,�Ҏ�h�NDx����v@]���@��܌<���^�����,+�j��;�	DG�d�փ��f�G��Co9�7�$��W�:�2��C ~�?�U��T��)��uB��c�!ߝoy����͌K���:2W�7A��y�0.$G�M�(J�a�[Bו��~��N�9"�Q
� i���O�r�ڍ�k�+�/o-
�n |(�_���W]{��Nb�����F��P�6s ���[�$�����ܗCi���������L�e�o�[V'`X#ߕz��1�X�v��!��X��G�^�Ɍ(&�O8.��;���Z9V�O-��r�Ib�o_$��6%�݄h�[p�G�:�(d+0Q�<�a����é�z�z[��K"X�������#��l����!��3��x�˃,���߹����Vզz{�Y�n���w�Xo�}B8V��N�*Cn���j��d�/D�o�yZK��:��	0�~EͲ���j���SȦ��˖���~��EMl��b��{��0溣Uu����	%*^���������.�����a)��ć�B�ʵ�0$�s~���EA�Eng���T.�x��`Ի�,< �(�"�m[#{dאAl0���uͭU�/-ȫ��6�J,�1*�5�惬R��V�ݷ�H/|�nf\��^���p����UO~	n�d�B�5��+/���h3���ȢٱI4_)&�����%ӈ3�kew ��د)E����B��؛7����$#V+a�Ļ<)�`o<�� Ld��&[��[t=cP0�$`#�`����p	y���Jgm�jh���a),O�+P�w���<�}����|�����*�՘:�K�{,fŶ�(ߖ[�E�a��4��R�S��P���B�g�-�����
��½hb�[#��&g^aTyMl��	��n�?{e�X��̀��vm;�~N�٧�}��𪶜z�w�	������*��M�x�|�s��0�޶g�_�eh���[˙/�DDi�t4��lt�2J��e�X�߃J��B��Z$�S1�dX�M�9��mVz��c7H��;�{�梄Mg:���ֈ���3��b�F�y3�ޫ{�E5l7��׷C���IJ�B(��br�,Sv г ���a+�V�++��Iמay$��j����-�^�X��w�9(�f���6�LNz����t,G5���<��K� �D���!m9'^���t$�[�씇8�6ħN���M���v�&�:��N�ш��N�g�Gky�R��*��g��K�>p��N�j�d���g�*��L���G_�3C��e��=Y�A�'7^WKF`�/��ü��Pk�'��Ӫ����	�i�f	�g�w�6�ۨ�H�m�B�(��f�M��F�~hy��3�CQ�ʈc%���Ù�f~����?�/!���T��c����'腅k+68�^���6�^�?�G9�3bU�˔�kI�x;��S�����1�.�%�ۭ�> �+�P�L����t4oVH}r�,�E������3M�(��oJ��f���Ub�z�z��;�n�=+�z�m�S�'�k�$�t�e�,�M��/1��v`��%P0v�YO�ʤ����1=��	�W�q��ۢ��8~�-l���˾0�H�~�m2~�p��Oy䒓¡7u�(��¦�'M��|�5�)�n)��9�Bѩ$S�}����	�j��$9�C'?�4���� ꙡ�W��:\�|�����h#��Y	v�P���?�����CoN#���E������}}��1Rٶ7���k<�ߩ�@�����O^�"w4>)D�8ql���%�H�V�; W6brJ
T������Z��N�')�>�������=7+?�LBa�q�ng����M���Ϻ�`�x�fU,D��%˧u��װ��AZ�hdϸI�:�}H|��d{@�@|����V�7�~�vբ�aFp[+�C���a*��SnY�0�1��ךZջT�e��R��;eW���R5�射R8� O���i���_p9�*<׹h�s�vH��t�U4��S�^j��຤��n�4~%�����!���@��v���9��A��6��a�x^��Ū$��g|�,��S�ъ_Y�7�چE�����x��iP��0���xG�=��GN�`��6E��ޛ��fc�B8c8 �yi+�%n\�9iɥ��]��8���Nd �
�p��_+Q��]�z��m*����ڑ��rR+�����Fi9[
���!9����4y��AaNAš����ZM�����e��2z�i_n���%ȓ3$�3��g$����s���FIb�u20CYۅK�s\�M� ��S�r�6n��;������z�@��>1$�Cݴ�3�D��pb�-��D*=�ֺK��v�t�}1�B�*�4/����3�R) ���0�Q\,��D��Ҕ�l[ݦO����k�4��f�(('{��è�kŬ
�P�UJ�+W�C&�f��4�(ǔ�dʋ�DA6����xi���C�fɋ�v/o�R���RHy
����f�%3B�=����S ����F���e�+e HCV����� ������#8�a����	�F��\r������7(��S����H�,"Z�:��_B�m�������tv� �R�PS�$rXE^��EAX:�b1��q�p���1�ev�V��g��f�\}^�є&وO��ª���R�`�st�i���`���;5��+��m�,���u��糛�Z}zo�6}tlvi �(�=!����:�V�Ǥ�?�n;�zlR���9$��O�5$��}��e���ߐG�:���}g�G��Ir/;�F�1&�$������>�����?���D��2�b�/�`K%E�}��pt.3�K{BR����fXYƇ�A5��/k���H�1(�L��l�f6OtU�NW�12�^��엖~݂��n'�S �k��C&�3&G�!�"D���4��,`�o �@����򫒛B�4�_vN�����y�aי7�	��U���p�p�e;I��R��r@2����Rg��d��t%�4���v��^�\��V�<ږ��s�1M�$�J�.�b�2K-U�㦈�E�;@O�8S�g/�3�6�7�Z�LA�c��q�j����"� �v�ɺ4_��@|��G�ű��o[XH@�x�'A�m��.�%��9�
%���믧[��&��d%��u\j�ED���@Ŝ���<�z�4;�"���qn�9:r�)�Ϯ���1�)]�
��p�q��ݝ�퐯���;�3��pU�9�`�!�=G	���cX���S;a�s�U��['dv ״�-�kQn���{����>FZ����Iُ̛ꉽ�_L"��0O�^�e�ybz>-��i��Cz1�*]Y�Zx�16]���P(:�oa�������u�I�o0��"+�̮_���x1PW�	�K򞟦�U�&�@����Q�G�9�PcWr�?��~P��Y
|�FE
���\؇�f+b3m�ʡ��I������b����x�U��Z����3Z����C�5{Gw#*����5���V@S� ���I�+Y��N�K&O�l�	5�U���T<���<^^��|��M3�(m�V@9b����S����˱
�FPԩ/P�8u_����@��a��r���c��v-p����İG��&+.���=�|B�bz��*�������gƏdY*"������A?Q���%�"=]�xN+��~�䲃c�������������p�$U�h{)�+�D�#29%\���8XI���!��[@�!�Z.cO�0�U��sm�S���0k�&��1���}�����1Z�d����Zu��ME�lg+���"�����<��*L�+������+8x�¦):��B.R3��>=M>�c`�
gN��\��sc��R=�
�A�ur�̝��P���wC�iN�2����0�8��y��v�Y��1*����� %�
�a�����Í8�G,AO%wh�(,��p�G�(%q�Z�C�������%o|�=�5Q���I����IA��$r�b�#����.y��V���VK�^y�>��T�;�k'W/+)��%`�!q��	Ժ����,9YmYL�wm���^	A�8I؇���_Dv�I��w	#�Yi�t5CL8Dj~��m�P|7m��8Ji����{��1.�|uc�6�iU=�]�j�B+zn�Z�lJ9m]�k������ßtvM�#��,Z���{OJ�W�d����_-h����������4Y����c�E�at)�:7�w�"O��A�~7E\�G?U͙?1�$[��!`�r<� ���S�A��=Cd �iC
a�	��op[c�!���Ӿ��7�Kv�Q���Y`xe��y��-�4��'?�'x����}{��\v-���rN��|f�Q��.�ז�*k��>���2s��L���,���eW���1.��]��ĺ[�.n$��?j6��	���E��h9�N/�9 �)������k�B�N�"��oi��F;����+5M\��u�@I�DF�C�}Yx���C��м�)-f��g�)�O��D���zE5H/�'��d��E4�u�ͨc.V�]5|���R�u\����]X��$�#x`�QR��YFV����s�C�$�i�@x��BԪbz�I�.:���W������7/��,g���Q��lR�lQ��	2�9zʒ�D���{�0+������>�n�ͩO@��:�"�����ĸ�FC6���d��x�Y)��?�)2�O����ǊD�Pl�
��?��l��=�כ��}z�ѲUeZ���,}bYZ�&\���ط+��k���)�Fu<`˅�{� ���0+�('	�܈��. FL��x��<����;ޟ�>~�`��a���4�<]Ĝ��]��J!b�p��D�;e,��]��y�󿕷��f�n����%F�3����-�3ȏYB��µ���@��|�5r��h!�?T���F�z��A�v��/��P��D����V�q|������K#�@-De���[�M[�#���:�FM�����l�C?���1���5��.�T��ҿU��������������m�m����}�$�:�С�d�������bB�F9��H�̭9�J~"��RE�1�!u>,���PO�i�}�dȔ��`�zf褑ϝJwR�����\:]��K�T'ηS[ϼ�*�����+�YӨq}���8K|���s�XRt�#oI���L�]��<&��6���hG*�J����k��K^x���g�}��(0*ܔF�^~Ĳ��8��F|�z�#�7��-g^�!]���7S$U��M�	H��>@:��Df���{�[���7�A_-z��B�`&�~�3�0�m�&���f+���Q1���s���Gcd��q}��Xj6�P�%81N@Q�������S��G�Fm꣱A����޽̎�`�)���j����L�t��� ������ T�Z9�ɐ�l��z)P"dO;�8�6�ѩ����!� �-�v��,BW�Fh�
o�#MT�N8���k�Z�#� r3���X8]3�4ա ��;�\�� ���D������[ϋ���<p��N�Y���6�o���%ng���ѦpX���[�aܽ�SC	���|Ro��V�J�=W�핛��C����>U�{6+��)IO5*����\� ��h�1��x��?G��2�Q��������t�~�Q����x_n`�h��ޯ�ӞE��.vUs����_�,�[�dO���7�]h��ay�H�侮 �:���Ԡmt���Ȗ�r�O��Rr��璪t?��Ġ�>��9��`�0��쵬�5�%z���Hkl��!�f��ޏRF�
�Nל���n�1Xo�,K=c����ν;�ʀ�����}�R8���4�}x���-�)o��W��#o���cj}�^k�Z)-.��U��|���8,a{�ihoS�+P&EȈ_fdH���Lu������Q%qܨw����5�i�=��[DVRe{��i��U�~8 ,f��M�1��F��|❿���T	��V�η��
+����B���%����D�9��̔��� z�Ğ6�v�e]��<d!�c<ޮ3?h �F���~E[�z?�_�Ï���zSua�@}E��lqT�n���Zg���b(�:�j��5�8���������7���|)��y�w�]�ޞ�o.�/@���E�J��{CO�y
:��?��Y��h>�T�q�3�Y��,���;���8�o�d�g��S���6|!Ļ�Q�&�ѫ{U ��ju�L�덷�0�a��0�	�y5+-؝U�¸޸K�X(ZOh��]p�$I�t�,�QX�8�#�NYr�kXq�y��A��{���囻P�3hE���x+t��H�O�'ʵ�(M&�8M�Di�A®x���/�(��G3�i_��k�?�40�<~&�p�SaK��\���:z���a�G ����P~Z#�k���� Q��P*	P��cG�V�����������.;&$٠<k=�w��Rz�Z�|�~Α��H��OPsz���F��<%�OX9Э��	vs�R���9~"��l6�<�#��= hq��뭆�F6�f�V��	}�I��jm� l���xe9
��Y[ğ�o}j6`�����()ұ-!dO�����[ZC���p��z�Z%\j?^q��_ww)�paQ*ʾґ�跻v���%���tQd��h�R���mUl�e�
��+�ּAll�[<S�9*�:��d�_�u@����݈�'�g1V�7�������C+k�v��QȂE_0r���E�ƴ�	᱁
��U��
���������6Me������A�gJ0If=� ,�%�3��<����Un��W09�@Z���vm6T^1���,��0R��瑾�4���"���?
W�+t���U�#=pv���Ig�a�n��ʐIA�,��f7&�&�6mU)��w:^ph��	R�G�l���h;�RB�K@r� *���!>Q�����+Aal�b��l����Zn� ?�mB�ϰ�,6��AU��)-��`?��,h,�^�i��@���-/*�u����ڊk.�3�����m�L7���Nx�4+@���j#A�}���Խ�!6�v�Q�ћ�[cV�Т���] �V�Q	�ꄘ����Ȩ�JLLL���ƈv���7��k0�#���)�WQ"�Kf�����W���aN�wp	�-Z%��,Ea�ma���؟�!'��/%W;�X�d�zEm�GZ��=.%c&\�N���n��6CڤaW�� a)����!t,��=5[\���xξ��� ��+��`����2R��&v�������m�g�#�>�:H��~���|m��l`3s�F�AEy�:*�}��x������Ci-Χ���iU~��;j����@"b�u���N~G���|x�T�Ã���(�:0ɵf�gk�oe��k;���"��.��a��r��?�n=�C+�u7�����deP�!H�.��Y?�E�;l��50+1+
�~��SI�O��:I���^������bw�����th�|���mٍJ;����$o�ϳEH1�^�14��y&ش#�}Q���k�n�x|1U�����r���g��QcySX�%�z;���lQ��o׾Mau���n2��ey�Ĝ�Z����0iT]�MZy�b�b����!�m�� k����c>x�Z�vTפp�iQ���4G�u��M�z�<���8$��K�?�$pDQ��,|A�f��L\�M�y�@v�����ݓ�gW�]���'�*n�ߤW�L�*���-�e�
t<YA������h�γŧ���%�����#��upIH��>p���F�<�Ց9}�ɶ`M�i`/���&&q+4�6ܙ�0���~o��!��f���s�l���8L�@t �,�
��-�B�����P��-��I�	�����d�ǘ�I��a���!��"jt��l3vkJ�'Q��Tq��y㮉��he�e�X4�t��n[pL�l`zƏ�⛒\8�>�1o��<6�|RҖ&��$&�]֟���  �B9���bu��!�X--�k.�e\�2�n��vr��ʂ�m�V�lb��
�j��%M��8���OI��{Wc[�_�ewq�=��ĳ�p�%L~k�����s}�2�6���w�>�zA(�LZ��F��J�����x@�o����B�����	�U�Sb:�|<%��.P�X�ڋ6m/����4��W�3o.�xdե��c�+*0�7�p�����|�d�;�Lb+7�t�!d"��ϼ]yΑ���vh��pE��c��ozto�m����~U[�r9ݮ���M�o7����8�ۤtZ�#X�Vg�3qY{1e@x�d�nT�v6Pϧ�}�:&�v�'�_D�d�3��\.��D��S4��x�`�
��ld0!qŮC�����%�}��ׂ���U���IZ7+<�!�������J_()G�4^y�fk#�ɔpܧ<��s���qYyd�N	�r�,E�z��yx=
�o!���<���!�|V#._�Q�k%em�q'V�������-nU�׭*��ٕ��΅��n�4�mi;�W�6�Cξ�.�N�i��A��`��,t������Κ�r���]R��[-���x�m�=��}�c�9���vho����߮@�S���;X[;#]��:�Z�o��c�#���D6LgO�W�z�.��7������	���3C'3�
F�X��������>^E7��J�̕���������-j�8A���wF �k�N�8�<�#xlh,]TΥ��sXK��x��3"�`t:��_Ro�
yܗ���M]��P���$\!�\�П_�f=�9$��e�-����Y���:˘���&�.�9�aY�������瓁�Blԉ/w����ڬw�@����$d���p	]�4�8w��|	K����ًl� -��<NH��� �C'oۀ���3Q��^�:Hf�'��[ОF+���n��/�ntK�����-�Ǳ�rَ���*���̴v2������Q����=�;���i�1���4+s�g�yv����;�Ⱥ�d�О����`tx���p�k�@"�t��S4��)�~�%U�~����-��a%�c�Ai_#H50P�K�����*�����Rm�9�&���;�v���*������TJ�^�t�_�u+�"���=�^�hG���{i�r R�"Z��$�|Мzcn��z �Nr�y���{K����s���e9�gM�M|*�KW�� �z{q�>M��Zy��.���K�\������g�`�Q^ޑ=���+i� /gvQ�a�vl��e������E�}l��c�ZTJ�^&gi(8yg�nSB��k�r�z����{px�;��9ϭ�ֻ>|2K;u;��U�wD�y��J���Ã٧��7�7�U�G���k�Et��oZJx�5a Ӷ�B(����8FÒ�XSU��^b�嚁5:��������A�x���8�pհs���8��G�<I2�"�H �Uɳ\yF:�V�X)�LWH�ɲ�ZF0[�2�q٥t^/�w>>�'����S�Dc^�D�R�v�6~��vJ<-|�f3��\�&4���w������^SjR�u�B���yk@�� �.������vD�g��}���7z&���e�R�`��:�F=dݰ�F'�����u����[�*�	؄�}0[!;D͟��n��I��R�
�;����S��	Z�b�Ղ�hU�Z���1M�#%����v���7X�,��k�Ƕ�.J~㮐�rj?�j��-0w���t]�M��iSv��C��}$���G�>�Af�����k#|�P�>,p�N:�T���?a�=j�Xi���s�/9�^��A%�J� �p�k��~.Т�c���=����o�̚�	u'��=
�B(P���8y~��yD�oF�;�q���bj(���N|*��ײ�p�o��zy�u� r�L���Ks1��]��> �s��@�<��{LY���R��#�A%��L�&4�/�e�A�1�%#T��mؑ<��V[8��eA�A�e��O��^m%%�M���x�M��hl1�e ���,O9�n;?�t-��(9�Y���=mw�mk�;HZ�hGR����HZ��7���h)�ab��`6-�N/�j��׷K^�5��}��y��}E��%�(��6.h�.:}�媒�X3����<F�Wn9�1�tP�X�d�͑Q��9����04�}
Ȑ���*�5��e��'-nB*����S���D���p�j�r�fOvL���LO��+T.�#$Y�Ӏ��}?���c3e�|��s�Dџ�T��5��;ݨj�;���&�7F�{~�n~�5���s����%i[i�������Ö��;�`����X]<�XT���*0�.�:���3���ӱ��a���ڑU�n$��G��Z��)R�1��r(�b/��=$�K��w��W#x�����!�=�!��`���j�=��LZ洣�8�c������!i�BnW�c�z1�������������U�3��#���/�@p���e�N�푥����*w~���C{�2[#�D��N�����\a�+�q���Yu�'!�W ��=z�BO��9�B�r�|�ԓ������t(y�1��؆�2B�w����9��c�h�		T~�"���L��Z����I�Q]ϱ;N�1��/)e��D?=���Y��@���H����}�6�vZ��q;�9h9������Mf*�^!���ϩ� GI���C֝sk`:����[�@�"X
����_��<OOm,�����yn:�)&�x���&s V��:#
P@���n�dh�w��Ad0����_��x
n*��+�R2:����6\F/�t�QN����p1g�X�Jy�5	�F�͟��1ɒ-5�}�Lbf �Rt9�M,\H��Uү��E�h�(��y�kɇF�))��������`py���R�ķF�7j��'_Z@�)^���5O�=D�9���ʩ�`M���P$�t�?01��%㒋TXjf���bH���3��G>�d����>���_��Ud�6s��(��#c��ۺ���1/s1�OFaF����f�hҰ��`�1ľ�1h9XvN��OLc�Bn��=�>�,:ՎA�K�]"��cbˬ������.v��_�U��G@s'X3������ED�.��y͔ҭ�N�X��(�����C�m,ݍb���
B����bY�T*TXFe|��'�%Oj��,���Ⴁ-m�y��kUc�\Ɉ��0�c�.�a$> ���ւsƆ�oI�]�v;j�.W�����
S&\���8�޵�
Bi��,��D���̇��cDv�K�$�+���+��N�W4L��k�A�e�" bJ�;��E��/���8^*qxl`3H��ivZE�>�� �\����5�ph�.�뱃�*�qfL~�&'�=�8y��IP1�"���->�{v�'6@Rg �3�A���F����L�*t�������YyGz��M�#�TU4���}�ANEϦ���,���<{H�M���`�GXLo���H�L���r�V�E̍�����������̓��0�RՖ%K��0a�/�!Ɯ��z
�H�2�3�9�"M�2��/�!�~�J�Q�a�'R�6��,��ں�	�I��
�(�Ǵ3݊J<�
�n��\�Nf�3�F���F�ݏ��z��9��IZ���x���:}�e�'i3H��	qdb�܍�L��E���:-���"3��!�"����dV�xrX�s�G��7 *�k:�=��1oGGQV��(,cW������Sv�E�j�!oW'
2�f�6����Vr���9+�T� E�z�*��LK��������)V����+�I̗��y܄���:��I�ç��iȹȓ9d�.q�wv^V�e>7�w���p(bl��{�o��燸���y��ڝ�F�B��J�[A*���{f�&<�iքK�=>@�e_ﴨ�=;�?�d?���{�c��~lY�)���zYr��3���(k>d���a^Ȕӯ��<2�ܜ4W��V��ݏ�m��ga
��u���IH<Ey����=ς�ŧ�a�%��6��&��%r�F�p�n�[uCGtX�sl7�͵�/'�|]�#�$��c��/�ub��~a4cee�c�֫Vv���I)P�'��w?��i�b��X���>�C��>G43��{�����_�j�FC�CVz=
�p$�ҙ;-�+��H>������j���dl��t����a�,��#W��	�������/ve��#���o�;Ǥ�^���3X�x���
ܢ�!wBs�x�!ĥ�n>���>�}��0{w&"ʊ��,�9ӗؖ���N�F�X�p3��ꈱΤ����|+0V�m�ޔ/�2�Jf��#u��A�yk�^���[�f{��  ��p�P�=��15p����� ǀ�f��c���,�&c eD����B8�z�W�È�0�l�	�	�D�=i_9q�7C��L8l�5��˥��B@�'2�e8� Py�.r�\bvE ,���A�r˝������_[w�}����!3҄�y|`��7�#y�@�,!~�m�Lm~�p�R��1�����K��.i���X=#�54����Z�uQA��¶b��I�l��͍EW ���$9Rt9�P���3b�cƑ@���&�šcK�"��n��Os��`�<�� ��;ɨ��r*BQ���z��Z����o0���	$W��JS,Q��(�������/=�A��	�����]epejZ~�.SOi����r� L�1lGmaQ7t�:�^7>5�y�.��Ԟ�9�]A��.�;�Ǆ��:�����>�.�Z�7T�jjQ�4�<-֝m����+0�a��jǄ�1̯�E�?��h%;D�W����)?���U��8/�ƫ�~w��~xP�5�	����d�O���ȸD�i���B-@ R�H�D|<I�ksRn�ct��h�yN�,��r�},k�:_M+�4�A@�^ն/WR���%q��h0I\���P�������Yx]c�eާ��,f�,;F��MbS��'�&h:��x�v��ރ�)���/Fo~�
��J	.'��bЛ�yV�ˢ$㉶\�w�������s�}��7�ϑ����8�ۤ5�-i�"�ҽ�θ6�����1Z̑J9$�EZ^c��ó������X�*��0ᩌz�����A�'7�XN���E��>j��m�}Bs��:�������������58J᥉mx_<�E�P��4i�ZU��8V�^鹵L�!Mj�����&��Ώ�]� �8�8	�N?����+��-�Z3����vIWF����QsA)p��ۧ9�������<�8A9]�	Љ�v*���	��7�)�x9�F�t��wWem<X�.S�R;�BQ8+Rd�����"4��J���V�տ#�X�K�p������H�b$��*PCN|<�2
P�X�k~�}�+��Zc�*��׬�Ex���UC�%��k�/�/>���Z�i�fe�HV�I91f(���?�xV�N:q]s�� Zs<��âƫ�w6\ a����E^+3���h@���]l9E���2�#�ERmr�����u�;SD��6>?e�J�1&�$R�	�����j���ҧn���]CD�΅���	����4�F*f��~>.�K�%���x8I�z�D���X�~&���#]9{�4꺙��em�Z��{�%�y�p�����q���u�ɕn����[�A�;ܜ���q��N�Ϡ��%c���	#zee�^w!��CQ��,h�
�����qz"���!@�o6v����M�f�����I�1*E��0:ٮ�B�Է�,� ���t;�Y%W8��m}�_� �Ϭ\�Dc������V�S�JɔA�y�4��̛k�&!X�������7+*�����}CR Sc���m���dE;���goNRMDzK��P��kq������%�+��q�i_�v�1���|h��/�Qb�����Z5j,���k��Ԅ#�K�;�+X��P;�dj;��T�l;�����\�Q�:�C`��8�Q�^�Pi���2�N�i�5Uk������,����;��>�5hq�mc�U{���Ae֞"4�5P�q��(�{���D�{_e���ὰ��4���c���%�>:.@���KE�|��4����l٪�Ŕ�CLq�å��R���6��G:��T�P�N漁=Ij�"b
��V�g9	,���j,w�9�����QhH�s�'��,G�U0�Xh��Ϥ���SP�����Tm��3l?2��X~*��G`9��JJ���$'������:�����!��@Q���sB����N6z<��ދ䮎�'ݕ<�p����-�����������8"���p�Nt�+��Ha4�w=�Q��I-����уx�۸o���M�uC2����h��H9���M}ۃYE�(eJ�=HP�����!�X�2�xZ7�����ku!S���#��,L�V�K�:��������2�<�9�K��&���4GPkd�MU���Z_�� @��x���?�x+���9�'���OUs�h�[c�$�e ��()S_TrS{���ۏ0���#��WZL�m�K�^&l�o�"�%n���]΅��h���#�e�\�_�z;d彩FR������ā�%!�wS�ˑ��PJ�ϸ@�v�	bYu��V�n�Iځ��[P�D�2��"�|UWz]i�@���'O����F���G/�)��h��H.}R=���`3�PtP���#�JF�����
�n nK���?���T���	$�4�n
�@/�'��y���cBF޺�� �V�U����7e�t� ]��N��s�5}>J�H���'<q1�L[��GZ�} d�r�%`v�]%�NYHdt<��53+{[�SB��������E4�(���0SoOƋa��I���	��2{%�k@�p��	� �I��y�x���-�e=b��y��MS�D�%�N룘K03��Fz-�*�tw��� ��IE��Ê����h��g�7�S{{������:v'�q6I���]$<�o7Rgã���'�&x�}�8�g㭪�y���v���%̫�1���l��|�Q��*�Q��\��9i�\�I�H�R$�ўr̕�M�p#� ve灺�; |{�.��OY���Y��O�b7���u�K!������̦�D2�F#�G�q��W(��L�����
�scdꋟ	>�M��nl���N��>���4Ȟc���Hx��ڥ���ƞ�Pcy��c�Z���Ȳ��s:&ѿp�4�Bt�d1�Tagm>���T�wl����A�ɏ��B�_],HO�t�Bɫ���0�pخ/�A�3���?ֳ�S��I��X�/C!\辣g헖&�o�ш��E���pq�A|2��t�x�Z cao����Y��HO$��ӣ.y��2e+o[��"���ل���Ī��ʿX2��0Iu|N���D�6��R���k(7��=�Hݺ�p�,k�ֽ�)Y�Q�y&(�z\�[�)����.�P��zv6-K�?��{��4�x��*��S~�p�x�ۘ��N��c�5��������{�a�mn ���}�ޥ(���HB˷�سE&�G[;rΠ�"��,�C�7�5����W�E� `=�ƌIL Vc@�r��U16(Ĥ�@%��s.���z�zן��x�O]L&Ʌ������]�o�9�sr��_������9��9��|V���vp�M�[oZPU
$s=�[��|���_��c�b�^��-?N�ǔ|�	D�+�D��'�"�Gں<�g���w�FO�>4@P�����Z@���V���h��2�jL��!�ڱG�ߖG�����[�>�7�;������.�J��G��&��.m~'����Τ�n�ƅ"q�k�lL#��'.�QU�(�gl�P��bR���tq���9C��x��Հ�Z����Eī��W~`��!H�n��!�k؛8%�tx��샱]���{ީq��3Y�������2$Id6�pKd�<�Nj�M��«[���0�C�7�����e�x�r���ǟR�q�*#��WԾ��om���0�f���e�cT��do��t�śkf>�'��8���%�n�I~�V�e���H� xy�$��2Qa�f�U���	�X �;B!.>)݃��_V�J�-�jόN�0J'���\�❿���}��5"�f��������9ਜs����1IF�Вw6C��g�����rd�GLe{�C��rUz/��v\�h�3��+G,�`z��� :7�2-�0AxerX�a�B�KOD��iR~���6�ѽwH��Sn�nb��/ncb�]�4�k�	��)�08�n�T�소, ������p}�q�R��a�d�ܐWe��6�6�����,�m���|�/�t}��f-��S�j$��2���=1\I�'S��,��:�4��7���i��HN��o�V�$�]_q`\-0s��`��&�T�n~�Q,�^��3w��u|�1u:r���VL6�o*h!x;-!� )ذ��s�[��G����!+9�~��e�1=6�N�ЁX�}Z���Ɔ4�U��ܗ�H�ѯ~C�d@��G0<��J);�zH!�7�(���Ou$k*ˡ�)�°e�y��U�'[�w�|[ n�k��9��E�|�'"SQ�>�e���(������>\��W*��2�Ü9ֹ��Ψ�*| !��y,X�Q�V\V�xVjQ����p�����?�fb
���u�Jǉ��_�V%���'���)TR�����5I�8���ĵ��;G��Q�*y�s��a��\{6lk/���#��`N/�*_��d���rr�s Vq����+B#�9�� 
/MH�G�!�-<�K�P,���E�3�
��̛�v�D?m����6��f��;�Т�f�V��ut'W��Ԗ?��L�����7=���ӣWQ��+l~E��YL�hj�'M��uwͱz:���i�Rr�dP��99�咈���3�$K!s�5g_�/��/��S��Y�ؤ��\j
4�lC�z�����[��d�b���r9�o��ZM��Vъ�I03j��f�q��F���A�:���sk5y�ԴQ3��{�|����/F�>F;a���x�ھW�H����Xk�d����e) �֙D�o��	���ޮTC�%�uk���0:-\�wK� Q�'/rX�]$eD��q�v�a��+��f���wS���Y0'� ��t����J=Fd�
[W���vK�o��=����{t|�94�a�H���#f�A-
���{�(�F���5k��۸#�z`�feII���$�w�$���]��']�����z��mo�:���,9�(D���+�Ó���`���_f�����Qt�)�'���ܤ��p���HcV��WX��NF�ˢ�aXs�����`���|��� ���Y��M�L���OO��
Z���IUҽ�J�JO/*�4�Z�q�1��j�K%S�<��j��H�i[��*>���e�˸��j�'&��ݺ1�g�?oc.H�R��)Ë)&���㰂P/b��
����ϔ)��K�am�Gݚ�2e�D��X5m����7��>��_�v�]9��_HWZ������a��6KJ���� ?�ev��g�z@95w�1�!�
��5r��+�	]�H�'uL	�ĽoKV 󋶇�ೇ
��ްT%�$?�PI;�^�KC
�������&/������\�o����۳V�ōg$5D����cȃo3��2E�3�:��Փ�3CE�T�Lc
�81�Y���ذ����o1���\�a&O���%�Q1��c���Zrϭ2;RtGe!�Z��K�g����NrV���a����L�ԇ�i�(vc�@�6����Ll`Q2��i,�޾��TT�!�a��s�b��m�|%�>�����* �Z�k�٠�V=��O>�kS�^�b-ƨ�z��!���ʟ;Q����S��)���@X�NSd�\�m��=���X�V�Ijf
)OK�$\�7�J}"�,�{.,\�f��H�rT&zy��]��6�*�=����6��7��(L�v��buB}#���c�e�R�d/��ó�̓S�5�����H�-�.�;5�*��o[v?��l#^�j1o���A���L����2�KG4���(̕SG�ZHc��j�r藣5E����p[O ��B�3�l�}6PO�:m��<�Y����9WM���G9(K���@�$꿊�Z�֥�j�,'�8y\�����!�Y(�ˮf�#b?��+J&(�+ˮJ�R1O_�����ϘlI� 0P^���y1����껄Q��̀�ƿ-�H*�':{v꺐uUhRپű]��I`�Wc��q�����FX2C�����O3�۰�-��s��h�"2����	X^*Ȋ����U\+Y%|��Ě�՘��E������rwˉ FY8�z��Q�*�M7]N�Ab����.֣�*��Yz��.+:��:Å�L��Uw���XN��I72pm�q�Ù/&�d��A��5o�8�Q�2�<��ր��2�G�m������A���_��I�o P<�B�,%!�]1�5MBi�N?���.�:�Es�}ζ��H���A�G���9�>���Va-dcT��P���2�l��'�^d#4Z������̬��x������9��gJ4�D�$�g)	�s�B���eſd�12�Я�dt}�ƪ[��V�RB
�Hcc6�<�Vw�#�g>l���rb�������Y��OКSV*�ZOf��t��I�ah=��b�=�zPi'�����|@��A����
D��xƯ`���Y>�(� ���r�)��c#,��৾>�E��Y�+�*4;5�����K1g�!�=���T��+&�.��;|}�#���ժ1MR8 ��Y0�(������]ڄF6��NqF�6�dᮠ��(5-^��L+m�k�6��%�T7���:�{���޾��ard��m��t����]��%њ�ښU�/�tU;ȏ&*ý�����Eo�c ��D��gs����HQ�)�T��O������	<"B���>�);�',���.r����0��)�QF���(a}pkC|��R��C,s˺l�K���%0.</�x�kqhN��|mo��E��RϷJ��g�N��޺m�v������Z��$��3ݰ3����otř�Pc�6�L��*��'���G�0� ��	!�7���H'=F��C*�n�j5�5)���f6>
��$�2h-GE�H�j�+�����ũ�SCK�l�	5[VӴW�aɤ�oJץ��b�֌��.͹2�r�� ��<ds��%}UT���={_M샑�R_�i7�ˑ�ݎ;cg��4�k�NW#�?�Z�M��
���gwXM�ִoO�<��E�2�"A�1̦%��H�&I����#�;�&��kHc��qRQy�6p�~��l�?���t
e��;��<1����-p���Q'`�]	caO�!w?H��dmR�rE�/Y�<�;����I	�������oR'��W
��dʗ���Ӕ��U?�P��iKX���g4�%�Y5m4}6z�}��(�E�-[|F�b+��vt�Թ9����[#�U�j{?��'�s��F����/�669~�J6�O1ԟs8yd�R4�����f/*߁Y��_�.]�M�nO[h1��v���#8·�a�Vw۝�����+��͚�dK�B*dC��p���0q	��'r"f��ɬ���=���W�l]>xR��u�#)��ә*җv��=WSb��P�k��XE�XU�	%Q��_㴽V�H���<S����oC�����	�q��<1��\��s��C�EopX�t��zq���_N�5l�4Lc*�ԑ0� ���'��kyl��.��`I��a���C5�j�������G_��P����8V�&,_�<��J^��8xЖ�VlF ��.ů*k�j��:V�X�pt�<�z�˄��'��~l25��|/�Ӛ�����r��q�k��c$W�� Y�+' �D�_P�k&7)f��̭�a0�ј�g�	K �z3�:�}�Q�F��7�?�$̼�����1���o�F>���U�brq��=8h�B��va1`�0��Hs��wr�'����*�3&�%�(��S��m���H�p�b��CR�3�%�Kg�&M��6�(yڮ��,��HRU���9a1<܆^5Y� ���-v	TB��Du>ݡ������/�7ݽ����~��ʯ/�ϳ�xT[�gY��2��o�KݜLד'Zw|��+`��7oD(@��|cG��3�ac��6�o^���Y�I�w��Q�ng��R=5T�#n����E G%2��N|���u�������g�ok�5)<Y�$�f�h�8����v�G�'@;g���
��@��y�Ԟ�H�?)�8?�VÜȝ(،M���B�v���V	2�A�F>�X���V�u�nK�i��N�B�C'�۽���6�
۔'gp5:W�M&~�H�� \��R-�&�̟"s�21�T�v�d�T/N���4�t���Mk٘ ��L�r+�����ZfCD&��l���ۤ�kG�-ϧ�y��6��[�����C��2b�y����'���Ʌ�����L��$Ë�Mw\�@����\��~��|%v�<BW����z0{$�B'���*m@~�mxw��un]��}	���#*~J'J6w}%O4x})oҋ"���^�,�b�������O\�����3�%e���JA���������4{}�3����kd����GSI�Q����u섃�������ju�i꬐C�?�KE�GB�ɕ���ѯ6�s��""Z|u�X�w�q������@�l�?äj��7E/K{)pĵ*��6��G�΁�n���jE���hSy8����p���RR#6M�Gw��f�����^�"8����q�l�F�$fŦn��gz�U��q֨�����O�����W�9��=��wH;w����̅�weWL�?&3#$M�L�x:~)�g��*�'9T"F�>g�\9(��a
�c@9ޡ���B�&w�������_�U\�2β8�E-<5*(c䱅{Qb��gNA�]߭Dv����
���'���+x9Ń�����]��qa��h�%��-K�M+U�v��V�a���u�zLK#�
�DJ4�ED�q^�K�YR��W��,ɔ��ꪪ�Ncwך������:T#��S|fݩq�.12��x���c$����4`9�͉��F��mw��f
Zm.%�/�Z�z�o c��4̙��ot��֯7�Pq���_eSxa]�C�t�QhJ0�.?&�D�t�����-�VO��g�m��'A%tYYX��_�Ǘ\�A��oI�/΀
�d	����賧I����s�?�o��/��l��$��ۭi��>���w�Uh
���ʀ˅��S��K��mOP�U���O�n93��gn�cv����s��I.Hj �@j8�OD���<Ol�tGx�3%��m��*j�a��SZ���0V�+�Tz�����@��d纜y�K��&�a�De�~zi;�ؑ'�������<؉Rc���x�+rd��!
PDk�������9����l���q~㴷gJ��5�F^H���)ѯ�[��aߕ�����8<ʾ;1���0��@�ɧ��M�$���&�ܘJ��w+�����H�z�MB�����- � ��Z*"����V(If���q	�}n0�x­�\��w� K��ٵ�����O��bW�a4��k�͙�I�;�����u�`#ɺ@���`�m
�X��*i�3o�T:IM:ʿ�I���<�"�,RB'K���(w||y�;��p�M�Ʊi�4�iH�	]`o�c�l#7��=�<�
o��g��VK�d+L��)�YYh��k%��P���%8���FIQU`�#�{S���W��8���e1��l���[&�q��+����U-�(A����s���Z��S`�A��^ѽY��\���=��)���0�t������F��$.�XS�y���Lj���ǃ�D��A�#��#����>;$�rM&��������[u�X�K!���F������.ỳ���f��9�a?��N,8�đ~vYٻƖ��Þ;|2J���N+!����Z�����IMD�A��yJ�gڊ+%>чF�s�`�a�k/�I�����R�T��3f������ߊ��)� ��E����21g���$��1e�A�����+�,�w�&g��cV�m�"Bd�3\��Um�Y�3��v�'��g�0)3G�L0��FXDU���0��ZR������яАЛ떉�Q��Rxx�̅��k�Y�X�ٙ�=\���"�0�����[@#x;S�
=L�5gf��(p��]$��"��Fh�A�G���
�{�Ҽ�p� CP��p?SG冂���h�[��L�dd���3���S �y��E��	�?D�+��s�l}M��0M�v��k��z+���t�j}U�Nf�;l�z����=�74< ��q��z2�����e`2�D��CLQ�C�hO���k�L� �}%N�����_h�5A�`.�����y�~V�9�K�u���#��+r��٠ڮ܈�|M��(+�E�[��ן�y�k���Bz5?��k�{��Vqt�'=��e�8[YQ��y��_a�|=TL�/[D���F>�GJ�fͨ�1/��r@o	�ppZ�q���{=3,�[��o�A z>��Σ\���WCw(�2�ՙ�C��\�<�e!�����izI��c�;�$(����GF��^�|L�l��rC�����}A��5	�y�5����7#�_�=���et��R�%7ڭ�x�￑<����r���8:/�^��%�o��Y�f��E�U�%�oNW�䨏�vʚP��>��Cԁ���b�'���G��2�Gr��w��8�X�����y0}r������y���15YG�����.<���g�D	WF�@^\
���uX�,�����x����9<�SH^�l P���	>��.�E��@�0K��ЮO¼���,W Jr�[�+טf6u0�����%S������쇌��H̼��v>�v\�����
��b�x�%��-O�n���+%�~L�W��?����'^�`��|w?��}���b�r��k�H�A�����88Q>�tF�7����(��К��]�\�+�i����Ͼ�w_���[95#=���<�FC��VA7���x:�%�ޞ]@�I2e�[(�!2��r�,�I�-	�x�%��.��M�H����g���B���A,�A( �Lmvb�7���P��0<�H�]Q���~ɥJu"�a��A�߀3�n�p~�J7��0��=�?���O���)��|��aj��kL�-G����D,X�uy��UL�7��I1�Μ<V�v\�Q�����F@�Ӈ�0�Fٷ��5զ
�tI��Ą��e�Q��#�7����t������ӻ�W�#��	��	������~AimJ�;� �F~jC�%�Ƅz��LG�v}�#�D�gV~�q��4ٿ����~'�a��Пe���+��"�l-v�r�����P���i[�Lد��/��z�HɒP�M1M�u4�R��48<^G�^��{�F4ޖŻ=�j}�yN��nP��N�߫(UY�����'R����VWCIy���,��FNgHy8�QXģ�]�� �� QF�˫�bLN�8�$Ǥsl�ZhU��^��.g���� ">a�Hޥ�g'���K"dۉ��O�����*C��b����A��l���FJ�w���� >"�IL���J}}F�#O�ܺdD�>�~��do�o�&Un�4ٰ:v����'"�}g�3b_�յ�sC����� ]yP��n@"��ڳL|m �~���X�O���<�M�r�ׄ�g�m��M�^���KmVߝ���k�5g+걱�LA�(�/�5öBc���q2��T��J���Ͼ��~VO&?�BO`^tC� �\v�7���Ū>�hՄ���i�rq�.W�������w�|��N���\��5Z)�'���A[j���p������~����Q~h3ϟ_���� MK�~�T�7?t��<nz����G �V�jn�c�y�U
{e�v�b_y���3OV���!<̯���zq��Yؕ��	��ۖ�d��ڬ��u�"� ���B\�K��GIDON�;|�|PA,9 M��)�}lE �bR�ZN���[��}HQ�2?�d���矆,d~ڞ� bg��[�i�ؓ$�QnML�`%��O���hΎ��>�ζp�C���2����^qD}�ԙ�;ε]t|\�\��͛��О�$B�ϑc�F�c�r���D�.�{ۺ6s�=��SpF����m����? ��g��I|�U~�`��,�`%���͊�Z���ꕗc�]tnJ�dL��ӄ�-��F��Ar��޹�#C{6iu?�2ɲ_���{�R���?ǹ5ِ��!�G����M��9��Kw�¿�ꅜ�}�#��|�O��p���K���jsS��73ct��̥��	�p�T۞��1J�"7)Q���7*/ZC>.U��z���������<;��(�� A
��Â@Y�E��\�r���VY�!�M�dHb���)g˝�����$g�4y�E�@-Nx��t��3V�_Ѭ�@� �I���	@��vu�m=JTU9���q�fB�}�2�S� �G���zNI�@�EH~	��,Kty�4����C7Q�q��~�y�8Z�U܏>��K��+$����X9lxqt����M�*���T�e�`�Τ���@�@#���/X=A�}ê%�X� J"W��k�!���K,��o��-�qH&G��-'��u��Pp(��%&#@H|u���V^�N#C�,�W"����5����P���kB���@��^��7<O'�v
�U��M�D��b`t��rP�Uzry��1eY�d�B�3;��9w�b�N�M�]�"����+Sve�'���W��}ݛQj�DVk��t����Sf�cBp����{~`�xO?A�2P%qA�W$E:%�9H-Ov���\6��XH����������9�)8w��fQ�n/O�9�?d�M^�+�|��4R� rP���xF#�^�̝8�$
�'�w~��ݧЛ*����,��������"4����AL4���X�惔����9�lӎ~�d@�$�g��da��Mq������?��a?��㳥��N�m��%��������n{5%8W*�tʓP�`�{��t���Ҙ!�֨k�kHu;U�u\;6p���IV�lŃ��"���_�]���X�,k�P�R�R]����n�sh�h�v��
Kp]�/�����<*�	��k�cO��.������Y
P���u�+�Ձ��Ԫ�=.�}��^��,6ǚ�@W�_AZ�be���V�Ȳb�SCW���������z��Z׽R��H.F�#!�d: (�:lg_p�s@�Nih��sm�I!xoh�L�P=��MwG��_d{�y�t�[W��������ң�>�����l�,w_��d_>6��l1�CͺyX�a>�~���ZÈ���љ�S�r)di�b��lo�jq�-����LaR�]2U���h�����6�ޝ�ۼ��ז��W��a������HP�*���S�H���+�덀��F��ݭ`��GA`�G�n7 !L�{�F���+C*���s�j�@���E��>&S@�vJ����=�'%�,��Qa0{(k�,����$W̐8e��<t+�����6��mk��jn��6�����Oe����I�^�DB�q���;���j�;.�t{��wtC� |�a���"�$?�:��N�έ��ȮqG"�-�e
l�νf��&P9+���RnSO���iJm���v�35�{)�!в�m���q�]�>��]x.�.{\����wu�D�a���s�8�����`���(v��\�@NC�9����+Q�`��r��.�b�>כAiU�2kKK�4B����3�\M9v���S��1�yץ�BZ |�#��U��+'yuk�-V��ۦ�\}��VO��S�b��;��VW6�Eм�.�nP�����KL�6E�`z'���s�|9�������m����"#-�d�rE���p
�E!m�jJ�BqoWQr��p�X�s�L�Iݦ7ZO%��󛶍�R":�sP�_�v��l������"����r��З�5����r��֌�XC�������`�[�� �6��jR48w�~�T�W��Dī��P05^/R�S�1�i�G�
��Z�(�|�J�V�|��?-�:��R-�����?��7��\(�Rb.K��=�wb�K�ɢ��1���[��} p����`{-:hٺ�j
2�D���-�Zuq��nj?��A˖4�\�Hs�M�������e_oP���3-�~n-�m܎j��޸r��|8�O�t0�j_N1��пOü���6��&����c�e�f:����������Gy��X�[�I+�r��32Re������$��9�Ǩ���/��j�������q�+=�����W3DD�rG�>y���=����h���ŝ@H�8��@��E�:���+�+��H�a��ߩ/B�V̩`���.ơX��p�$g�{�H��%�zo칺 #�IMV�t�ߡ�4��;�f��fi�K���B��R�H �%�c�t��6d��khf�kJ�2`\T�!��Խس�#@��wgr�%�D0�Zh@./Ƌƭ�!�PR'HuJ���.<�]��D��i9�y;ҷ:����d�]M/��*�J�4� �씦G�O^YuBԶ�qI�3����V�J��%8�8i�V���ږ�e�l��ű�����3�����L�:#�����T�Y��bB�+��_t�:[oe��*f �<0=T�u`��
p��˸7�Y�(/P���?��%
��T�I��Z��o�#�x��^���q8�������$���m���E�k����䧗8��x�n�b��S�R0�
G��M��ơ��ס{�<?R�KU~+N�%Z
�yU�m�*{�LV.h���+ٻ� 8X
�dη���an,�����D�z���Ǻ[f�%�j!�Ӥ�4o���re�T�c���$C������5z�NΏ��IZ�Ә������d%�\Һ��&��ҩ2�	7㣩�*$h�HY�H�aPN�b�A�m	� 9����5��F"����\-f0�+��^����|+�ˠ0�9UW�~������1t��(�"�8S�fT�� �=J�\1�?�/�E���6��Bƨ��ZW��9��;��|V�q�K(���(1���H�>r��V�\�	��&�զ9�kMM12aݐ&�F�X�`Vt"��$��&�]s� �Eקէ2 +���7�d.�/�f��j3m��3v�u�����(����"��Q2��a�,�G�X!)��������3D��%��7ř	~��`,r�=K��P&���,�\���������q��.��|�-^p�3x�L9�V�δѣ7$H��� J��ᙺ9H�i���7�)�^���~V�-d��wq�����@=$���@�Fx<���sR����ݙ;2h^dP���CZ�Ju�0-?�C�@i�Pϖυg4����	���?�dԓT8��%~*;	�2Cբwk�R�.�����*jd����2�<c�o�o�M5�+4�[j�Y����~�c%��d�H�bR���:%�w���G���?�]|�7��3�$����K�����y�6WƇn�a4�w��~��Kl���x1�~!w�1&��m�$&ٞ�9hq	{a���䫚�ǋj�G̈L;ƪ.�(��JU����	�;|�K���u[�_���A7�>3@N���Ј8��6l��@�5\��}}-v����8B	�}�g9�$D��*F�e�i.z9�ѻ�����1���B=�9�Mat4X୼x�����@IV�ݘ�<�8k����"������	f�(5
��<��S�iGć*ԶΤu(�[�(�w��d�bB����~V2!��83Z��Qj�tҡUrG�h.h�ϥɄM���Wb۬�ƚ@`�T4�[1�Кٗ���,��@�Jb���z-�@h)C�4/��Z-�f�S�r����|>��W;��XZW�����~�s��D8[q�(��Z��6=#����P���2�WUiO�f������}&
U�<<i���2�~��QLĦ
�\K��_�m��5c�sV��������-�Їc7ɂ�-�U��zPf�x�	�����|Q �k ���急��pF|rP�9��/0��k�:���[�L��%CN������d�`�0�J���$*G�&<^C�EhY.IG�M�[�m��t��D��^�'}���Y�����$��Zj�o)�ẖRs77T?:o�1격�C[�����1NfJ�<�gŋ�S���uXNC����zd����I0m�&yR����J��Y31QҥC@r��wp��y%Ǹ ��^V�2Xؐr��$>�y�����������f��� u�N��]�bYM��59�N�c����y	 ���6�w$�ٯ����஭�W���L�����R�j���3� �h����?h@(���)q84�w�Z��G��Ѱ4�\���0D�]���V�I�?c���T��<�m���[��c�`�\�^]?����T�ݵ�X�~�	u �Lo��U�q�4�v��eu�f��?��ߚ�*]z@Rz�pw��to�F�G;�3JPz2bJ}wه�J�lIB.���(��ٺ���קju�h��Wܫ(-���~.C.xl�{���c��
���xD���	Ζ�G���'4�+ea��j{M,� k����C�5oGI���������BV��K5.J��&$��c ���%_)�������XL, �6������9���D �ҲM��ϔ���:4����O��r�b(������˫F���#٤�Q�W��xS��O%�Ch�ް��c���O�Z����]6k���"�m���Zu|hAIG
C
�58�5�/��i]ZW��*͘MF��5�����wT�T���r��X&I���Op�9-�g�d]S/>j��}f;�����z���CC��o0�kYg-���^lù�X`Wd:Z����/��ͬ�(#p7�cཔ�f5�1�!'�����M�p��;B��|Vł�Cd��m�͞��l_�I�G����]Q�Z�ɽ����_z$�8:�2�ltQh�,Ϲ��1�M��8�H-.��S��9���9��:�����^ NH�Կ��2�+�bh��k~�a���͒�1Ke��G��Χ����e�u摭E룀$]ra�S�e:b��#��ƉU�y,�2]S���	�h�ª?��pr�Qw�)�"�}��du�=�������-��q%�mc}Y�	��`z�"f��,D6j2w�m���x��O�+@e�W��h��Ǳ���Q�1G�x�/�Y�.{�ԿH�T�=O�I�l;��8��y��`N	�n�"���q��*.џ:�޹U^�gk��	�Jl����R+,�M�P���f=�g����Y&2���w6�Z�g��E���~���$�n�q��-+�*_,+�#�E@S����|ڟq����s8 ���bUZ�L�(m��
O�#�٥�k�:ae��)3�:'�߈r�2���:�g�%ҫ�*erO���<���L�e���d�ڢ�.N����Z��ǒ�_�q߻�'����4�/~U�a�N�9w���ȥ�D��2�.�?
�k��9�FP���5N�b�0��y0��m�}G1��ۄ\2��(ﲊ�����ҫ{z	��z����bfe�Y�~#B�o�.a�n���;���\�S��5���Ex�E���*��p�1�8�q-�ka���Z��^�/h��z���W�>�� ���o�ז��斌�E�7d��P�O�I���O~L�Gd�&u�آ�d�a�)�k>[�챟P�.@
���E��wR	���)�Սk�[2 �'����6C� ��^��\n�O#��)W�WŇU���}����[���e�(%'�B#:@���C��x�Xc���O���*]�칆H�AgO���L�+]�0R�#/���x�]^�U�`�GC|�ʚ���,J¢���o�$����|u�H$�]�A�7�U���R�k��:�9��}�}hY���57��ZHd�5�{w�4���˵������Y�G���K��^�X
5���6�n�����B��)�ⶸg�= ʨ��b�J�@�+�A�Ǡ��2j3�w�No`:t�~��=�����xA��4���i��ĀO	\7=f:���t2��d5��e���!��]/i�s�%��2&�E��"��w���p|Wk7��+�V�c���(#q�g��>{�i����ʹr�0G�������0.�����}�Bˡ2B��љ���S��"�ִ�&���Ȑ��b�3P�,a��"?�,C�-T2�K�!��0[J��J]z�ъN�翫E1�._>�e;�jDK?����[]|�ɬ(^RL>Ϸ���Vyϴ-�:ܙ��<k7s~�FF��=��wz��y������#�Y��K9j*L���:�}@u����yox��j��..����s_��$��CHA��w ���{���'g*]d�.�F����0U�������`N_��/�{&��eQ�����鮨��[���a��:�s��ow?�CDo��Ⱥ�V�2L�*�J?Y����^gqw��qk�AݵU�;���yR���!���h�y���Z�� �Rph¼�em_��B�j�0A���s�jZ�l1����`8�]���YOivi�������3k�֏�~�����?㏖^�/�e��Uh�l���d2�Xe����~��H�Z���/���-�b��,;'�����*Qڧ4��>\�R��[��媎�]�QY�B�w�� Q\�⺯��Z�kFa֌´Y.fF}�;����
��߸vA	���T.��fI��z��5�6%�&�J�z֍xk(n�5#~o6`��*�N���tޚv��@YR`>~=��g��õ�y�z��P� �Fb��L�}��Θ��EW�P�	����e��(/k�R��1�����s� ����Lԋ�+�(%0%HS�P��h&hb�og*��F��Z=n�(�{�x<[lw�tյ�}�	qpԄ�Q�?
"����M����AM ����7����� �8��Q�*�h74y��dT��E̮ehb�V6_�����lG��I<�-�蹊d���\�Vg���+�&� ��x�ۥU�Js���_y6�(A9�!��A�"\a��Tr�ҡ�#����݁���<Z���}�{��g]7u8�󞔕,Ge%9�$�hak��X�Y�f�(EX��'���N����V��#��H��f�����Ĵ
u�&�HBOXno�DK�`#���B�Y�0At�Nj\E(w8���pԀ22Wn�Z�mi����6����nF�a���e��M8!<bPw睗m� �J0�T�!�g��Bd��]E*���)��۔f:��	�J٨� Lw8c*i�=��Q���^�0o�3�
ц�U��<^'���Ŋ25٪=|i�N��������S�GR�"�е���OZ[(��v�9�t����(�xڿ��}姩�:ڝ��m~/�b:�G��LOf"Z���������%���	#���s�K���5��ʧ�&�<���L�o����h��l����6W������a�=N���Ļ����ķ��M�9�ۀ��g$�̊H����,�V����ں =�w���pBSS����jt�M�ŖkO裇½hQ6�
�k͵�\q�3.�h��iު4;cz��ٓWu�i�jN&��
7���z�(�tv�;L��מ�CT���l��|�R��̻��;������f\��#�#0��	�����w�PK�Fa�c���Ǩ�J�w3�uk�J����oQ\��>�Ѵ��C�s����8�ЌU�� (z�?)��i��XZM�*aSB��ș�Z�? m��xI����2��n��ܧ��I���b�u��~>���q�EKu>�(Ԯ>(H�$ÆW�w҉�x^Uaok�������#�h��-������9��ª����Qo�n3���˰��fm��Z�Y��m����oh�*g�Y��G(���Ê�����,r�U�H���@>|�%�4m��Ά �L�-v��4�]�����t�qGQ��i�`L����L�T�B*���,Z�x���	ȜunE�,-qp�a�Xu�!-���\+�Ti�R�cy�1�h���&��.��f��sI��(���$*R�hM�k$S���&mh�"P���촯
݅�<}L�>�mb�dtH��t0���s�<~OB��p�U�_K�Q��8̉��M�C4�嘎k���*�y�Q�'�'�B*7@`�Q$������B#/W�:(�w8����3(-���Q������ ��{�����H*Y���ʣ��p���ꫜ\�l��R�#S2�L5td�+�DA� }����X� ��4�����Y9L��'0��p�e�>�y�k��jRt��UQIOCJH;�*�ʻ	;$u-C�`4�)�V���hm"[0pk	hY��ٷ�����^�W�Cn���S��3� ��NB�ϣ��=l.2�/��9� �EtǬt.�_�H9�O�6")C���͘���D��7���/�ʯ�Y�(��� �:+2q�� F`����JS���y�N�䓃tw�2.{l�7�ei��%ڈQ����k��pS���x�j׹Ėn/k3t�p��.e�顥�A(#���#�@o��� ~�F�J�_+,�~��A�D�
�NB�̪�[��^� ���'�T D��~���n���������������6����k��'M�Q�?�b��E^g?(Y*�Z��3��}⇤g�U'EOv5i2MW�q�z�j`��֦������^I����6�
�n��E��򐙒*pBwlW�����%+�04��_\��y�`�@�_du�rFޑsf����
C��K��-Ը!�"Zyf�X�� �=蛞;����W5r��3���s]vb���z��_��c�fOЯ"��KB�\�U���H���;��j��J���"���A�?�����L��f%#���z@\{��ۏ�(F$on�X�W��Ds&�V�o����}�#�� ��J�X��+\���Ǘ�݆�!����;���4�u�(d���j������$�R�6�s���V�WO9Tٷ�w+�/5�hL�x.St/�h���,�r������w0�������N7\�#�J�m"w�T@�C8 �}m�d�#&��]� �r�a����e*� �5�+��݀��-1k~��|!F2^\��z��y!��<�"��3���
v8�l����!//��<��_x����m�t〩��r��~6r�ﶍ��c�'ɷ&hz��-L:��Y�'
�+�,��oy����D:Y��H�n�i?}����q.�-d	2��GJ�[��c�w��[B(���8�։���$�;Zt�2#+�I���YF�_�,rox��s)��D�!�cȍ�p��=�,L\S��M�:�'�G�y�w8���u��5<�����8��f�.��Œf)�a^�!s����_�x��LnHm�Yq �-�w�}ٶ<�	l���0=�R��%� �ӷR��mZpU��u�����	�5<����.*	�3A��!ϭ��,����SN�t�]|64�I�yq�j*0��@!����]�����x'U>���mb�LjfFW ��2��#�b��Ɯ�E���Mʁ--ַD�C-\=��A3�����\��i�~�Y���]G�rQ�.�B#)�
����M��U��n����E��{�7S��xOnPu4fٸ�1u�x]�U�	��W@��'����TY_�����Z��JȞ<���w:�(��<�؛`��P3D\l+�}E똅�Wc(J��C1��Q�6r�����S��?���֛���s���T�R5��4�����aP��5W��� *��|��@=�o�S �>�z��P0Pk��g�����(�"�����d�K���i1+!u!d9��so�@�V�����<���n�At͏V+U3<&�dɁ���!#��c"Oa� ��b�����W�l��x�`�����E�l�u�y�TKD*�L�~��+tt��FFm�C�w��+	�I�������C^����g�|9�����ݕ�1t%Ő��%���4%�`	�d����F۟:3���I��1.�;d�d<,�N��[�*�ăb��
B��X�^�z])��d5�,-!S�U�I\�RQ�]U�PQ����:@��h�Wx8���Bby�N�B�o��
��f����Ÿ��o�����E�Ep �CՌP�:~I���5���!�͓i�#\ ��U�%�G�Ss�)a��5��e/J�9/����&�1I��'�����gb��ʠ�-�1�ZB��zq�+��?�\���ɝ��q8�(\�`�<�7-���|��H�G`D�h�Qw_b��5���K�!�������G�4�L#� ���Q��RHX��3W���r���U�82��_��	x{�)|Ec}��M��˚�!�7y{�Tܨ���|6�E����Z���0�yLk��O�_C�Gx3��0�[z�M��8ޡ�;ڳ
�1�v`���rtYFI�W4q�����mXLjX��=`��I߁.Lw�Z0�)��=^s��^.H�5�-a �].��L^mg5\M��c�T�2a0x�ڄ�~�e: bf+
fa���'z�
�ب�4-{'����OQ���<���h�en��Ym��c�#I孖�N�1����Q?-)2�@���f��� � ��\S�[��ɶQ��f��;9K�Q��L���e�aHH��k1������#۲2�U��#��$����@������C� ���n�"ydg�����@e͉�|��9��� ̎�m�>���S�B����º?���-NS�4�VR�v�҉V99���?\��~V՜�4�,��<�O�9���$J��������Ikܨ�X��f���}�4ota<���a��)���@ë�B|�������(nK
._qY�U�{O-U!`MV��-\��BL:^L�%l�����3)�^��G��֛�h�Y��}B�9��|�խ��b�q�ca�Q�Y��9G�n{�8�cE!��hv�o��Y&[[�V�ھ�=Ѱ�MO�����Z��#-��O���Lzd��٪%�Ҥj,A�Ln�\��F�0�-~y���~���!s������/���$a�m�E� -���8��̉5����z<�[d� O�\׊�A���FL���Կ4� Dg���a�9m_����p��h��9�v�c��� <����/�t�Aj�)�z)US�H
���%�'�������=�w��T{�Oށb�b�Cśg��[���`ݷ�_�pq�w�1�w�ռ0,�rY�K�3/�3
|r+�ܫ)Q�Q���N��s�p	l��WQ6����-Q�5�Y���G���!�q��	�D`�`����	ݙ����\�/K@9��O�@ϓ�(%�4I�!�A�L�e�	�C�Mƌ��F�V���l��t�r�v��8N=��V����s�z¤%���9�S�xnC�K��p��gB�&���g���
z8[~kv�kG��ؿ���{ౌc=��>ʇ��k����j�r��c\�t����lv�.���S
'�3��k�'���
�>bBxI�m��n!���E�C%��`I=��Y�W�d�z&wd�J-�k���gC��׬����t��q;��wÂ)(ݫ�#�<
?x)����8�Κ��k�*0�=�qz'�lXܴ���gWwQ@@?���:�Y;ީ/=�K+@��x��9v�n��|�J@9�s������.4��hs��Y���H���(���%���.Ų%�����C��k<9h���e� Dv!����"�T!�x�Zl	�'�y�??U&4�ąu�6	3t^���PV>�hW]!�u��F%��=}T��)�.�ܧ<�ԍMԃ����_<�7�/�a^ �l9��F�S�#���<�١����]��՗����Y��ޥ0Gh� �z�	Dr}��l�r�Vo���*�~����nM{�3H�<���@s�`{�mn��ruOw�M^r}uG�U�GEC�DG�}��E��|���rX���ѿ�����ky�j4,U�hԑ"r��}�����!l���=��!�p�^�ib�!;1`�g�0���C%�1q�Z�ץ�Jgi|��1���BH�G(�_�2p�1Ʋh�> )��>� W��b(�Ǳ|�~ЇY��F��a9��]gD��vQl7�=�Ô}v'P��z�[޹Ge@6�R�����5cM꺴��O���\3	����5���38D�Ǫ -�Z�v��&t��N�jl#�@ժl�C����s����wOh��(��Q:��m�ԃ�o���'D��.W���Q��������@�����g����d��B��vNH���1�aK��N��0�
�L��i�˺{i�V�AG���bM��ȏ���7�'�1Gu`̢�d'��c�6��lƯTΦt�5�Y�IW?0�̝g�|������y2�0>)Ĺ%�M"�����r{Sϒ`W`C^����e�C�E.0~�ִmŨ�I(�Z�J�u�|�OG�/�|�:�E����d��Z�����u��ݑ��J�!�:|����&J�4F��0�ٛmk���li�y� ��ݬh��e��o�>��)�(n�q�R1���[�+h�� �����"ԡ�&wiZV� \҆�Q�^�\���x��f�l�N��C=�4f����G<]t�P-�R��j�U��"�v��Q�,@ �pa�
�2��@P;���8����,��GK̠a��� /	ZT��Q��������,�f���Z�߃(՟x*l�k��������������:������ܳ�ZUbR�W��h����{���B����Q�Rqg����[�-J�O?¸7��nQՑuH���j��RW�.���d��CO9��a�� ($�NQW��pQ��Q'��M������'}�y�Ⱦ��$*Z�𙾆G#�b�d.)�k"/�R>r�;3����3�Z�2")���y���X�F����PP��W4XZ�����J�<��M�R�E2`�����6`��ؕ.��p|Rи�%)�G���<�OHr���"����c����
�� �	�?`�3��O�T�L�7]����Y���O�_$���7I��)��%۴قÐ�+�O�ˮ��Ԯs�t����S(����/	I������ddq��cH=�%@I����ɤ�,����na�Xr}Efs^�M�ͺ�|�KN]�1��%�^1~��߽��-� �]#�~c�*������\=�R��B��p��'��P��'q*.�A���<�g����&��@�k�6n�JvM�YЪ�zda�s��o��7:m������7F�b���g^cd���ǜɛJK��B�ѱ_+Ǻd�ĚzAϼW������Qo3�R( 	XB+��co����R�F� ��a�d�j����]���\jq {+����yGr����>�10Ac���_'^f5{0m�b�s��.�+���׼ҋ�--�J�x`ګ݇�u�y5Iw>��'X���@y��Q�H[�7�Ur�ٽR�r��.��
h��4�c%��|2�̋�/�B��+����z��{R���P���MucB�o�M���m3���}�q��Pߎ�	"*y	U.�g�fc��}�ڙ^�\���l%ؔ������%�j� �/M��$�x���[6��Z����a�oD,�QL���-
R��l!A��������B��&p��?�'��ϐAAMKɛ�%Z�Q9�>g���Cڟ�DZ��=�-@��_y��x�J�)��/��S=���*�U��П�2잭+��O栉��'[�h��c�'<�V5~;)�����ݨzӟ ���IQ�Cv� 
g��f`N弇#.�S��@.��*�͸]i|Q{���� �Г�-0��c3��\H>�Z�����gf���D�x썕�3.P��줐d�Ȑ)��#\���ei�T�LK�`��J	'��l|	�dԣ�5�=�Tn��������f�Vǔ��zF�.d�3�ZcL��l�n�+�ZӔ�b �Lm$�K�g�Li�������aq/ǈ��ۧ��2�?�A��E!P�����ENQ�z^��Iӥ���p$�b߽�2�3p_��1c�~��"U��>з�h>A�yMwҤ|EzS�K[��E��p
g��;1QZ[�!�8E���Vʪ@�?��BٜRI�q��N9)4�t�T�V��Nw�"�䕨��
�3G.y.S@���(�H.K����X�fp-d��:�k���(�L�>�W����gl�l�Y�\�RVף�`S��� ��z~�u�_�DPe�W����k����x��L����V��=c��4y��#��bd���x0�(P�_�2��%��������f	9)9611���.���9�M���v�Px���o�Ü�E���Tg�/�J�a���?f1�]��d0z��=�{E��si�r�T.����]R8��XT�P�:���
�6��<�ߗ�1�[�v-_��y��A�k인�O_"��i��ɱ)J���y$/��:�B�*Q�w�H]�tu. ���iӼ~��yvJmeQI�S����ڎ?�T�0�����p���>���W��2paT���l��6_�Z!���w��P�OL{Jց!,wtD�1��r����� M�H�:��PU�R~hWR��]�s�j3!J��"��4�Q�>ҋ�\�]���o^�Z�3f9�A9O�O����Y`c��;hubᤵ-�@��C�Z����w*��/4W]#���kav��nS���ⴰ��4��f��	pv[���1�̗�����]}Dé��\XB���vu��pQ]ix��%�t��1]\O�ps9J[C-4Iӽg	~�P�!�q��~%���~�z3'»4�8P��1�R�;��?W
O��'�S@6C2�E�Z���Ei˓���0��@_~�ҵ����d�t�m@��kv�����3�(N����Y��⾫R�ʈ�1-��i{�CM�Y�hcٽ������o��w��k"��0�ʽ��*ʉ�u�!|C�f��9�)��,r)�)`5/MU�?����X�}�Ѷ�L�*t�u�=�"�Kq�<_h�1�\#���~_���hpJ�J�I��ؒ����=3E��@��3�|6\O��n�%iKO	>l�NA�8)]�o�ܾ�D8� t��Jb��܋��=�3����cꉾ񍔬�Vʁ�y9�)�nG;�5شS#^F+7���!���J���{<�I�#`��"4%-�I�q���[�پk�h[�UZ�~p&�gRSֆ|>��������/�~Ǵ�L�`�5X"1����=
�H���J*�c��k�*��nrV2�7{��5c� s��A�����)ɚYX���Ta��`�L��h�����Yg�Ֆ@΍x@����Z��FW|�F��@�}����lü����?�!�AG���~�����w���ܘ�:��p��Euqi��6�:�[cp�s/����rON��x��-F`�|���4��4��!�̕HX�.:1��7
u��d5����]�(�;]�]����Fx�ĎAj{��>���+%8Ԯ_6�Ae`\���w���V�&Z	���D����
�Tf8��uKX�h5����o;_JL3����M�3�-r�G"stQ!y���N�G��f���	�MRZ[���ə��V5��a�#3T\P�<��V<hq��s��7@k�O��3a0F�k(�f��顦��[�����oSJ�rwUc�m5���mr)�$��wRŞ�������<�&N/�90H�K�a��j�*i�PY�n��%ݐ��b��o����H?��=�֤.v2�BO:��Σ�ڧA	�t��-��n�����h�Õ� 2�s�}��*"�� � a����'?ӓE*v����NX�
Y ��Ip��@DLY����U6��e��a*\�{�zV��,��<��ݭ���g��(B��X<���v,�F�V�U���m��@\��Q)!��(H�PCz2��@qQ�N��	���Z�g��Nz�5�ޣz�+	j��jL���O��k��
�%�����Gɑ�t��h��@�z&���u�/�h�!�����N�)��FC�B��E��-���o�X�I>;u�LFc�=��F�]������D׊&�|"�r�q]w�.�)��wG�C��������-��;��(`�R'L�5�G��,<A#�>�'n;tX�ާqF���ަX9�<<����Y��^X���K=˯s7$���>�|�xo��J�YH��_$�����L�j���RUr�%���z^��L�d�1��%<��	���`�
��W��T���\�Z�+��	w�E��z��:|}�"j��d֞�M�)�{��]��p�b�ĸ��A���?}�������B�z=)�$N��.�%�{q���o��=[ �h���!Pi��O�}���6���8_�u�e"f����{�sDlV��k*N���E��]�X
��˞�#���O#�I�4a|�\���^ Lq���hm��q�b�Rls8D6mh��F����$z��X%qm2�!�P���ñ_H^��a��"y����/ȣX�󭨱���B͊�Q�F1�!��]��¶���|�^�񾵼S��|�����ԩ*�,K|�_�&A�ݐ�5�݊?��zH�*��3Α;R�����/p��6�=����x�p����RBe��͝�D���:?�,���tX̖��2AEܴ�+s�@���*��P◒�����g��?4n�Q��y��8��{i�tO�Sq��x�hA��<�z��]qL���G�K�8�8J0�yר����ul=���C���-Q<�`�Q=y���������?��W.��qý�s�N�Ѽ���TQ�vĉ��Ӱ	c��
�4ε{#�$d�2�5Rƍ�zA�����Ը*�@�/�������5ֵ���"4�56"Sl�'��|��Tv�_�i����z*�w|m+ e/�����\�O�-���ǯ~@�Љ�Ԉʇ�xx;5P-]^��8qO��P�CO����0}�gM�F|v���'��E�p��b��H��>`�4�Ѥ�\5�#��2�%~��k�S\��*���?z��K��4t��^v�^�z����% ��j-t�l����p��&��wg����ޥj��s�����\!*7��#��
M����KB�H�>CR��C�;���� �Jc��5b$�p�<�v�S��]�_l��EāD#��I,�W"!�w�%We�7?"<H,��p��Q'�+���F��I+4@�u�ə��g�<}J���$��y���<�
y�F�Ͽ���_<�YL��W��9��>��{��on�2H�z�W�7�h�7L֛"V*Y�-X�S�l�����}MXN�S����2�Lm���H�2j����ᭃ����~o7v �K8Gp���"gd� �����6��3�8%�*U:uSߒ<+��`|��$|ͽU�88t���QR%o��p�ɐ����d?�0�,�2���)XY�|�dGڻ��HVh��7��S퉵y�~�[�z���Z�B)V�h$B�?�&ӥK|j��3��i��z�l�$��=K=hncX�V�s*�
�ǕX�T���-I�i���⹘�������	�M�)���妵�A���̋�3���`�+)���ќ���of�X�&�&��,����@�b�t9�� �=މ3U"O�;�,�w�'ګ���zi'9X����u�i%�B=S�Q׍۟�#/~�b樋������1�sz��V�hғ���%`�}ť�dC��}��q��הּG�	s#�O���y��#랹	�;w�.�L���KU�uü�s��^}�e�h�v+/��b��4�9�V�c��ύ�jL�$<�E]�8�m.~�(�P���n�e��;	Ch��&��`8�&�;��C����������fKU�3&�c{�U�&�;����P�\^B�h<��z�ɥ1�߰/�S����Y%�<|��p���ޒ��x*�P	��#���mp|�,�/���6������w�귊��q3X:���_���#�c&�;��I�7<�9��ǃ��2��Ӣ��;����6��d"���Zf�&�|R���ʘIc������Cg�+��90����[��[l���Y!�����#c[CȂ��z�k@k�o� ����m��5�a҈`�=qK��'��A＆��Y,Vɐ*sL�)�!y�y���A%I����TB�ͱ"0�㜸��gk	��RO���Y@0C*���6d�iS�h��-H�¸Q���������5Z]��1���KG|~H&�hqʢ�� ��WĆ�{my�$��'X�a8w�����Uw�2�,2p����	F�]m��=D6�.�#l��F��§�%%͠)tu�� �D`x���P�u�k��}�"�+�3���7H�aJ{�-��b3�w @W~0 �F�L�¦X�$U���c��!�QL��!b=k�����A�'>?�	>JӚ.��|g��Դy��/Qγ��X3�ۮ�^�5��є�44�H���ٲ�"����wW�AE�4~Zo9z��5}� sQ������ ,���M
c7��+����=���E KY��W-��k1nB{�-u/�4�+]�7�N���oؓ�%��03�7�l�A"v�> ]J���/���]i�r�k�D��~�1]�������/ ��[�z�I��D�b	�0f?���M%���,R��8�5�{ڑ+����Qm[���B�/���9�Íoa�e�� )q�A37����	��`�`�ɺ�Q�0��C`�-շz��"~�13i�!oS	Ǘg�ytOJ���-RvX�\�b<�#u�R� ��H�c�>�ܣ^����[2>�+�ܺS�I�֕��~����?J~ك������~:�*3��5��{[�I��2i,U��ϪJ����v*�S�c��me�8X�mmX��<�N9�q5���u[<w9+yP�Dӑ�1e ~"z�s���`~��G��өtC�-�܀i�56/����?��ڑ�	��iWH���N�G3��d�RKc�Be�ò�ZU;�Ё��/}3��\��2ƽ��;�N�X1�`�T�`E��=������>��}���}ͱʥR�y�;�kn�B`r�R�t��D4�,��n��6�e�$CV�=zh�W��j��.ϴ�|S��~P)���g�FO�n�-�-G>@�T�;K�kDB9���U)-m��/�3�H���1��f��a�C�3a��"��Z�Lw�6��	���B��f�P��J��v�^�Q'Hf6�/��ֲv/S��R���a�P4s�3��N�hE������s�þ���\P��G�g�?w��Rm[k�υz���&�#�,��4���b��ׅ�Kr'm��X?k�d�X]4��ǩ��{�g�����z��M����X���/k�����>�q	������gw��~�o�L�{/�_Z��;ygΘ��˯���Uv�����B��ZP�7)3I4qg+�.,�?���K����A�eV�����ۚ����5r!5<ۛP���3�ȭ2��ŢJ{|�E�.�81�;�z�r9��E�J��/��=�����'�&jL߂AVe����4��L�F�1G���<[�wM��MrY^Zr6B*���6�̣��h�uT0�>�Ox4�01����s']"ؚ�S��f$&w�v`>>a
hߓ.N����R}5V���IS�E.U�AZ���m��$x7�g���>7�X_s*z�����͓TRằD\cUܞ�S�o��?#$���il�m�4����X ���([��~8�b)ޠ�'�w@o�D�}��nb�ـu����͎��1z��枯(S��h}>�[���H���� �ɧ�Gk=4�y��]d��Z��Ѡ♗xj9G�,�]��z"��/���\ų*"����tV<���"���"�����Nk$-���H,>/��a��dq���n��aR��Z�хL'���Vl�R?[�U�	��y6\�W��N���eɺG��,&�^G*��*�W�Q�������M9U��8&�T��k���qzW��Cv��F�Za�bFw(3o��� �[k�ҷ�.�۩�&3��1�B���l'hx��F޳����>�T42�TO
G��*M�妛�3�n
EYťCI ))��%���_��AgТ�kR�բ��N���b�����{y
$D˰�N���O�2�5�i#`���T���"��Z	�k���<�'��XiB赘c��)~n���H�x���ח��W�D��R}ۋ��%��b>�JypUnz��v���<�� h�+dj�S^�{4�c���2�(��<���şf��B�4��+�p���y�w��A���^u�EbȂmY�~�y��e�	�!/F�H��nN���+�HM�Η�c���;��MN������{�p�?o��)�p���;�s��zg���龝2�o6�K�K��]���������N]U��5!��ߖ�#]���)�O&�aKG	��ɬ���/=?�h:���*���!�s7~��Vf `[M6+љ|x�(V�h��"Y�����@�H�N�/��*�ˮC3|!	OM��d������%Gqe!����0�����秩�p[�D�@��c	�N���$�w�Gr\1�=�kX�=EJ��>d��fe�8��N%��8���Z�����ŵ>Y1���b �3\z�&��]9�_TI��������r�٣-V�9Hċ_�X���M���U1o����[�huC�46� c���u��\2�ir{{��\�PEC�cp���>�����8g����1K�ٲGo;������Υ�r@�]_]���C9��i��"�kݯ�&���K,�­��gL�E(;o r��e����tZ>)�ɟ��W6�PnCr�]�|�tT���n�z��!J�T�Ϝ_���ǗS��!#�`�R�0^h����U�
>��p!�(�S���%�K��{N�p�t�qK��jI/n��C�m���rt������H��t�9�C���o�c`+��iL��z��.�(�M<tV^�PC��v�T����^(*L��A�)�kZA���f��;/[�1�=�a�}"�?��}�4�*�r�&�OQ{�t�dniCN"x�O���ra�(�1�+����� �1n޴'�+��.\bR�-hx�nprE?̫���@���Y$��_�,Q�{[Y�3�gQ��iX)�h�J�'�n)��%dd�Nil�F��d_"V�sğRv�
�}9Ԓ��p.^��;Y�֐+���L� �㇀��!Z����H�[��W��K����q���"U�s�T�Y��,mjw���0�� C6�zq��6!����,�{Mhv�rvMG!�6���)7Կ7��>׋L�s���ԲSP�e�� ̃К9E�(ۭ)�~�R�R�idܜ�Ļ���HɃ������O�}�秦�IN;�NMo���"?l�a���#8�ȤrQQ�Ր(�0k^xBJ��Q(�`M�vp8{"���[�,���{�; ,h[�i�&\���bS Lm~@���zX��0Y R��&[-� ����jU��v�5�q53����[d����{�}���.Jӓ���(PTY��G���wI�������)�����;���p$�]U�}�7�Pg���W]X>_V��ԫt��5{'��^�ŀl�)��g��-�N��d�]��w��P,�ۋ�+�'��-'6 ��$?�O3l�B@v���2������t��)���tɋߘ{���"w,{J����3>�AF��V)�JO��c�NP��w��F������Y�Nk���P�.
���o�4��liP�r��?����*���D8}����Q��I�B��������)�F�Ӽ[���lj}�e�E���p�f�;,��<�5�P�&{U�x��P�l���lكa�@ze~����XЊK��K���/�P_&��j{!��6�M�uW}k�w�&�£PY6d.0�������ȣ*�e��eݎ*��Oce,Ȃ�}&�W6'F\��3�9�L�z���wR��Hا��'����HR�KG�W��d��ۡW�e��y-���������B����o����� ��8��uk�� �U-P2,�ֺ~�z�Z��8����!��>.�J^h�n��3�tm���V��'�������Qf�@w�cN��ǂ!a����K{��ơ�(* �pOj{��.�\��٦����D��4M���� ���R�4^d����Dz������T�^}�BU��E���"��,�+:��r��R�0i����ph>"�Y��	�-&j�?W����6���2���T �R!6Bdȡ<@Jd�7(B���W�U3�#�"XE��c�T1Z�GL�UK�]jCs�X;5�b���f���A��y�`�`��#��dQb��=�h93�j:��=:zP����
�<�2SJ��_N_$Â�4��ӏ�Ol�e�M��N�ab�ĭ�,�?@��� ���7��[�XȪΌ�0i#z�~^�Ρ���DlP'jf:t�{�iqZ)gy�-}�b�D�t����vgn��sp��� ������᏶Ss%J7����g	;��&�R���w"pՍt �� ���DuS�G�s�)�*ä#�cHcЬE��Ovq��L���i��|�@�/}�H"�Zl��Mj��&-���o�]Ӯ�1{�}׍G�A89�w7��О���50B�K��`?9�U�L�'��a�c �F~ǬC7���:,��Sy_��މpAc5}-,f�؎�y�\^�3��2�%:&��	����%��)�ۺx4�I����MT�g�]N̞F�R=��9��IG��SMuۗᖍ��I�G�ӭ�*0��O]��%�@N:�L�l�?5���Ѣ��/�J?����h'�ה�������0��{Z#8f��|�m��B�q� 5 M�� �����:M��I�dk:=�X���`��)6���ܭ��%��t��ڍ<�#IUs���|��H�Iv$`и��皭�%VG1��+���7n�XX:�o���x�v���W�t��x�	���B$�,��UIb�X;|r���E���A��do�.�O�F-���]|��l��I��H�xu�-����ߣڬ	����e��{"1��~���IԆ��E*���\��F�L>�C�ۮ��Dq/�����3�uA(����,��|ؗM��@M����A�<���s�|�g/��op��x TX^��W#�+2Z�bҘm���ڌF��[���T��+��
��UU�����!1y���M[�I�=RF(s�[+va��qc�A�i��0��#�s�Y�}�bXI��V�d�_��O�Q�6=�����F�Sbx�m��J}UWqO�`V��J��}�b�?�'���7�%��qc����=��**~p���/���M�M�y�)�_��+���E���i�/
6���i�4�l8L�P!҄��[8u�X%s�5(����\a�<=n��?gc�����Kz��s5�kŹ,���O"�Is�f�Q�C<�*y7�kh��S���g,(ְ_��Z�%���`�f�з��4f'���Q%Γ�F�����4Ǝ��@����_�6��ı����6C�4S�����B�G��9<B^�$@;�TŖ\$t�;�p�a�nt �#����u<���P�\5bY�����R����n���b<�4�@�X�N�"��Ⱥ6�Zc�9��]��S�@Hu���/�ۢ��"�cf�|־� )��ћs��X;M)�cKNhw�w�J����Fc�9��nr��ҷءY�HZ�I���	�U�D�H+s�[_�
Hl��٪���:�*�JA��gh�&�T���m�> �����6ϋd8{$����0��ͷ�����-���c8N���x���֛Wr&����|yϣ�b#�����
*��;uH}uT�K��vPO&�(�;�@�#D��V#1M��l��5dW���f]��D>���M�g��ir�Q�p��	��M�����b��MT�d��.Qh�ހپm���դA�v�y�֟�Hm�b�C�h|Ra�a�0/���7�یv��'���`cQ�I��:E���Pf�����]۵_>݉S��d��ޡ>[���{�1�ӌMn�Rm\4�Y�PLT;�[�t���6,�����9M���0�л@L#M�8~aɭ�>�|���,�i�� �f����X�4�'�@wb��Ey=�F|U�1�j+�'�����g�y؍�}�S7"�"E�z�t��XlB*:h݌�u�eg+��	�Yኵ���̠��eJ8jv����ǰp�n�U�+�a�>]�{��lLM��A���Z�W]/VY�Y�J����2�`,��R��>J	��\#>Â���|5�����u��DE�G�,AeW�����2�Ui��N�w�6�4GO@_�p
�}i
A��u�Ne^�"V1�r�9?�-r��2��૦�pHa�M>�T۽�i��]ȡ���7Վi��iP�Ũ��(���g�]�Ep�;��s�`�f�C I9��-'���pr�&����H�сR[A}A�{@&E_��3��992��l�]�n�wP`��1�	"���f^:Dر�-НꦛaQQ�6Q�O�iN��1.g�-g=4�t�C�2�B�)����s�b;��{�0�*?ݠ��a�|>`����`#�ưI%�Hw�AFt]�SiD�;R^��53��[��70��ۥ�QI:>�j)��GCԑ D��6oN�iH6P+d�>�)	ڙ�x��;
̓��̡��}�.'p���R�^q'�yj�0h
_���x����B�%�a$�b�Ad�iN
�a���ɑ��ǰ���B0\nE��uH�B2fl��YK L����sqͭ��4�b��[���+[@XЧ~;}-�54��g��> S
W����	;�a1E�"���Ѣc��r���6������"�Lm��dxR���1aLⶒ@�F��3(wP��n~��lw�^�EG�U)w����<ޣ	c+�-˪'��>h#)�Md��p��Z�%x��׈\J��%�EVŚ�r%s:P��Be�	Tfj~K��-��-m�.K�C۱p��X�2$
���6G-c� jΜ@�`�;������������,����a��h��^]�A���T���!J��vy�r�1�`w�Q6��=�L��py=nUˊ�r�9�/X`�vC4������Ի��3�c��C�tm�%�*�����D�c�U��<2|�K��]�c��-
��.�1�$�`�6��ѷ��t��L؟�Q�-����Ϫ��)�y� +5yJ��&V �YBkjO!Y�=�m	\+�z	�eXe��f u�2a:2�M�յr/z(�Բ��S�	�I/k����~q�����A~2�(@P�p�����+�2*�7�/fO+��:�Ӟ����Ű��d?l0�u+\+��-��LK-��"B��I�c�6-Re7<��g
��a�M�cZ��_�LE.:ᬩ�w�a/�IX�[~�F��Y���eqGw"���(�K1$F�&{sL%su�e���uf��ü��ƃφ>z�YoY)w�dF��3�b�M'9��e�
鍅�u�`U�5����=B�O7�����5r5B:*�=��9k9��4ըƂ�����������o&oؼ.X���H���Syq���L���Ǹ�k���3'y}�����{���,����j����;��[o�V�?7<K���"�`O^2� �&�\�	-�X3*�0�w��VZZ(:,����E9՟��	XQ^�!$�/g:[f���%j�뢉�t�)Ce.��4�lOu'J��Ez͸����U c�I���b��^B;��ul�	��#3ɦm�H�0�p�(@* 6�Z����E�e�\W���/�ڦ�G����ޔ���BjD�xE�xǒi�]R����:?��wnW�i 6�t��D���Myfڧ���e4��E�%�}Y3��'�T���³�o��n,"��_l�E=��::@���+�]�K譪G�ߒ~���`�35�_�UJ��Ka�)w#�k(Tx{���:q��wB�Ov`�!K
�B�>=�(��>D'xQ��!���B�Uc�������k)���u���ʨR��J�)��bR�};0)�	`nʴ9��J�Q�H6&�ȃ @�ks ���o��b�-��>߭M3�����Y��Dh����\[��� J���0��'�A&­�o�J��,	�T���L���84�.��Nk�)f��8�)K��i��d|�1~�£2�-��6��qօ�!vR�ם��%T�����-2(�S�'��OtO�ڗ����Q7b�{(>j���F��^]��,�V<+�O�W(���y�Ep�M�N0p5���M�����ǴL5D���q$�b͂k��@i�2>K�2��*��I)�A&[3ύiߠl����Q4+�Qu���",�Y��ϼ�A5��Tw����0��R�@	~�̧y����$`зo������9���o]��=9�u�tZl*�hℶFF
��1���k�ˬ�������(hR�� �z$�Ϫ_�˽�8�B>�U���o]΃dm��(���_۪iM����B���߸�*� ��>6�(5�J���S� �����	�F<`��d?���r���
�s��V9�_���7���i/sM���%�u�(���}�HT{�p�@�u�R\Ӗ���C�͕d�$'�/.�!v9�]- �m�g�I��D��
Q��zĆC@�n�%�,3�}�0�%[��E���E�x6�Ͷ�zw����]ta3�z/8�c�m=��jo7��V^7=���#�1� � �K��l����5�f��{���g��*�����g��Yr������fh-k�J�7\8�޵/��m���6���%.ۀ<����!�[���e��-��z��=?��=ۍa��c$BR0}�Y���Y5i����ڰf�}B��W'�V�m���,��8�/�Vv��9����]�����̊?�!�,JJm,�2�%}6\��_ɫk�C���م�i�����1X`!�mO%��5{���F�`�ELlv�z�C]UU.�4ޭ���xz�<��h����Ď�;.d�ԁ���tq�L�wEyk���t���iS9; E���G�4i��y̠�-� ��2'�$��N��f�?�S�a�s��5�Ԃ�v�p�2��7�?,Q��H�-X��yHM*�=Ivp�/�jGe
�#���YdM:�T]���Ru��i��c�PҔ2�8j�;�!��n���!�\����t�q���B�N���]��+O� ɀ�݃�;�&L�d�R)�m���Τ$W�t�jj���'�Yrs�O|3~G,�Pk7x�?��1)�Z3�g�KE��Ճg2�q�,j�i�E��^Ps��{_��K�aO���lR��1�}�"��*�<��~s^�ySkβ�h�}B���2�,�頝n�ٯz^��T���D��h/�!2�<�����]����0�����`��y��0Rڮ�`�cj����L/� 
��F'�Ӯ��d�*w|L(~���<��1\�;ی���+g@f��$Y�oR5�(ru]{�"RX�{��*��y�7�i��(���J7~z��Zy��}�2��;��%��� 7�FZ��Q���N+��U͗5��Y*�X��';U4�Kz�@ӄ��`A���?[3�'��N��g/ֹa��"�.|,�
�������d&��*�Y��q�NJ�e�5N�
�{���e�`<�p���A��Q��2od��'� T�z����]��)&)G)�:�[H�h�/����W�̓Io>��ա�f��x�ߕ�c|6�u�S���{N51�*��S�/�(���(�=A������r`T���&I����x ��
�~$�' V,��¦l^����OAN���\����	M�����7Ѻ����C�p��ìjj���y]}l:4��e�E�E�p)��{a��^N$i-�Q�GZ�-j�������K��Ho�i��%4��f#��2R���~����[�����v[�
�̃g�&T��c��0���@��g��A���j	t�<�O��C�#��q�����׃�]��fޜ0ه��.T�Q5[�����9�F�t���^s:�N�̾���l;�T���l�ٔUha'C'>[�:��ϭ��,s�:[V�Vie !�#�5���pP���lU!e����O�k�;L�|��o�{��'-N�5A�]/"Q\����z�uKm����;��7i���<�T�h���A&�A�@kD�Gy!��т�:(���	��}����rf ���[2
#�BK�*$��G�43xjU�Y�{29��t�'f�VSR�[�am����	\H:���`5C�J����E��@�l؟�;�R�Ny�����Hf>�!i��E�;�:�Sx87��6�f��1w3A��"�6�`��Ĕ z;����+���Q���B������+ݑF��6����*rT�x���7��u�b%����#e5;��8*�m�Y=�x�3�υ6�C���� ��#�HPĨp;�_�n�صn
m�v���)_j��T�ی���I?�1���Q .���Ɗo�'R!j
��6�B��	�P�XV��,��Χ9�C<�����m�� +m�b��04(X�4̵��{��1�O@�LPup�<ޡ�M�b�]����T�Fl;v����O�Mj�xe�GԄ�F����ƣu�sXn	���6�Z6��E�´@��w���'�����J&|'*��Ҹc���~���86} $:xo��7�8�k$���C:_�Z�%����PN��V[=�Ʃ�<���оC�S��>@��_hI}���5y�6:ϝ���0'\Y]�7!����u�B�|q�2�>��lT_���'�A])!�O��Q�M΋q�^�@p�,V/������LD��ǳ��]6��l�gm�����7���0n@��5��ȅ?�sf��^W4�5�B{��7ŧ�C�P:E4^���@�O%���� h�fr�He%�sl����9�߱=�ځ~�H�|����pw�t2�om�HW��'(��cp���r�L�H�ɍ��IV����DC�!�g0M�������5�0�N|�nK�d[��3]a�ȾWg8��q���!$Y��_`:AK��L �z;4��_HүJ��F�k�ӊ*Z�����h�P��4�e���,P��<��S��\Y�rk�y6����zu�3@L�"��`(yX���SmO�
P^u+�$���;;d���g��}�,�y�+4�\��|?=�3���;��b��:*�dxX����<w��'f�"�������?o_k.5�\R��a1$�R0��o�� *޾$�y����k3��)_#��+�
$lsc��C%�y���j���T��R9#�d�~
_����;�!�c+M��<�,	�-n���<N��8������wң}
��<scF��6}[+�>< �����@�2@�y�)�_�5�3���5C�d! h�P\�G_=�\e���	���:���/N��9����(|�/�}y}J�&�s/�D4�ȅl���s���O��#[�Ϫ3�^A]l4b$��'��L;��FFE{������8�W�%��ii��	�t]�ZqSM�:��/� :8٢��x�t�n���A��$�c�|��G���H��X/;�ܯ���EC�.�м��/�BZ��!�k�]�˭og�ʙ�U�h��S:	!l-�o�ui�!��{F�C�����k��}���3�~D���XE�^*ӕ�ӪV���5%� _v�J�	��M­S`Zm�/�y���seckK��E �0���Xt��W�z̺� ��X����r�h��T�9�3 =�&��m�X�Q_N��b�d@�&Qk�*�)��u�X�j�3�:�w�}&�'���9�k�s�V �@^������C�L�� G��&�����F^��#V
*{�Zϕ�ﳼ�W�0?�<��-@�#�ԓ���ąd� �?�To�~��N>�F"�F��_>vL6C�`f��r����ʛ0ή�#�U����OwIk�����G�ƫ� �~��?r%�A���qb	|'粮;�"� � �����~C����7��:Mi�����RZ"3`�z�U%�nF���1�R�)S_�O�x�T��˹=�~NMkC�JU����$ ����҇��=���8.�G?�3�@��-$m"�h�u�"�V��wG�w�$����ݶ��~y6���s�I+��s�P��^c��_=u��O��id�c��s&[y�l��q>�<��kt;7�YU�e��uː�GŢ�������U�)�$�0X��W`�m2L�d*��*�������� c�t%&��,���3�z�O�����&��x��;C!~��Զ����満�Y2�x�!�G%����t�a*�W��ѓ�-dF��Ʌ�࠵ �j+���;�v8d��fce��.0�c�4P��wTJ>a<<Ҧ�'�ճ�E��}����%@���5��R^��&9[��z(Cᑆ��U���)pf�5�v���B��:w������I	`�s��v��~Vu�$� baV{~(6�:@��â��y["��B�d��<�x���"��b>��1L
[G	u�q����L|9��@Ln��%���"s9Bk�tl~�2,d�@��*���]���6�X�h���st�-SK��,�TU��`Z{�u:*G��[�����a
�PL�-G��n*fLp-�>���z���}}B��0�H�/���&,'>>/
M�[�޾�Y�����	X�H|B^��馻Y��io%@�������(̨��23�m��o���I�oMA�y����!��PE�U�[�����"z�Ͼ+��RH;_�����uTHB	�ښĉ*�fk+�I<"��Qq}tks�6x$uh��6Wq�-����J����?�A�TN��Cף�p|����m�N�weH����N���J�KK<2�` ��W�$jbgm�+�H�����Ŷ�Wuw6"���K��8��'��} �YDLd��������w�_HL2�t�f�T�zCY3��QR�ǻ+���36w���Ԝ�zqq�d9�/���6p����S.n51������7G��w��p�L�����m8�NY���f`�T���y$k��i���?t���p]�l��cIU�PCKlvLŢn��t����pj�*��HJ{ �A>u�5���9cG;=��@8��������Jk�����h�0��Hi>���6�%�I�8ʡ��$,^DX�/}��Z�dƪ�T��k4@�}#�w�==�S��<4��N��O�U\�Cs��
�J<Q~�̠�V�O��ͤ�N}]z%y#���)!�-ˣ��y�YQSϜ=#��M�61���&���3X1��s)Z�TG%�ܗKi('��&1�y	2ei���R����,0ϥJۘg��Ҭ�{�Y�Q.-1��w!t(����3F��kK-���_bY�>i�fhJ��]}��8���ݳ*��y@���ACn���o�Oھ��~��
��� �ԟ\��/���g�>P	��qoBg罵���W#c$'�Q|��R�'g5��գ|��>$�����ău�몜��:�G�.,R�Y�S4[J���w�)A&<w[��ĠOMt�O��W;	���6��߿
����Y��FZ7�˨�\3��dj[7�k����i���}��7�Bu����. �]/�& i��	h�� N�>7���{'"f3��wH]Bo��̌�� ���l���4�"�\o���y&f��x�,]�.����To>�~ڷJ����Ƥ��T��X�m��F'� ���gzݒsi���d"G���m���ͷ��<��x({�e��ME�[��|�YF�4�N�'G�B�G�Bb���>�$�4g̅9fwLE ����}`��M}a"P����f��k��*[��̅��#|��"S8�uj�D��4@��;!�����e�1B��$d�B��*̡��k!&�aRӣ�����*�A�X�X�+�Q�0�V,Qs���d��B�	4�]���'Mk�g6K3� ���������e�)}�}&K���2=��Ȟ�t\��9B��-�Iɬ��`k
;� ds���c&�͚����<9'lC�?C��)A�E�n��{{toՠ�=�ʃ��&�PO8Wj`h��O<\D�S��?K.����/T�f$?�)p�.��R���(�4�@ǚ���S:S�U��
-E8�1
�%��yq���mev��"�y���]�n� �z����\�(�ʏY��j]����A�U�޹]�,2)�� ��F�?B6a������7_���G�s5PyS����sG�?<'4���ӷ�u.HTA�U����<="A��.u��@z���pp(j\�Z��U���>�ɥ�e�YHRc�]��{����B�TO�=�7> ;�e�9��J>�b}�9g�H��ۈ�fv�,�Fzv!��O�T�<ɹ�zP���A�[%NQW�����C<�:�K~d�_�/l*�"�2:g-Ộ܌��%Kf$��c�]�N�E�*ں�Y<&-<r��y�dQ7M9/)�@V������0���+9aIӼ�v�Q�UH��;OC�&� �5 �u���j���K�)����!��>Q�#?�7(�Z�m��ю�Dc�ʮ���S��)�E[-ʃpÂ��d�d=�ט�Q���|K#GSc�eQe�BQx[��7s2~���(��&�������9�ǥ��N����C��n��c$�U�bo�F/���˫t=-�wIܞ���n���R����b�{j��q(=t;��jd�$�	�V���~l�y�oz��k��<��c� E�ݏ*��w6���J*@���>F����7�/�P� 1�����84��TS��9Gf$C)��0�$���d�Z�@!5C�nI�Q��;�QJ�A��eǾ'0�����|���I���� [���i2����r{�
��[�H>���3�?��8c�je��C0N�/����Cp�1ee~��M�/��k!cb�UP�e�W[C"H�̾B��}NtN?�|d����i��3���*���7��&��
:���R綦N|��QSj�8�e2g����/�cwQ�`9��tأ殻��^(�9��ڬ����PqK�|H,ӽŅ%�%E\� U�8
+�J��ۦ��E�B�,�m�m؊I�-!�u@>��%�M*E)5x�RX�Z}�(�~kW/?�z��MCI��Phԗ���_�x%L)؜�?��7�ay�)�&����n�:����W9�R'�6�4����֧�վ&Y�o�#n3�mG�w�3��a_�׭Z�H�C5�K��7x�_���D�w��S;$~3�G�\Qm�nVN�K�"%�А�nkGS���Y%�� ̚����|V��5]�=����e�,��`8F�֋��V�c��`Re��u�گ����v*I�
��!������o0-)py�o!3š�6V�,1���+'[�f���l�~����n��C�wO60}9����x��G���JP��wZci�{����jmq�^��<��Qo\�W���e.	$������M"#Ϭ|��@��J�{E�ʏ5r����R�y��xޖ��X��x�PF��,���f47�Ž^}��3�F�H�2�9w���u�u�a���}>���s_'Z�Ҟ�H�P�M<�'��� ݮr���k� �&�	�]ߩ��O�$�c��k��}�t5�����J �F�fhxC<�dV ���1�"�����&� ��	Z*g�O�QW�N���ƍ��VB4�]3ieqV}�	����j}�>ݎ�Ԛ]��^k�,au��� xxH"���Pk;6��cJ�����)2k(���+!��]��ȡP�
��L��K'+��A1�R��)�����:���$݌�ݭ ��������Sq�F1���$(B�H	)�c:ѻ���G���Si�_ȫ͓H���6#�ȟU�����	�*]�ɬ0�h�#�u��EbN�Ԧސ6�V�8e��n���O��>�*I҆���n)�p�{�ҍ�x��t	�� �7�1T���Ղ��.��VT��]=�M��x��o��x�[�ɽ�>H@���4CЭ:��'��g��C�N{��N\�Ԕk������.�'�,�.%��G� 뚠�uK����(m\����昃kpf,�m��v��N?�9T-]��%V���D:�^�"c��.������PS-�2�������s������ݽ>��S3w�� �̸ּ��G0���M;C��).)	�y�6��d����HoJ�Ls��vx�S�\b+*ܛR�cē��O[T�W��i'��D���4�Mj�`��}���٭�z7��2�AR��4�����B�?Nѫ��v;0���^x'�eX0��u�j��W_ ˬ^6zR�t�{�����Q�%	O��I�4�H+��ȹ^x`��}<��B�Y^fn8-�#.�F��=�!��b��:�c-R��v�W��tg��9{���4c�תߙ���G�?���es���=�j���R���U`�
>NQ���#H�Б-���ܙ����� ��;kϠ�@#k_�7�*��F�H�>�������C/݂?�Ļ��8W��%Ǡ%��.:��>�T��B$�@O�"/�y�����L�v�gi4�Dn��͊�p��L,\�"���c���4��ָ�=�A7�hjX�_jz٨t��m8��T��%��+�������m�bm�~
��������3(�0��V������� /��o��@R�n��t���	��fЭԪuB{�Z������P;£��SGŀ��4�q�6�R���m�n�x��蚩i��`9��h����Uv��|_�]~��R�q�o�3ǩ3��=�6~-�@���/^׷���=@�l�X�oĬ:��м��6���p���X>Nbz�2��@���n��Z�������c*�t@ȅ	��U���w����
l��Pg"��oWI*!��)2��*V0͠L�O�k7S �6�����,k����WP���(�;�?�9<�!-����'f�(|�T]]��45$��f��l�j
��;^B���� �;EE(v�ݫ��X��͛^clTPY\���^�v'+_Y�R��Ij�a$��m/�+��ȿ�n�y)��k�Y�WN1�0E�?��'+D�ygm�A�E:=�w���-}�� �0���F�MI�����W��r�I�rw�cF�%�)ً�1'.k��jT쏇빉GD��!�f���]>��婠b2S��%	���wb�,�,t����N�3F&�{@�+��㨼=.nϱ���&Р�q��'��/�HYn����6��N���|ر�l��<�ܦ[_���'����^'{�mO�x��fޅ�΃��dR���EThc.s�y(c���$͸H�;CR��&iqR��*
�/f�W��E�c�xy\�@�&�_Y�r[V�&�4��W��d�J�{9,4C�Rr)���Y-�(	=S��kʸl1��vM��c,��]���cƸ��#�Qο� ��?�N����ر5�2XIt|�F�Q�Z��{��,d�1��vgr�@ǹ
`�/�B���Y�;eł{P�r�s@-	أp�Ű�|���B��|��x��ʁ�g%�S�w�����`��Dߕ�d��C�~�o^?V�Rǹ�Zs���0O_ڞ^s�@']��^��,E�s�^�>�0�
3�tXq3*�{|%K_b@f��v� D?����B
1��,��üc����b���≧G��'��#a�!Y��ݛ/沄P�$�i� ZA�E]�_3��
.�fIR�c���.r�<IΉ4�E�Oǩ��i�,s�9u�ȧ��˩L�)�d�ܟ^L�ә�m*��ʓ
���lc6�?V$S�к�v �����x8���r�%�ŝ�H����
R�^���d�e� �>v�K'���}A�*(�;G4~ �j���o��\?��[0p��8s�"�R��s{��,s�+���r*LQ��V�����~�P\�w��TSӃ`b�4N�!*i�Mx%����5�:ych�����dGG͎4pܶ��/�&��N��\��۹�@'�lD3�0�������{�*Ge�%o'Ov���
O�Fk�f�pW"1��[kZ��2�K�K���ف�z����!z�[��F�dE�rް4���&�8�UN��9Z�q�-� m�c c�Z!їM�ōa��pS5����8��s�OL�W�
U�4M�Z�V ����)�`���?K�_�̲Z%t�S�6K���JpD��Y~HQ�1��2��0r�EoH*��wI0KN}���f\��A!�ۉ�Qb�(���)��K;���>����ooC~(�W��ne2R���k��3����it�V��sa�J^��"�`��\����U��;�^^~�<A�`A�$��q�K�N��~j���b���|N�&f��C���i��Nkż҆�������[�K�-�.hm�V��D$�������J�Ϟݚ���ܢ�I�H�M�D/�����yG/��a J5C�M?R|S�2�1��tQ.S�3
&�0�w_�ϯ�;����J�/m��r)�EK�I��4i2h�J�VOB�W��*����_��@�v=�3� �]/�޾ǫT�w:�3P8�ĿB=G�<e�	N�B8|���F��~����Wn�t�J��g����I7#��l.}��=�K�z��y�B_߂�d�-�E)+@�.C�X:,D�*�Ϻœ�N�������v��P|��(x[a�f�	n#�����v��� ���b���j��pʨRל�(�E�;��ͥfz� ����@�*U`$ ��S�yQ	3�3�_]��K���e��^`Q��[��\L� @�7�8����&���k`j�j�!��u��CL�vP��A�+wS�EV{g�g��$.�Ǣ�ÕJL���"�'��Wߪ�nkyI��ԁ��.ag�ᥛ�hdѪ�7g7�R?k䏂���S����Qj� l����Uj��I��=B(Q���Zʛ���K�ӫRk��_|�v!��(5�}� ږ�� ��TRg�YL[Ve�bz��l�6�|�=�D�3��64X��D�B\�2���ك�/�8�u���mL�
Y�����W�˾�zf6%���+��A�:��_O�?'|���<c3{��KDwF���~Aǹ�wO�)�"$��E�"��	��Ƕ�	��϶��������5a*�����"JE�ɪnc9��Mг��!���$$��E�R���}1�+�W�����T����oL��O�`ۄ�ۈ��LI���#JkTf벫�`mg7�ho�c/J�<�)�8�ά�ѩ�N�6P3�^EU��K{�i�sO���K�ܟ����u3ӎ��u3� H\�❉�/:��&���~�r?`�q6$��/ ���
����|�Ww�&��11��hŧE΅�Fl�VuQlF_��#Tu�{�/[��f�kOb0�j�)u�\��,�~��%o������f��<��jW#oDL$l���5"b=�S1��c6�N�~�>�P���|4~:C>��J�CˋԊ=$��]��SJ�`��ע���l��6����2!�ٙgffiߕ-&	1F�_�nb���:j�r�"�EA��i�X�P{i�3�*:��s�����w�,�K��Hi�bт����b3�7)ﹳ����*4�ׂ#�����)���;I�����������{�;�`x@g���Ӵ��t+��5���랐1�z����Q�������@�o8aUڥ�M�z^�?����n�0�5���Rq{�V��o/T� ��n��Be�,3����1.C~���/L�ZB��nn[�N�Se���q�s��0c�,�i���	�",sƷ��_	�����_����s���-%�����n^�$^A�c�������	�w���xڄRG�)�(���_�������+*P�ϫ��v51���""�aQs�r]�N���L����Q�cqwB��b��~N�!��PɰY<��-���i�r_��KX��T���aC-2눚he��ciж��
M|˝�@����!��S�j��~���āV^oph�H�˲�teTB��_�(�_{Y��(|kS{�.)���T�.,&C��D����Y���s�]�oG����������첓K5J^�ԗ@� (�����BC\����ړŚ�HXLdć��9G.
l��2T�?�k��n�o�d�.qЛ_����a�E�TA@�.#��'oqGV��e)��1��N�r�m��L]Z߬�P		��}�Ԭ�ր$�T����{q`amT�5�K�<��,<����i������1�K̑���l�בH���ƺwh���QU�������piׄe��|�O����� �C��ڈo�_�1��g�و���H��~�����m$MFf��G?+R8�2���[dŬz��������2*��d;>�|���v�Ӥ��\���I?�l�5�L�Ў
�)�q�m]A��G��0)�������m���h��.���玱]/ZUTJ���`������@� %�<�%�Q� �����������������G�LG�k4P/�:�-s<=��,�2�� �_�����<�K�"���Ƅ��E��EY��`��~W)�Hy�W�&��5�ug,�����u�<[������pߡR6�В!}~��nf���~AR���`,u�🱏o>��A��҉�3�\��%���xX��yM�g���_���D=>���-}m��*<�X8&% u�#$�e_#�ݖBeV{Zrk��ː�%O�T�he5�`��äI�����:�8��΋2 7}�Ine<;���'� ���f�I�@�>�D�� �Y<�+!���|Jb�6Q"�������e`�B�?*q���th�d�b+�@��]��( yi��V�O���z�W�U�Cx�|d�� ��Ѓn��=�V�[(��L�2����&t&	�p��/W�ט��j�?�E��g�
pW!	 vU�S�8�pX��jpFE�4�:���C�z��R�f�sq)C���C#��~�8��ut�������Zr,�e��Ǩ��<s�~�MFV����&X�%~
Rg8C�
6�ΐ��.Tȁ4+�O�S��ٸ~m�	��n�?��-�^݈+�w]�����F/�_�!٩�Y-(��0�ޏA`Y��
e ���~�	���T��j,q5dZ�$�[��������+�N��p|tP�����U��zb*���!� n],>���7��VM%�����0�t���Blbނ��M�!"�we{Ƅ�Y���۠kui��чR}◟r�=�c��Qx@�	�0�Ž~A�����1#U�FB�T
}Je&fWA�ʓ�����S�f�L��>�(����(�b�x#e�Lc�Z�{�(����U�6���P�e<��Y�E�u4D����0!\Ua�'P�s���&L�����<��X{�Kuy�lҚ�y�F��e�~x�edŰ)�5�6���|��U�<��T%����6��8'�n�\��/mU�}���w���R������^�&ٍ�����6$2,d�թI�"����>(��C�*y��q��ED!��P�^�S.��M���g�a���9����A�gD�C
Kel�<~P�,�7 �+����F�c��J*`��!ĺ)�(%���.�3Qx�* 	N�.���6q��,t��6:w7?rq�fbhf� n���\o}�:���B#ބ���j��ߠ���Y�̶��1�J7 ����Oa�^�,��oR�P>�F��4�-�*]�y�ě�����jz�NVx��I|�ч�g���ow�0�9.�����z�\��*�SzRJnuv��G�x.X\�#�N����xf�Q�i!rY��,4�u�ڴk�y�/j��D����N�-��u�8�ټ�>����+&���9$�Vĭ�)�N�a�q�A�ZgF �ح�Ώ���|`�T����N�N��SX?�Pӵ�Q�I�IP��L���(��QW�1�r�����n�ԛ�{���{kAg˝~�Fl�Ɔ��_������|�� ��j�_�v�� ��!i�p�u���N͡k�H�P�%5�R5���&��D�����"Zw���N�|P�� NM��?�T{�����oc*y�0��1�i��l��tc�2Ra����ˊ~��z+LI�7��5R�#,};�lW�	uu}��Ov�w"��wO�e��Y�\�'A��K�(C�"�*j>f�9��d&5Z�X\vV�i`�?�p��p,�$L��n��"�#I҈r�4��D�D�x!����!S�����ڣ�Q~��{��_o�����7F���ݟ�.T]�t,9���K�,��C�q�yQ9�2�ؑe@ɹ��e`g�m���_c%!�F�^ƨN�,��/2�}KI���y�
$�i��R�P�>�n�NWcEiw%�,�Vo$\�P�!k.
7`���<~BvԮ�(U>���q'B&|6���e�Y�`I�>��-e���Y��=$�:Q��j>�h5��j�����dt"^�T�-7�#��޽���	#* 0�YUs;\�c�l���S��'Tj�ڠ_R2pQ6�h��EFjLcDsW��_nv>���CAa���e�����QT������n,�0ؽ;�fi�Ib�\N-ҁ��Fݵ������M�+�>�+�/,s�<<�SbImΜn�zg�H���kj�]�<y9)����5�?���05E���}�EB���B�{9B9�W8I�4�.�����d��1%QqIK��J!خ�֗QD����D�~6\^9/�!�؅��yQ�ot�[��=�g������>�Ix��<>�4��0;�n���rݓLu�i�7O3�GY�!����+���MR�/�d�n�6���L��>?�ۮ�� Т���?=�1���#H���'|���/�s�(��!a��$;�#��~#��K�_��4�}��0�� �T�na＂/8��aZ��(��Ղq�N�d�����aٛ�oA_�cp��j�;�[�)�RWj���
K޻1~E`����W�㓙���Ê��0��C����m�n�?�tr&�޹2\�-R�2�)iiH��ѡ�X���^����&�r�lL�_E8{"�'�/B>SX>��w{����C��&�?��/F�n��[=�A���	��؝��u ��3r�tR9�o����� �=PDs��w���w9oݒ|�s���ؠ,l���9#B,j���x|fEt�Sl<HܦJ��"t�ӼJ��
������y�؀8
8�������A�; �e�ὬN�'�yb�{�%64ʅT�M�k�^�N���*�)lL�wַ0�<U���q�k���&�0���w�3S�����{	�̵u��E���Q6�<QV[�*y�V���[QXH-T�H��s>�,��d��yߍR�^"��+��m* !�C�`g�r�F���UsSB.A����P��D����ziX�u��Nsڅ�"�>d�+���s�fA�O	�ٲ��c@C�;�x�>k��~q^�N��I�TJUl��[��+�@W�������&�E�{���ۧ�Ij���Q��m�b�ʜ�\�".Ü��<��M����팎���mf�#~�����(:Fv+i4,A^��9O�y��QW]��Y����'B�JEؕ|A>�}�W�7BMᙥ���96�9kx��H�{ϴ[ݟȃŠk�߱�r��K���`���xK�B4
�էsmlh�?�Ȼ+[wphS�|�,��d��܉%;�
��7����D�3���t� 7�@W�ۧ�;xnZ`enİT�6�П��X��(���O)32��li͊b.�Y�U�G"m2�<��{ۿZ��J$Dl�w�uR��B1����i��s	{�H�\<��F�X<�|)��{�o���hx�K��m�
qy�9{�ٲ���B_��?w��_�`�'q����^�'�,��^l/��]Rg��'�(����H�=oN44�ۨX��х�w80�\[`?;�S{�J,�1�N�x�sP#��G��N�����;H�m�Έ�=�@l����'g!"Iw'������^2��p��������`?� �E��Pl��F�(D�� �l��l�h���# s0���!9�t��4[����	��i�k좢k�qP����O1&���:�[�ऒ�A-H��t|X�ϒF�Z{RxK.lѦ�N����l%�3:@{�xG��V�v��(�d�(�T~>�:��Y�=x�����T��Xq�z~&�ٌ��X���<~v=�H��g�$�6�|�F
`�R�I̍:)���'�U���J紺Sy�Z�!�!�l�(��B%=�D���S#�G�q�֖p��fR)��� �9�54!�.^�]�2w�6$ !Y��B��B�j� N�U��_Od�ۂ2�u2������1�r����"��r� 
��+sj��?����`(<�q���cy�?��s�V�;�i��u�t���x�-:&��=G�(0h�������I�Р�ףڝ�$��n��]�6�L�.���vӔ����]j�AO��F�̸�x[��9uy�W���/�~U�����H�X�W�P�M4��@����v�>�:8H�z��p��0�]�a��EC.ʪ�ے��bRӓ8�j��v�liw^a.�Kx� ���"��W
�B��g�z[���<���Ҋw�e�r(w^���AT����v��|&rV/\�H:��A|�Yj%fy_�D�ېk�m�Zi9g��2;w����Oixt2�Gb��f[�_B,ߖ���=�-<�5��E	T��qO'I����	LT����NJH?#p�26Ԡ8fi_�C��x�O^"�se�d9)���\�_�=�G!��|�}4��6YE>���ʋt�i �ȟ$�z���݊����`4�-�p@�.*�)vx���R@Z���QM�	e M�A�_�)�^"�7��F�Ӄ���G��P����e9J�������p�/��=8]!W���x�]z��V.�)�������W��b���'앇��n��ZЯKn��@a3�G<|��9Ȧkb������*�z��ŷX�y�u9�U��w����a�q���y2@���j	_�߬0�0�+c�d����>��daV��;����62�ci�~��kF�x��T�"�A�/��,�l�����ǣ*���k�8w�3� ̓b�{R�� �J���O(r�D����K@�ΟIՌ2�4ֆ��G�Pg��fX��!t�뱵��?A���K_% ���Z��+���l���;x�����4-r={kDQ��B�����4��k�m1H�Ҹ�G�9���߬?�j�N@G�&a�n�I��l$�@����W4P�'2҅��IE���F�S��9�i�㤒�`�V���Ym u�X;]7	k�������SD$�N�]�1>�+,9��h���4`XQӗe��v�P�*�Ld&c��]�vb�����+v�� ����v5���upv��>
.�)�bn!O����W�����H�o����$ym�=+��#f�:tod��s�勒'(�@���g�~�򰨷Iv�4�W��G.�f&�:d]"�ϲY���W�'Z9��A���Im8,��6��� d�o�ϣL�7���I<f�;{�P�$�+4�F�q�d��/�v��N�Hb�\�]����T�f���x�ӽ�v'��z~�`k��g���'�����3 }H�2�"2X�~�ޢ���&�V�h�4u#�!QT�<���*e)5۱� vLk��5�ů���)����"l�D�v�#y*uynx�Y�C�?���4pw�'��9�@$���.��@�R�����<�B����N��As+`к�M����vH�T�4����y?��lΎ�׭FDǂ77`P>�j���f���1�����S^�8��8|R�_;�.o-f$ɐ�p���W��M'��W�ɭ��a��:s\f�6��\S(�>
��׾�S�G��k���fjK�hɚK�EFt���PEˬ�X���}܅�?k��3�/�2H�$���~�$5E*�C/DN�H�g76rU��U�f�+.���lH�vٲ��C\<�MKS��q�9Z�I��c���SH�v,���ޗ��2��o4��"�\���p�����3Nz���øqeZ�Ƚ3v��M:��T�GQe��sU�S콶[t�ZUU�5%�
�E/���Wj��l���)���Z��i,���^�=�*�(�ֱ�F����i�k%]]��,���(�RDr"z�6|[�t,���TA���䕅&���$��^�J��2����P�\y�f� ��}�~$]�F����u;�;�q�����kto�鰽��RX��*J\�8\���|�g���@�
�h��K�ZZ�f�4�	�d�j�2z���De�HKde�V�V&�v��׉-�W�o��Y@NF=��Fg�I��r��Z����qyPp��������r����|l��R��ȴ��p|���i^n��V���F�3��{aR@s�����70D���D������>�^L��J%H�0��z����S���J��+�rC��u<��"�ܽ"��T�&H�+��h.,�22�*&�D���V׍�,8o�Y�����g�ףS���Y�}���A�L�����|O��i�s6?����$�a,z�5̒�a���X@Y/ңwD�ǭ}漴�����tɩA��.n��D-.)��j�4��3��,��(���W�6�7���V�~;Ĳ�=�_c8��>�+>���W��:�ſ��/��6-��z�Ƅ\(ɊF,a��)��v�����f(�ߍ�	_��-�������j���iy[�_���yR�+bl�P�B�>m?Mn�`j>��z�23m�¹ۓ��q�%�^[t�\BA�!K8��gl{� �ܩ��&ݱ۵T���o��>�0�U��y��.�T�#��e_�T�f/K���~��#\gs�:�}L��������~(i?��Ւ*ʒ9=U��}������n����r�љc_����~0����!阇 ��6=I$i���T��8Zi2
�y6��\ҁ���P�f-v�Z�^>&���>ޕ��)c�2���9�[
3�(pA=�w� �غPᮋ���1�U��3��;�
���2�XQ�ޅtq��kd�e/e<䞁��`㲩���l*D���0��ƿB���]D�McOS�"ܝ����&�8��U T�v.���"w�ވk�*�@��l6��bkP`�q��
ġ��g��\�|� __�/�	��!-RS��a��E�^�D&,ԭ���>0P��&;�IiR�ūb��[׺U)%d���eU��)+Y���S.Ś�]��ĺb�T�r�&Z틠��T��я���ahIU^�?�1���=�7
���H�x�[�z��ɣ�G��aϵ�S�l;���4/rώ�V4���}L򷧑 1r���.'?�V�.Uʝs��P��pz�ۂ�mf]K�����+'?�~�vf mں���rd� ��S@俳�_�Z9���)����T���!K(�?�Ҋ^㫭4|�J���}u^��\3���h��B%�l��ى�f^`ф��K94�8X��|���?O����^���豯UE�gS�ى�%6+v�;}��X��~����i�\T����CeVY�����o�z�i����.�yz��+ٞy����+��XEnz~�*2�z���̎��=��1��f�Z������,ө	E*�7=/M;��@7;-Eb����I	�Ǟ*�~HO�fs���r��ȳ�e�0�v�p��j2zl�^��V?^O螮�C��ؔ�5�&��8o)���Vwh#B�AAc&�X]���E��Z���x��\f�d�^�	(O/�=�Nõ���C�Gj��� ���[
i|��!\*? �0��:K�����y������|{	���)%��q#61������P��SOP��S�7��*��Q��YK�R�ļnz�V 0YC �������d*�7����{��n%AN:=h���"��w{�1��Wlk ��~����۲(
:�zo����Nd���]�8�`'���k�x4@\
:@�=�k����7�H��)5!.Q�&{U�9_��A�mr`h�E��	(웿ٹ����	�j�˰mL�X�Ǘ�����$��h��.h�%��>�RԡL�l�A�P�Wc{d��SsF�X�����M�&� s�˘7{��+�*p'�w��]-ɐ��p���ⷁ�n����-����FP.f�`O�vV�̆��$�ko�������.��2�{��d�~�J�-��* �FlC�e'�C�,��i���_�,��V4"حHj���f�cBy2s��n�bu����&�2N�ĸF$����9vL��п3�7*������q��u&V?�n!�0R���csP�67��Ez�ҥ�~󎨝s�/o��������`����	+d��X���T�ː�0]/@���Ξ�b��m�E_}o�n͖�!��e��4�!����uxSpEZM�<P��5����
��&u��m,���Xs>�`ނq�P̹��<V�_Yw����ǔ���)#反X���*Q�p+����T��`���OΤ,�$���1o��>�M���
���m�qpC�D�w��ğ`�ɟ+J���I�r��d4���
,=F�S'�dW0jA}S������'"�ġ��t-�ɑ6ٚ�Ce�rF�/{�����sf�L7�	E"�1a��;�ؗ��U�	r�m��/���h�I������a�SD
lX>�n��-�vdA������\}��(�2�7�����ش-���Sen��6���pJ%�D���9ߑM6c�*T߬�js8�2Rܨ�l����)�Gk�D�,�G t���- �~�w����y������z��HXZC��%�/v񁶎Q�#�$L��� �O�U�dl@Y�-pC��K	���!g�`�YE�O��4����W�_+(�Z_'	��[�m/�	�ܬ�9?�d!e�f	nϢk"BQ��.��AFm,r�^}P�!Ѻ� ���L�8b���TH���3�i�`�i��[)�N�-�V�e�y��8(A7�A�\����� �$0���5�/��=�RwN���A�M�3Rٙ-�����VEF;��5
��	��䯦NC	d��[\8h��5�nz���ks{J
���=�������UP��jˈ���K
1���8u=|���Z����&�t#|RjA���}��R�������!�f�Ҍ`zd�P�	J��$4Z���2)�}q,�H�v�(�ON[>^���0��4i�E����Qmmm�����"���G�� �!��rnדZ���=Ǹ抨�9��x�䌛$�K���
CW!,;#���_����AÚ�C�+A�@�3��)}��GMUc�Ӈ��6ҁ��6�׾�CQ���Q/?��b$�&�VU}���o�L�`9���q�S I%ݝ��T_e)�'!�0���TO, ��ޝ��46a����.]�U=���r���wԷIu�$L��}A�C��A[GྲྀJ���ޏ�IFK���-p��bq�3��C��[��)��ݨ�g&;�g�qOʱ�.qix���|Z��]s�O��;ǹ~ �������(hH���g�}��o�0)z�6?�f8@����\��y��Xި�b�4RYd+P1Ct2��jh!D�E���k
Ng%�r��0�S������w�UP��Bu��Բ���������^�E�D��ռ.�� �y,��D",�e�J�	~��s�M�_�R̋E<)����nθ��ˍ $�8��R�a��C$��X_��n��:�R���.�"���Yo�.��WS�!\��AXI혩�O�YB��?��C����"�����$�����]�%wuEV��*[C]�*aM�I�nΜv�{��&�F�U�� \�9Qt��H��ca)\J
]"p��e���誱6�d�hT�e�4iB���`�f`�5�e�e+
 ��׳���$��8V4`�2�h��ʭ#w��/o��3c�g�ۦ�`}Owԑm����c�����ʛ�;��_.�!���6ү�:�(�h@�W��/Q���=��a�� �hWҎ����)rS�����ӏ82�>���N���F��0���qF���W����W`ؽ?�OI "'E|F�a 7�Y�[��ـ��Kie/E�5�V����s]�ij��AW�[C G��6<K���'���
l� �&a9����#�I�4����1��I�5�1��xr��	���,��m��:E�(�3�������鼦�,�Cr-*6p� ��5��B�|�1&�K���$���<�jE��!�n��_C��D�#�m�.�Y���<�.@������D4}R��ݒ�5h�Ki���DS,8z��!���>�=GNN�@�ڲ�`F�j6�����vg��N),�Qg*��U�����j���_����4 ���N�_��t�A�1��xۉ"ş^=X���p�Tz�2UՅ�\~��
���<v��L��pVeT7ԕ�箫�Nn��u��n�\D��$�������a�]:?d��2*�(��E��m-���`�(��!ƔY�e�XY�P� 8~��]��8;�&@?� Rf<��͐+��ZY�=$OB�9u�MB�5��B��D�M7ܘ[F皗Tښ�����|E?�T���f�����I�ӎ+Ҡͥ���[#ü���E��;{�@�!u�IAC���u�y�=����J��kB�+Oū;���+C}2J¿=Uz���$Vn��;<�3:!���1����&!�'��2��DS?`Q@��)9[�����.*�ƣX+�*�#��&��b�a��&�Ef���Ω0�ah����`�t�c�o��h3���L�=(wF�&@�]�;\E�D�ݬ���P����Q-�e�^������`��7����g������#�*g��^m ]�9��"S��%�W�]u��R�_h{�ʹ� ޹5ŵ�fA��!Ră�ݸ3��/XG�UY�BV��uO��r�s�).h|��K'�b�JP�ka�-@�T�������\��he���Ú�U7V�~�#]��̀�2T]zL���È�]ӑj��V:)J����C������.�����y@����o�8$]<0)92�qs!>�Iֽ��bW�?����WDBo�h��,�f�#�����U��*��(���DjyeIE�h��x�0�|0�0���fn�Z}1�vg@����.4����i;�zV�XͱO�.A�'������|��n5-WD�΀C=��|��SVq�ˁ<3�����X���ls��[��ȏA�����+��kت�e�8�x�c��8�ʜT�Qb�.�.;_�q
Oc��N���p'}��LX�XS�K��8�,7k&��2s�&��,��P�3k��!c�Lb�o���>�f`��.e!��D�n��}Q��);(���vI��S8�cI�9��Y��H$�ڃLU+���I��0���Jq#�.'. ��+-���2J<�(���4� -}D`
.��{��:[߶
�P�w_e�4�"-�v��m���Z�Y|�����W7L�\�A� �/#�g�ൟO�ڤ���I�*NJ���x���~%��b^��ΌV`i�2h�F�}�������KL��l��N R���3�2s@�>c�S�N����iBw�q�������>��US=l2h���ݡ�2A�����v��9���O��z�h�ACj5�C嵪�@��>�R�1��f�w�	��c�v��,�}�e�C����`�-��d
t�;Uf2&�Β/y���.i^��j�>:���Mv-΍�u�ybx'�kC1�8Qn��o�2�8��6�h�����/7���v=�������@\�+�eE,�OT���ԩ5�JNlR�q�?y�H}z�`��q�K���ː�*����דy�p#�V�¶[oK��bUY�yMV&{:�t:�l&�_�!�$V���[� ���$A��&�Q���R���ss��[�!��1��Sǹ
�@�ՒV�_MDo}	R2D��q�b��v�Y����S�uP��)Ջ��H�)��pB�"ލ���>o2��
8�"������=l��f��[�3f8�w'I��@x�6�����H�rH�D]�^:�Ը~kLN�2�i/PK�Ǐ����ֱ��n��{�d��	ZtO�xSEf&X���c�����	?�2��ZiO?է�Y���8J�JT�F�O���"/�
*����6v#���v��ɸ���c;|�ت��Y��2΅�P|�xĳ�/��ܒ��b /俺	T� ��^�9^�'W��޸����jT~�Q	��y��C�в@|�+!M�s�!ͺ@QI�HǸE���x��m�Vӆ(J�">�p=b:�?e>(sa �o�?��agHƚX����4�e<��xtF�/��|��� uW�S�-7X�����S��R��5���Y���.3�˴T$�R��1��i�{
^@Z�j��0����� ��PG]���32,e�,�1+z�NLo־�N����Y�Z�W�>ו�\v }��9�Z�A�2`9��=�*yS�ͅΨ���?��c~�Ŧ��?W�Bp�j4á%G�e�]�����J���Y��Y:/�'c����x�\W{�,M�e��u;���r���3�/�n0%���3�"s �Eԯ<�`��S�E���1j���-��*o��5�iD��U&o��2	Al~�pQUc����Xq(?.��H]�1�(Vׄ��s������0e�q�v��T�|%�d�/F]05
�G�Y3?���3�wc&���J}��jR�r˥�lw��CEQ��,ڛVv)0%qE4^�B�J��!��>�5���.��&l�;� Q�F�f�?�]O�+�򝝚��:�=���fp�b隌�]m?h��Z�.>JU�q<�X����Ǒ�T��7��w��_c��z
g*�����J���|�H�B�	�2U��y���v���)�/�6
*=2���٥��-���iȖ.��N6\Z�ȸL5q�"��Y�K+��	q�O%�7	�"<��E$�F�*<��}�¥+v.	.�n�Fa�0��ۦ+����g�k&����oΜ��������߫4���UBސ�4Ÿx�q��5��8PY�CD!��W)��A�M;�a��G�lƐbN�� ��aa݋&�fɚ��f��k)��gʲ��-�夋����q����:˨�R���c�Ñ؃}s�:.�Pu3���N���0��z��gg�x�#��9á<M�
� �fMO��� 4!�Ҍ�Bh�;�5�,J=R5��d���!���T�CCM]����ԼI��/���r��ݱD�#˱�b�6�yl�L��_���
�:Շ4(̶�B�NLO�LL���+4Q�]X	���E�����5Y�֖"1�\b6T���P���{~D;�4���z�w
�%�)�4�U��8$?�,����BS��b�-K;q�c�2�wƊ=��aA~����WS%Od��"��g�þ����a���
L-'��=աҽ�8��*�7�w�T�qN��p1�R���V������������<ȓ�D[Q�Őc	���`�����QWBZ�(��������s�?���J��1�¶| WY��k�`�Q� J]�=�¤&���y��*'5-�%����I'�Ӆ��.I��B۾�B�*fx|��h���O�mm��-�$���A�U����3Tw�[�#��fA5d�M	�
�zT�|���?�X.Ž��i�"���4��$���}x���LK�y�Q�-aȄ1���K��'��*E�l*\�.�����/VX� H�)S�
ěs;UW���M4̵W�Qϥ�n�/Z0��节�Q���%I���:o}�'*�C)���?YAWک�ܑDv��D������a�
/�>oV�8�e���V��K�8ػ����*B�,$�S�~���a��q�Q��pR���n o��e@�_���Ɲ��f�i��� �
ww@���ל'7��z�M��+�6��D��3�9@�;4M!Ր^o5�E�/�Q!��5rk\i�fWm>�!We��\�'��h�3�O.��`Q�P�S�t��U-8,�����nR�CY�J�Y�/mP�V�{���;�����E���%���vzelW����<���~�K�?������iF��2Y<�iI���K�(�_;�5H%H��Z	���	c!�P[p��<�ŗLJ޵)~��sm�{(����f�6!�uܮ3ޙ+Ev��i&3��3Y� s ��������4� ��T��DG�Ђ��.�eO�{���hn�Z��O���6�� 9�w�C����#zA�;��xC�9�fy�����A"J�����������d����^,1'�+�Sq��K�ک���п
��Ϫ;h}��{&kZ��
4ƅ�a>N4_^Vͧ���������X��-�`[�����}�&�)���bI!�?�l�����0+.ݥ����tGI�2�S���t���x]�( �o:������X 4d�둩�-DIK�%zX:�y�{'����4.@�喸o�5��P�,$KX��F����m�|8�4�!�b�@E�=ǘ����d�yT�4W9�Җ��~�\�o0f�� �{W⮁��CR�c0��o�F��9 �ki���5�~i��ÊN�:�^m ��.���+S׈r�2<�)���9���m!e�=� ��o\ �}g���s�NsK�0%�x��3��G�Dt��!O��������~(�����o���t�
m��⺚;���]d��lf��\7ǮeqMr�ܚ��;�G�FI�L�*M?� 1�|�Y���Ax{g:���)��Qxz���6�_"ȃҖ��|�O@�h��w��ګ'V%�K���c����@Fy_~S�f�W��0LX0^UatH�N7��J��ܔ�r����`{Lh/e-9eN�'�=��k�rr3���ᲳG6�Jƿ��\�$�Lau�
29>0������Z���@k��׿G3H�BeǍ�$��ݣMO��_{�$�,l˷�G��h��$C$*�<M�χ����������:�w�Bi9c ��AI�$o��0e;���D4�e�c���q9'4�e���E�΢�I��;���K����?.aF���ӝC���i�$חd�G�c�������u/~s}�;�/K�����`�smAO���;����&���V
K�ki "ll�'Z5�*�W�p���%�<\3�5����
��g1VxaT3�2��3I��4�wW�x}�)����Q�D����� ZB6�L��@�/��f�_�J���GR]����;�L�!�Y��T� %V�D��x��o�.�����Fý��8�"�g��^�T3@c5�S=W��82:C�y
�K�����KT���ωÝhަ��)7*��{�Ջ�E��E���OX���
|�@�7`��oW�ՠ��:>h퇴�è̓��'Ϲ��~�172����';�}!날���������v�OG.�Ig��4���'�MO���E�G�ߋ����t/{C��V{<W�aN�͵��2�%ssШ}^��r�+D�U���5J��Dl��p��aD���>�N}?K�&Fyׂ�B)��!g�u��.G9ͽ����Jo�R��q�њ��Ɨ���,�����~6�D0�p`"���W��R�臥��5q�1���0�kBV N�O�3У^Wq+n���^@���a�ྶ��Q��\�ą�@\ߋ&�99*����!�Ds��4�8��3�/Iׅ�ɤ��i��_9�[�|��(�o���u���x'�[`�u<�H?TK4�*��-����==��%�|��v�\�t��9�M�^�Es�Թ9'��v3�jJ#�E��;�RJz�_5��X�|��������b����#n����Wvt�>����B�g�Z�Pt�<2u;b{�J�zT�K�0�Z9q���0�$����|��r�,?���f�`��y"u��/:N�T3�7�J���w?�H�_hP�O���]��P�WO�
�！?e|����L^�U�u�7�N�覵�5�r�*d��v\6����6��t�|� �p��h?9
 ��q��>���͚B�L��.�@:)��h����Z��+?-��壠`��� ͓����S:Rw��:���M�
,���,{q��k����B��}%e�P��r���@.�hm�a�*�Z�?̶��&���Hl�n"\�;=��i���%Q7��)�9 y�ܸ�}�F#�:[lA!�>��Bf�����8
�;�ƂN��+��e�����"�D!�hG��F��[�&�C���������AgW��K�S?_��!K��Ȗ��/� π�X�߮����S9P�>U��?�T�zy�mꬼ�G��M$Q��_|����h�7%�T�>��\���ÞcV��~�D��"GF̎{�h�jV��J�m��/I�˪)�> ʅ�N��&ݓ���H��C1�la3ri[��S������9����w]~�)�`�J9 F��p=ހ�ӏ�>;Cg�G9p6����-4β�J{�5,}��2�����_��f�w9W�8gY�d(u\���ZQf(JQP����$y�p���Oy>b���(� �Z%����|B���P�LO���c\��S�(�5���9�&\6֑��&���u�?0;Y�tM��Q�~Ӭ\,J����(�:#}���?��ũ��J���M��}���ݱ;dj�����������q��S'v�̺�a�y�ͮ�@�Tb�z�秢2�."N�1�9��#�F^��(5	m:7�ϙ��
��Ot'�)�}��j~9Z�l*�x�ۖ_�]}>��E�o��W!F��k�T+�»���hoa1��1��sy�E���P}�%�3>HrSr�������I&M�GǇL��פ֒c>G���C�"���Yx���=���aE�J%�u�0[����ʏ��<������@��!=	�`C?�*��8��ub�Hi�b�}uOi|j��a����~F���J]B�8!�=���YB._����Ph/q*Mp���I)�
��<������G�j�,^����2�����ć�T�3��a㕬�B�﫪�>�k��Eܕ�).
��.�糌�9_�a�V�B�P<v�_��<�9���3�����-Ж��g��R���h�|s�F�Z�����X)�
��X��'����V�7��C�_�r��U$�8Ih�:�E��0���?���ݔ�.�o?f�d�f?Җ+���;�Q|q��Ѕ�#P5G�RFQ^U!Xq,�ʚ�X��K`acG�z}*}��
�o���"���/�m�i����ϻ�,*K�[0Llc�b5kI
����c�À7P(t/9�k����qG��'z�VP��Wˋ!�K�9��J���\��e��Q���~���P��Uf��wp��g���txOb�����AⰘ�2֕IF��.�fe�(�|��2�sQ��U1��x��]F$��z����
���Kٟ�Z����(W#&%�d���LhY����RW����AҐ�9�p�<0��JR�_�i�w���mδ�ʠOo���4:=r�ّ��.u�5�����?hd�&��3�yM���<�tiϹ6^�>� �]�!��U���������~4UB
�m>s��e6a�&�ن�^��w�q��b��k�1�	�1 LA�OBb������ҵ�Xa�U�hM��|����ɀ�0��X�j'x�e�l��0є?+�а�������,�zG=S�Q��u0�I�m���6U��[�i;��EY����pe�̫(G�g?]ɁU�,+|�pM�;Ђ�N[���Y�b:���؆��|��b ��ǆ�b)E�@��j�f?�}�y��P�X莕Ʋ��0����� |����K$
� 	��v%��$ug�O-��,�qm�"�伃����o���?��$�|��{�ϋ���s�Zm�/}mj\������LmH l/�����N�+�+pQ���[���/L�S�+8���hY�y����;��v�-�m$�����k,qV?,z1�Rqo��-fd�\��#]�X;��;Z
=݋�����6w�	)ߞ�0�<�5�i�mD�U���&?�O�I��c�JMM�:��\�V?2���Z����<1����ʏBO�;m�}hs��PS�����@�b�,�wVe�Ɂ`����v}��UY��%�sJ:�q��SK@�2��/3W!yK�T#+Clo���x��Q3����5������j~1睥���g5b�Ne͠e�xU�F񚱙&)~�Ԅ��z>eԻ8��q,���k�dm%�u��x-��&d�0ς)��H��Y��yO/���-�d7PK���a�J��C�w����p?6���g�~�^�89iRz�|&*]sD;˶y�S�9NhA���V��4N�	�NQ�(�R/��]�M���	�ȷ��j\~s�,3	�]l�E��3C㧡?4������u��ʯМ@���T�
6���a�D����ZAh�����OⲿSIJ���6'BV��mQ���+����x軱�Z"�Q����	����-�cp���iz0Sn�G���#v2Y�!~���(U�Ze�'�R�ߪB����Mx�m�夓�_`ᩫ=c�x�&�E?�,<�jӠ���pZ>�~w��S��Dy' $��>Ѝ'��za� ��((r)�P׶Ĉ�]�Y�����f]�4z��@?*hZb��;`oC�w)���zj�l[��=��1w).p�3��b��-�Ԣ����2z�w�*fwB|�Eg�6�Եl���(�sM�L�w�+}�~��>��h��גa_���?S��.����R���⍄��H��|r�G�"HG���^i�]�f����w|�vw���%�@pj���Yzy/U7��\��߮ȉ�#�sc�P]鐡�|��E9����My��dml���Ɂ]�k�E�X��(]�L���t��rA�>���6S+�	�nUNy�1w6dS�p�p܋�̮�K둂5��nRG��#�J���\��kC�
e%ٰ�+�B��՛������>��X��'��y�7ڼ�'�L}`J7 �%�x�P��Ɉ�Mo	?2pt6�Rn�W*8 FBO�
�Gm��=7{�VW�}z,�{�r O�h.cf���%�)���ur~2N#V3�w���'�i�e���uXBF���aسjc�����ݗ��"�W�GC�s�n��Z�u:h
3}�@�h|c�a&.��$����x �Hp�f��J�=��C��\���W�[��;�q�t�,��߶F;-J�x'ꘅ�~����(�S�dp�?�[�O-%���l���o�29�6�*!����KR�g7���'�(ޙ��,�����c<���h��*�P��Ӈ;U�a�!^���|IP��z	5��������a�+y-����[;��+�A��;�}�¿��D㫚���PpL�{CN��o&�Ww�,�0ae��;OUd~���n�y��/�䇙&l�|)a�A�[|wOq��0�~TD�^�@�I7#��j�-}D'�f�ǅ�WNoeE�N� �`�����&�,�N��(�A��q�2Ώ 9�Ђ4̡�fx��G�,�X��p��������)������(�O,������+�=�Z�@��Y+|�N���R����p�-�l4j����,z������G�c'�8����QW;�(���aS�?��]t�$Pl��ǎ�O�]i7���V&G�U���qA��)V~p�T��B8�Fكh�5�I#��+&7b`�;���bd��0�&г�e$�U��<D8&�gi_�*�;䎚y0��L~��|�S�03�7�W{<�~��Ė���V��l�Q !C-��a<.�7�,y7�`(�	�P�i7�F���B`6UJJ�s���Q�G�f��?��Q[r��F�g�\�|�����TJ7�7�?�K~M�;7��Ԣ#����I��Ʈ�D��Z�іnc;DH��1��*�r:�]�����#�{U萗i�M�{/��Z��1<�)]�UDpD�Bc:��"��q�N%d��}��=[�9��`��וDZI���G���f(O�D�ɀ�z�R+�M�:���D��p��Mo�W��ϑ�;��60�C����E�p�[�Ȗc.b�ݔx���!�jE�����nБ������hZ�^�(3Aa1"<��l��"1v�Zэ�g:��]_Y���I��@��#�<�3�e.~sȔ�4��-gq��o�H�슁�����硧|ɿ���%#�ɂ�w����s����	c5ß����=�I�7cL��ݙ��I���I|%�x���5�&ǡv�[�y궞�o���!TI_>I���eg��j9�L��X�c��elj�L%�^�c�����D	>T�&6�c��{M4i���h���C�c�{<OՔD���KN�u�f��vh��'CP7~�fS��u�w��6ю�9 ����_�{MdNq����DcDF�p��A	������Z�A, ���.�bE�8�����_: ��gݣ�0D�$��6���Xn"<������4���J��N{�|�s����ɴA����[�,�d�TrA��JfO0�v"�C�1�V�Y�(c_y��# ����5є'|�]�M��8�5t>hy�!Y��hC˥��Q�Z�l��Q]A��u1�0�v��t�A��`7���K�����I�y��H@�\&���V6pO��z8�2��(�n�?o�U	��p�]� �u߷e:�:�^�拵L6�B���M�Y��y�M\�!A)z�qF�{Q����V�L�cQ��~��.��;4b1[��_��-���[p�����B��@���QlҰ.�g�.Ҫ�ay֑��1#3���a�\�Z :U���2�n�3�8|�6����|�OĘ%�o�F�|pꯪ�8T�Q%���Я� ��h�������-
񒁦Tt��$T��~8��A�!�r��Q�3��Gd[�����P�Å�|A��ue^���|�=�ӰÔ/`)�ΞX�6 :��R�8�p9���y��1ܐ��8��R��hV/�a:XY�%��-؇͛��&:r��lb[��)�cT��9)��H����7�2}�mJ,m��������f
�2��d`�͚ ��?*N[nU@��۫�er��CRt!b0F��e��Z\�{�f{��+��ѩ��ϖVp���z�����q�o�?<Ϝ�����1Df��I��}�v�a��������J��
Z=%�,=���4Q��!���J$�y����R�)�=,	�!I�U{��$���1���ֱ6�X]/��L�Ie��w�X���Jc�m�o�i?
+�����D^�F��`YΣ�k���\�Խp�����_��(���}�c}]�����/�r��9()[�{,ul�:���o;��	�q�$|����r֯%Ny`��t-��m��`{g,U�&Cx�2$2r�i>]s������r�&�G��y�񅴹~��;C���$]�)1g-S_����W(0t�gL[�y�H����t	$�X��;a�t�&Ç3�-��3��c��2�k���v;`D+a���8����0�ʇ��J u]㗮�Q�C�s�T�t}>�H���5G��h��������e��J����%�Г�����������}C�6�v0_��F�c0B.':�H3�|�=kղ�49zt �tfV3*�4�2m%��" S��iU\ms�����Fv#��xF-�pi�+S$�'=�W�`JV�*���=��i<�'J���ވT6�/OA����YHz�5�r%m	���#��.X�cϣ�/��O��.t�-Cv��R6�Ѣ�&����<B���rl:%U]�����r���I7T6�yç)F��Vzʂ�� -�]M���A�ʈ�q�#������PY$���7�B0�bm��j���1@���6X3��~��� ؀�ya@�;7 ]/����?�ֵd4�鳗�&%�:�gśB��/&��辝��)R����G��7"�J s�� d`,?�,��;<M7�
V5��C��"&�pR���H�g�&�!E�(ǽJ�{��,���%Mf���*[��tf�~��LyM
Z���`ӿt�Y�gv���%'N�e��om�bV(��[*�@8'�w�WN�������{Y/�"��y�w�.Pv�BTF9����k���%ݮz��������ID��\W���:��	\�O]��6G����k5`2��İQQ��/c��^��L:q`}�_,;".7>h�AhC��4�i�7��� ���;��]���]�[ry|���ݷЮ�\Q���:�3���m�а� ���FC%���@��l����p�Ŗ���T��I���'B4����!tsI��������J�(��'gf�[�������`�בap��(�3Z�-�o�l�稽��W��6*�@ĎO�~s�CY-���[�������M"@�p��d�ⷔ���ш�`5����Ρ`:� �Hos�4�aV"쳴T~��n�ZSY�H���줪�k�����NEEf�
���@�5��ԟ��T%�v�-����>�i��Q�>�hW�ڭӨ�}�x[�I�K(V�1i�D�Òs�B��䒄z��A޵ ���Sq+��A����4LLH��Su�dc�7�s�����(�-S���g�-��frv�w���0W�h�<j9`Jb���-0��a�(Kr������vbi��[oy�A7b|C2Ȋ��S�KG�7�6��y<O�<�%�y|�=g�(U�����O_�\�_�,�Ƌ�o(�6�Xe�T��_�tG�3 p�p�ILu����To���-���lFjpD�M���9�0�|Z	�XH����Vov�i��S!���,=l$<Xk��i��+����CZ걔�q�̓�f,��9�4~��M�C�P�4ƀ7��1�Y��F鳜U돽m|��6��]ޘ�I�Ck���Tz�%]gdE̢�1�?��Q���ʛ史���Xa�sʰU���%��A�st�ڵc��ܗ�[q�h&(��H��ýQ��\�P�e����������H�>�M�a���]��X)\��@*$8r�<�,ƶxJgSP�y�1wH��!�(�ҵxP�o9��K�@\��Rf����44�!\B��uC��i�/��6��wh��Cd�L�P�q����|��v���p�Y���pG��^�y�d�~ �+�)uqd���v�l�7?zPZ�3
�l΋1��\jӽ���,�=�\�)����2�{��OY�d�"XÌ~�����~������A��[%�z+�uCaE&י�Ao���̾(T=���$��w����΁��b���|��)�me�[�Hq6�C���
_�~�O�_ݬ\2pF�x2-;'Փo���_�O+�8!)�����w���[��4(�f4�*4�c\F�j���bO߾Wk\���r�ߘ8_������7�W?��~��3%�)�������&<���%'\�egK7�U1�ʲ���$f�R3�w3;���闱��b�JXdHk��y��z�ץ��0����@og�I2n�n��4mjAOyR9�MH3DۗP~B�!�,��W7r
������	D�G�ޑU�l�C��5˃<Q��4J�;������N�mWQ����856�?���	����NE���*��62��}�]�H�sw��u-wK�H���Sn���B�3�6�/�r�����"^�9#t���A��"AԌ������т�E�Rx��1��p?F8�dE�Z�����/&$/)��������v���J���a�|w8��<�~����լzU��bb��5�,K��{�x�Y����3����Px�y�A�yg�y�mz��(h�g���~Y����WZ�+���R�C���{Ċ��K	Z���i�8GZ1�Wc�-��e�I���1r?�����/�y��}D��j��xX������=x7���� ��O<>�?j�y\�.��&? ��l������{s�����	��Es4r�H�3�y��E�d<ѝ�J�����r+?Z�P2�!&mG[�<��ɔ�e��"������UϽ<��<��;^�Z��2[��w�a���P�;$h����_��C�*�)���;��M}O���'*v��Џ��
7�<��ipP���!�o�áPKֺ1�zmyļ)un-q���͋�υY��C[&/Y��FA򋭜n�����bg����
௸u#�ܞ�qW��I�ϦA%�q��C�D�v�M�����x�1�A��Hnc��Uh2,�eD
^��p�0��c�'^�C�u������D��Ix.��d�a�P�E���KI#�����<&��~'�?�Wv�=.������xk���µJo�Œ{H�C�&{�����xQt��en�+�w}�$*����W$�}"�c�5�K��z�+I�uM]�)R�i�̕�*�v���%���w�l��S��'�{�Jo�a�_�~.]���+1z�K,z�4$WM�e�k�o��G��S�Y9�}�M�[��~{�6-�B�kA�I�?"*�8����&㎟8�>�*ˑ��k�`�;�G��
A���Jh�����Lz�T�]�Ec�u?{�O���2l��� ��}*5=V�� ��Ћ�(.E�+*p��`�f	�x�,�/,ؙx9#��jR�9p��yA��U-�9��{ӝ�m��lOkƎ�����	׆n#V��PP�X7��Ħp���xjB�>R��!h/�e��/�xe��d�d�z7?��mӽ��A�L�ѭ�����ZNu�+������x2�ӏ�� =̩���_~ً�,���f��>�5�X'"Ve���D��,+�	*nA/�73�@މ	g��aa�m�Q��5�5�U�(>	!�\J��g�P���n��)�L���>�mNd� ��3l,_)�ͅ�Z����H�=8�#���&�IT��CM*�F���X4���>�e9������A�(���e���4�i���#�>�ۀ���ǰwP��g����a��Zoe�W��E��7�Uz*��iR�"(�F!��}V�,����.��W��5�E{��`uu�����h��|��KO�HN��_X̟�S0�{-����[|���_,yx*7ϗ�����#���Z��;��������X�X�������+��G ?��B�H�{5���@��qÆ)��K9�u�l�q�����׍��	nj��]	)9Ѡ3 �b��_G���b����Rg9b��E��,�߶�0K'�e�0��=LR�p�a+��\~�nG?�"F��+�|^���@>�v�	,\N򳾥
x�����X$w,:ՒYs�)ɉ�%����k��-�[$�� [��\�e
��.��].��z���? �ӥ����Ռ���x���+��K;K��YYd-0�[���:q�����u+�1�+��@�����X��Gzp8�jㅐ�J $�Օg*�?
+�wF�
���X۫�<��3;�$�*�W@a&� Obj'щ�O̪�Lv���)�0����4C�M�[�	���X��*�H������Z_ȉ��m��ͨ<��US�֓+��o&��x�k��V �M�%9i�8Ρ��O�}�RI�Z��,`}�*@����
g\��i\V�ZU#'b��F,VmB�aw�-/�	&�+xz`�7�@e:�>L�ńJ�?������lM�FL���d�A�� ��-������\B|�i\���پ�\��7ȗ����������}�.�_5gP�5G��-}P���/���,2 	5=ݫ��zI��
L�x�0����ڡ��_pjPv�# I�����(2�MjVE׳�z�zE�Brcg����L��%��Q���$��?�p3�,�j�ᆠ���ܣ����ݔ&��{�f��f��Bd$p��]q*�>�/�-'�.��F���q-f	�"]`����E�ɀq>��6�ʺL��IE����>�Ǜ��?��<�nvAC(l�hO:��sV;#y����?Ȋf�JR�z�{|���=v�#Vt�j�<`Bn��W��բL�_c�(V���[�> ��)d+���5��j�^�6�ֳ2_ͽR^,Bb���s�@�pR����,�ڰ}���]엄v�2?��~}�Ϛ�m#�"a�b-Fm�{R��V�g��o|��~̆����(G���+�f,Q��˻g��:UQ7K!?��Pt
���ՈyL�E�j�w���^�jLae���&Mۊ��R�
�WZG������X�����=rP!G9�cѹ ���ӄNL64�ZMu��G��[Y��2�J�	�� ����wi0�ED��q+�>�X4�޶���J92��z؝j�v�p�����n�l���'�8v�Ƴ��k}]w�0\��u��gj�FL�^!�)1��H'�xCW����ZE2���ƍ���*�'�>F$[��ZW^��q/u���Ɓ,����S�ȶ�hq�m�:`�ԩF�[vRHrs�(�#�W��PD^�}�LV���֔�N`��L�0��M��Yy6�.��^�c~6>t &I�T#��&D��3��iҫ@HŌEc8^o�I���N1Ն7)?~9���.��ܖ��jy�u�N�G��A�`qW����0\8�����w%<�&dʂurIc���I"�����>�k#	i���t*}�x�K�.�Vw�PEXt�Ӭy�����-;���C�)PZz&����_�N�c���?����E�32s�*N�CxsȰ�sL�F�&��uz��l�Q�	�bغ��^52��2�G�EMA�(hkN>��5^��o�͞�= 冔�h�UF����r��ɴL����wQe��BT���5-�'�G��Ar���=�ˋ# S�(�_vY<�������-�^�b�{X�0%��Hl�*2Kx 6����@�Ń��Y��X�lwR��O�\�{��c�p'����%������|�>��O����'��2�^Wp�#\��՚ɲ�B�;���!TP�����R�Ƣ���)w�΅cA��3-�<�i�~s���v��4F�t_��
��ϒ�����o�����s��*,��}�_�@��e�ZMYc���b��C��3J�j���Pw:3���Ԝ���`ԷG�:�����+���v�Gߔ��hp������")=�8��l� �Lr"ˀ��J�%]��PG� �4� 4����D�����\�	�T�C�-�|!b��Y��"����pB������F��>�7���dQŴ�����M0Ÿ|�e;�@�:����*������;�,��_�vP�4���pk<GpV��$�������"�]�P��Ț�ww�?h��V�u�IPߙ���$��D��D�4�����	%��|�!�"�o����)�xB�xG�:a&�'���l3��m
[������,�0A
B b�.���nm>^e0v�5�k
4�L?_u�6������=�vl*Q{!7>�������cD:�,M�PT�����&/R��y�=�O���Ҩ����7T�*7b���nąX�z����I��~s��%�h��[��ۑ+�J~ȐHS��7g�G|�~��y���a�; ]?��P��:|mu������e��^/D�+��=@�2լ���=�A���Y��~���{����h�[C���#�eh ��X��L��p6JZ^�X2�olH��bt�j��؊$��u���^�O8���;�a��q��IB��n,h���X�2�+� ~�MyA��f{�����LýYH�G"`f8g8N�S��=׻̊��7��=���9Z�7����X��0e��R�K�a��imY�,XX����KK�<�x[��0�`Y��?y����3��ҫG��~-�G?�Sjn\uښ䝲�oW2��Q5G椴/_���u�,��g���!QZ��A���B;�/����N��y��=�Axa#�_��I;�w�;5�z_#:^�f�<�%�;c����9lz�Č��/�\+�8~Y��U<�&���a)�������������#�tF�I��]C������tw�^�82^�!�B\l����ʛQ��2H��"kÞ	���0g/�(=�D1@��Y��iM�F(��Wr����2�m!��d}k]%���/�,��Y$��T<���U����3� m�at����Y�U߳r�~!]6 �8MuM_��I8z����&�S�Cم�%�S?��o/��{!�i���F$�PrT(p��>��̇v$�E�����{�A93Y�:0&c�`���>,2qLz?���.G��t��>�/yp�9��I>�1����BC!������#��*3pD���!�_/��D���6�߬�)��5a,@�f%��vj=�:�vQB���d� ВD�EE��~�KGa����[���F2��m�0���/��n���|q��#%J���خ����8������|3,1�"*�8&�W3]Q��(	Yx����s�M����H�5�jI������=_0�<����1xT���yL���cŚ�"x,����6w
�淴ƙ�j�nB#m�)�IG�
<-%�)�򹠃omF����B�i��t�!��ُ���Í@1������Q�^᧐�gT�s	o�`9$\ Y�Ȩ��e6� ����D%��:�#�Xc��s�%�T=��6�KS`]���du�<��4��~��9�<vf&�(�)�\xڡ�3�,��|d1���x�����D�2mZ�y��#:���\�Zv�?E^Ôp�3f>¢���=�83����p�7��
{T'Qm0�\P^`_7Ln3{���W���c�+.��1��0�	��}�oOl�F�1��'�����3�mB/ ĨK������9���� ,��>�Y�i�)d�����c8�����^Ɏ��^� ���59p���+2;i���B��نV�o�9��хi�i��AK�/避�4X2îʯ�S���`2��TA!�O�6��a�Bq�kֳc�Tp��~��'NR-V4s����2�_�+��YW���
�hj��XQ��$Z�z��fl�ns�Z�=��'0.Ber9,��-}� \����M\�q9R��Y9�R;���D��]ǡy�d�ٱ>^Lf��O���.��u������5@3]�L��n$&"۽����o��s���"�ݬ���R�[Z�+�m����t��[l).���W�w�H>j��DS��� F���]���`��~�S��L5�^@���Ha�t/��O�~�q
v�(�k�vL��񅧘�l��q���A�·��1�;2O~Fo�#)���&]w�X �$�^-�Y$<o��Y6�p������$��2�Qme�ǈ�&+��AX�HIH�fݤ�ի��͍^"|?AO�׉�r�y׺�p��<��:U ��`�k�}('�F��K������pY���/�k'? 
�u�y'@0Y-+߷���D���Z�H�el<a>���jߖ�Z=����Sisa�x�.�Az��eT�nem���m���;�-X񊏷	�I;�H��<G�x�k�v�g�{XBYkav�ƶE󣱁�
�y5��]pS�R��X�V�F���oW�huy�;�B:��v���j�c:|$��C'z`��.%�*4�5��őd����p�Z~�6��_���A-F ���l8=2�$��|i(��e�҅�M�{����`����/l>��e�r�{�BJٸ��Q�D�Ҳ��������,]�@+0�iD�����뱉�D�����^K(j�،ꐣ��5�h��_&�at�3����u������fh�/�5%y��y��	*%N��h]y�0P�%�H�����.�p=��!sK'������S��it�L��iRsb({�U��.��:�����I/Z�r0����7�� �-����7#*/�f�p"��\ڌ�]S���̕S�3�ң����0��+���$a��BAF��~�Wy������W�&a���v�^��]���U^~���w4�f��>�h}i�9f��*{�\�z�05=Ⲉl�£��z�-Rn��ZD�DNօԏ�]y�P�����ښ��VԬ-N�����c�+:P#����!��F��\{V���<���b@�C݉���A��sվ��};1.����b����N� �^z7���S�3F�`�L��t�FXS1�E
�4��\1`^$��S�j�D���c���L�q���v ��[޲A{�..��w�n1F���~�����<���[��c>X@�+�۬��夽�u�Xy%�gX����X�P�� 3��\�W�+�����1c���c*oCF1��er�=����S�e��v��q�*�~�4
t3��4��î1��t�)�άr3EZ5d�λ:�ʗ"�^V(���(ݺ6q
��J=icWPY5u��F�|Z��q8�aT�l���	��$s�JZ+�����5K��	-��1��
�"��Y8��"��`O��Ɨ�|�\/��O]�f�i@s�fc�f
$�!E���L�	�I�<!�ü�i�3T��%���q�O�Vt\Bn>�9x����y�� ���/�~U�^���^����lD'����:.ɮ)�ey�il>�:N?r20	�Ĕ5���A
������^c��J�&X>aގz<2$�ofa^��P��:����gw|du<U, �]Q8�~S��ᱫ���ީ%���1:�wR%�z�	Jo��H*l�|��
v��LeIO�#5���o�U59�z��h�8au�P�WK���u��_��
<'h�=�,�4hw����{�h{�Sv��3�Z�;�<:����$"Ĕ%�R�ήeי����U
�>�I!FSʪk��d\ذ�^��f��i\4���8*8At1)[u�n�!�E�n>"@$}�FˁU�w����FH���euA�]�&�MԢ<8�s�i�^���;�P�e�0ax�M{�r��i��r�B,xS
�����_k6�_��Ｆ��fx�+48���_�	A�͢�b��D��6�����ΏR%rT'������Y5��G�=u���k�sS��:����y+�wé6m���;�Vd�d����W."-� p"J%Cj�䅿^��:���� p���;�~�B��zP��~��[��d݂��.�
p�W¢E���d��!���UT>Z���Kh�8�=m��V����,3�6��	�]��q�~ ���]�پ�ȥ�% y�3�"܌7���O�u4%A}D��B4Q1-��֐�ۼ��=eSSmpAM���a��M�Fpk2i����pK��h�V�C�畧�&��k�nV4��H��u��Ll���hs`����(?��_c�&\��n�ٔH�՚����-J`��[$!h�܁��,[��|/���̜0dLz�r���/�zͭ ��90J,~��q��-O)�!t�V�n�� ������85�� ����v��O��Ut�v;q�������Vc-��q�\�K�����f�m=���U��t�4�/�Dp	�a#>H���q6ձ���<Q/�E��'�	��͚��4�mo������qR�3�5�;c1�g��[��L��SqJkԻƀ�	ҋ,r��Fd�ď�����?��8�v�W�Kr1s6F�(��M���XZ�-`�	h���O� 8�pI���1���(�oK��§Y2X�����m�t� C��>Un���*\&{k���=�P��7�����t:t��Y�3�1z��`SaȈ%�b�ڴ����B%J{�:p�;10����D���p#�Vs�%x��4 f�I���	�!���ˠЅ�/���f��A
,�R�H&�TLh�"igݼ5��x꫑U��2������?��sGkO�/_�E_��^�Z'�`Ѻ�^��K͎�����m�%��w:���k)CM[�k�[C0��E��pB�H��7�PQR���K78����mLNT|1��Mpt��)���6h��N+�vW���ZyV�E	$�%�mp�%��uQ|zT"Z�>����Ec��a~�+�=ё��L��S�0���͒�R������p�q����Jf&�mcN��n�X?���G�{�����,Mm�1_��`:�س�a�Mh_���A`��`�����7)�H�� Y�$�@��q��5*��*���f�3���_�>�V;�TN��;��F*G6��	��dkL]��0��O읜�=R��Yi=�[3K͎:BԽ�|{UJ�mqy��Ї65,_Do��Lg���cn�6l�IE��S4�w���V�.��2��fi7_�:�\G2l;��:���bi�ّ��C��@CN��nx��&Ս�.�xa`��sX�7B�@���fT�0MV��?��a���LN�= �z�w3��+�5 ���8b�.�H.z�l ��N=�Ķ'%#C٬d�c�\1�;�|n���=T��>�QObp�'u|_�I+�x����wĆ���Ο�n���$�R�A9��peR&������Z�a��%;���(3��w���*�15���Yi�S>.6��g=+|�a�5/���Zl�Qd����n��<���y�lE�:���0۹�*ø��{/;ῡ���� E�v�s^�������ZJ�9�e�U)݁��2o�!��%��&~� L*�ȶ�� �OK~����Ya�q�T�!��/}���z���,]���{�0�y1��	5�M<�Mk���b��3'��6׾ײ��������]�b�ڥr�	�����_gn�4���$S�D�+��h~Sb-v��H���
�I�i�&�VC�����ĺ9K�	�f%Y�kʎ�*��Wd��,p3�Ҝ~d2��6�41�~��g�k�/�	���� ��j6�A%�L[\�$C="{�ߨF��O��$�5�|����K=��K�;(Q���uw"U@�؎��q9G��NJ�g�Yȷ	�}�;՘7�����H��Т���j	�Z;'8e��f����0E�I�3�6��(���-QD�K +!�
��g�ciO��~i�}�}�i��64s�B&���q=��Z� ��MTc��3^��l�i����)�+�۠]��f!7��1�7�u��4���w*��\�@n��)u���`Q!�n(ur\raK��i�:�'���@�7�Vt|QO��z��3��t�
�'����P��JԮ9�"���ΠHn"�?��9�>���^��=#���
Mp�L�z�3����կ�F��e;�������`c=�Μ-��M[zB	�rك��j��L����&LѳbY;�r�N��~m.$�@�؅�AB�[�Y�xo�KK'�}R'Ko4.���6WZc|�W�c�J�ݔ�P�*�ViSP�H�|7s���g2���"S�����+0Ƿ��+�mĥ&�3��F�l�L
��qk�
�ETQ�1׻n���G���|��R�#.��kw$�]��xo,?u��X��p���,��3���+��,"0��n&�;��\���"R�4�{AM���K
@���w���`$M����;�k*3�f蚙�f�1}��4M�k_8�} .��_W.>!���f�-�J���us���h��D�ik6M��w�D�z��(p��� ��!U\��n)9u�d���5=��~ �u�z��I��tR� v(�S�!�����cҶ� ��/P�`��>��d.cn,HJ	����9-��9=�J�������"�"�:�m�����;��?�4>5y:a�<h�u�?���i��M�O]YYջ�����]'��a>��iɝ@o�������@��"6�3�#�F�����_�� YT]�`/'+wο��uk]��x���
��U
z ~���D��ڻ��}z��9TsC����_��(� K��n��\z�O��U��!=ڬ�eHL���D���/ͧ��5��I�g�-u��c0�@��`�C�7��}�Dł�Ss��0!�<�C�#��O~a�pD�� �|ٱ��6L�in��E���B���d�ƪ�q�o�
���Ҳ�Q���u�C��Qq +l�H�7�7�7A���s P�x��		�}���@v�0mN[��=�9�o�E�,��L�ж�_��_D�����פ�1xZ�^�<k>��E�x8QU@Pbd^�4?���Β�j���3�I�9�������k���F^u>�{�j��2�1=��[Q��~}6e.�0�l���xD�ɀ��8+��,ⱺ�<��?�k��#��Ow���Ϻ#��[��PcL)����q�$ ǃG/���x�����A��>�jc��!1�oT��[M�Nl0r�N����'��g�+hJqڳ��u@�[/	��N�q�cP�kp�͟���0���߃�ut�e��	���T��"oy3���4%P���x�g�������g��1s?�u��`��C�>���H��C���"�d��|6��@��pt���*�EmD���3���L��n�����Q���C(>;oj�^��'�!|qv.L�?�x[{1�3јAb���]�p��5�I.��[Y����(�S�ȼ~�AH���TCT_�`��sU����<:�ߌH-2�מ�\�/�2�^�'�wg:��l��y�&����C�&���+�hqxGk���޻լAMrY~��f5��8OɌT$��!$3��L�q�D�����Nq$�+܍f?O7C2e�D��"Ɯ0��
��Js0���Ӕ� ;���L.R騊�5Y�e"H���pvr+��^���В�H��,���?��	����!������@)�����k`��F���W#	�EX[4�T��8�x�eF�$�jd@�v	7'P�ߑx��2uYY\	��TG�34�{x��这ytZMG(��h9l%"�40��� ����w ��y{N	By��������֚������C����M��B ���^q�Nl�AŒ0wF{7z���Ut�K�%nK�r0\<DFb�e�Y��/�3����X+�Qj�L�������s�s݃HN�"��&e7,>��x #XT�%)�z��E���k���9��h	1
Xf���f��c˃&F柌�ߠg������k&9F� U+��נ�Q,x<�&�<�P���Y??M����5�M��f��MH/T�gJ��z�a4b���{C���S�rB*����9?zQp��
�*=T��� ���l+9r:��ɼ`�^�c2D�M�t99�Z���)r�@�������6B����	 m�To+&�W�	�ňX�̨/��<�ҳO��R*3�2�2(ߵ��!W+)Y��_. �%-�}�l!�Z�;k"/�hKi$��&�0=��wb���}�D(��^`o������jծ���XNE�e�k8.=�b���,S��m����ݯ&�_�q�{�ҁ��l���8�\���,�Z[�`�(�R�ر~��c:��9��@��?ݢ�i��q�:�B�*�lp4�
��� '�7'�1�`'<�v�h7N�:`|���3���/��=��݃���~$��J�ޣ�U�lKcb��vzf����D0
�v��HU�ϙ�Í@l)LT&Ml��~{1�ӛo�{Y�FUf�h�MB��].�z�c�UՅ�Hl�>?V8�D��&�0鼕6�g�H��r�ξ%���?u�-�h��۴Ț}�bw�-{R!��vV[�`!V�fW���M]/��V�" #0��~d%�#;刕�k��i��Tu	{���|8�|H��-�n7�q.XMU�υ� ���-&p���������� ��~�����LH�=��	{$����-]K2��%��Z�%Iª�݌:ſ]0��E���rw�7�!�W�_:��Z�����C��)A c��L����=.�����]�]��5u�Wd��� qvO�Jna�g6R��D� �lsb��q��Q�/�B`�O�-�����T:���	7���:�鶰hЃ� ^�a'��]�>F�+��5��H �~>˟b3꜡��v�'��#��6m/�-uL{����	�IX�d�c�	W��+�����N^P~_�PY�b4��3��]����$��3�%���6ff�۲}��l^6�z�˙V&�u��mxؒ`i�����K<]ㆀ7j�M�Z�l�@�� K0���j�����7kV��`,�$�����e�������־i�N]ƛ�����N��`>I*�e���#�W[�=����E��wJ�Rq�ȁ�ےH@�K��tf�F�Q1H�����6������`=�(��E���0��.V�u��:��Fj�*)*��r�����\o��[$kA���3�悠ҵx!(��?;5�
WR���j���±O����������R�>5|�l9�� E�=h+(������`L�p�|��w0�sT�S�8�� U��5�+̊�B�ZFV��\̊\���P
!j����ٓ��=��	����pGs�n�gp9�t|a {>��H�$c7�yV�	ZC35�����!!�!#�9[?����9���R(H��g���j�Be�*�I�d`@$ĿO���t�
'��C�P�=X�P��T#��7�T�� ���<'�IB�L�Ar�a���4� �|�\�Z�x�P�7�_wa��兽��X�8?��5�p��'�H�j�����$��R���!T���q?&�Y�� ��lr�zQ�п��qΠ�����o.O�Q��o� �-���ePy��1)���z�RǸ�~�n���	E�)�����?�Z7��b�
Za��*�#�Z���\h����-�|��/S�i��!����M��x��|?V���ݧ~]_� �R��уv��֙A'�2��-ԍ���=�@��GM���^y��|�͛�������W���D�UޠS�+��E��dӌ[�q�!H�����=�����-Q|/��Q���u�P_��է�O����5u��A����YJ
��4`>̋V~�T��te"IWE�:�"oCو��U˿G߹<��K��t'�z�-lQt3��=v,&����)������gZ�P$T��f��:��e�z�JXU�)�d4RN��hD�w��hgWc��ƹ�zw]|Ӧk�5V�U;[�j�(|O�{��g����m4I��,��-?��w��p�tу�\��= <�R�,��uG�m$�b�lz�*r�ج^�cT�Zl4�Nu��LB�Z��u��o� �f$U&8e�o5��9���,:i$f�:<�Ф-� }C`hw������N=�;̦��&���E��/Ѱ��V<�]ɚ��ż�H�4��78Z�"*��0hª�Qho���������d�7u��+"���U|Q��o�J[��-
��|(`�f5���{����R}h7�Z�t�	��I2A�gqt��%m��sݑ�9G�95n�@f��~�S�w�������I▃�Dytt���a�� ���Ťk���s���*3���ӟ�VCh�}��tJ��>��*���6ԵǼ�\������ ���f ��_3X�ڱ����E��HzJu�t]����\��[.��U�:<� (UGqb��ה|��x�~���Az�Gr%�����AO������4���x�L�kJb�����v����U~��e3�<�G�~��r�{��I	G{��H���Ekx�2�:Ѽ�9�P�MA6'�eM^��di�x�����F,�ګ��3��r4)�\�j���$> xrH�Y��\����ɭ[E|L�pbi�s��鍳�|�Z����v�H�9�'6_��[�>��3�;|_�Zk��1�\ ˇTA=L�'�(iց=Z�;�@�[��0��������x�#�ka/��=�8�Kmz7nJ��xOyߎ&�5߆Ԭ�A�Ƅ-8�=~ςIq���z��	�c���5�Z�ג/c48�aI,��a�%�<YEx2��)�ݰ��r��®�з�� ���<��Q��`�6�@�;�|��@&O����k�y�x�n�
u0u��U�ݝն�ڤLݏ�;�V1��2?�9e�9Z�^�ׁ仛dV[�!�9�n�1��w�͡�u��c�('S/N�/q�7pg�t��ߣ� ����/�E�n�� �M�tm�rr^���B,�Q���b���'��\N��3?[q�V�Z<�a�*Z�=�ƅ�[D!��]m��}5�̉�km̯�=���*�}����U�:��V����6E�9���̄���oA�)f��2c|~��YW��!�ީ�v<R�s(k�Z���oS1����!^�Xgy��[1(��L��읳����p�(��������C.a}%Uc��qU��H�POф��9/L��<�J!a�]��X��Mw)|���Rc�[�B~�"�4�2cu;N$�� S��`T�4ݲZ�e�� P����<���m�c��rY�v��.���N����ߐ���w��an!˝�/��� o��eqz����ŊD��˩#����,�5y���JR��#Cm���h��겡Rm8�9�z3;����/�)&���I��@���~����t����:Qo���Ɉ�TQ�j��	߇;|2�O�Ќz�S����{����.���̭��?7�t<���􀅗(�� ����Ѽ�E����B)m�A̕�h!��85,ϻ蔲Q�����k�i4�$=��v�D��>��FS�����.�O�h�ʽ^��&&�ƍ��T�\n:?N���	�\��5�����p�Pd�i�����}�ᬦ"��g����F���K�TX�Ϛ��{�bBsb�F!�H���r����_"���tL�F#dq����,À�+c�� s�@<��(9��J�N�ЫO<��2���V��� z�Ǆ7+48�o�X@9$�3��\��HGvq=�?���EN����K9�`��.�w0�G� 4�^����}�\��R�A7��"�
A�T��!|��8h�:�Z���X�i'R�U[���a�&�P��+���Ֆ�/3Z`�~�J?��b>������W�Z�7��D����n>�hE�Qi.�*F�5��M+s���2ʉq�>8�+�T�����jVZC27�T.o��H���b�=>�e��S���1�w��ښ#�,��y����u����m����P�,���QP�в��i��#�h��̨�eiOx�����u$eA�z8�lT;b�3ё$o���Z�.����k�a�F��QS�SW&E���W�r�9��ϻh�|��m����9�Ks�	D�(�oK|��-��4|�{�ǈ��8��AJ�ǲ7���A�|���Ɵe|zٝx�V��<i4��Jp�I�����:b�q+ʗ�NK���y��q��p*�2�ra}Z&�ԩX��	eڜh���f��	�Q�}��)���t���2�&��Ξ��l��{Um"[v�����j���8s[�3����ڄ�bz,���zyr�ZFe7��ޒAr%��`�e�@wѼ�8^�Ǉx��9��a4���g�^���~�QP�{���߅G�S�p��=��xth�����p�]f� y��b	�-�`&�OsJ6�ށ��3^C$�2�^]Oܲo�ȱo:��t���G+�������&5�"1#>�(R C������Z�q�ڬA��b[T�G�	>��j��SH�1�]�Cݴ,{Q�>�O��I:͊[ҵD����*���2��ӳ�+�<�p�3O�!�������\����J���-ؽ�����5�'���D�!�K=�^)�V*tG+�m����x�I�sl��R�H�E',�-��^b�Μ�P ]iz�E���ʓ��Y���'+K(���d�����<ckP;Q$I�wCB�d��� j�]�u�)-Z�W�q�#+�ta�+������H�X^�>������vVc��y�����#y�*�vj~�S�w������RR5ｾ9��v2�t��PE�D�	'X.�*A{�l��>���d�bϭ&kD+�
�]�4*�>@FH+�|�p@rG׊�xqI<�=~í�"G\O��y%>�6�79���h,�(�f���z���tɪΤjd7`[�Q�i�wMz�� ���!y�	����`��1��	�a1n�����ai�|A�*�Ć@0��/�{�$�ĢG�H���J�x/֋t����I��Y�����!X⤔�Ʉ<��n��J\�����Я�����H,?&I��7��:7Ӣ5rRe�;]����_-&��H����� P�� �}��sGaեP��m�{��2lZTo�Фhg'�K�{a�'#|�[��y�'«3����������>�?��>�8j�;�$�������65� �D�{�S��A�VF�J<��O���Q�$n�V��8��X_��:PQx���|'��K��=��h�z*��IgZ�\���Kli(g�,��\�G���ac�י�]FLʯ�̥H#T���bå�<�e�!R�m�8']�V��u�m�M=�Ca����J�FQ�L�R7�D��7�~�:£�/(ݩ�q.
�1�|�̝�R��)���C���8��?̱y}>z+~0��\J��j�6�0rITn4>�º0�L��=Gv��.�v�͠ss.E腑���E��8Uᇷ��ݓ��
��[\�r����v��2��p�T��'sYh�֔���΁�Y�uM�s�Ҭ.�j�P�d)��?%a�B��#rG{�`�>G^eS���� W��淩̦���-[���5��v�D���$�"`�4���&�n"�8E �#bTD����76�=��X���WA<�q)�h������K�Է�����,?����wDɺB!JM��#��,@�g��D	̶
����bw_�$��a���p��#_����~i�1��&f�ՉDA�����?��k|�V���q��f�h�qD41���! ̆��})�B��LF\�$pϏo��K�f��v�%���DN'�����V_\�M~��I��2b�t���+��xSo�ó��
�@��{�y��F�U�ؤ'� H��s-���D{&'�~�Se�����h�\g|����|:6�U���z�T#K0v�{%<D��;Ŷ�M=���F}�^���&g�v��'i0�|�m��L��>S���G� �&*�}QhX��tW	эΠ���-1����M!���-�U!]B%�L�K�����0��S06���!œ������D��(��a�4�;Y����=�Y���A�Wl�eY8W~t�:6ʂ�y�x�2�F� | �)��f��Z�4�է�-����]SX�~��J�O�,#66��S�%B�^O����v?k�Bʗd<�xjR_�E5���uT}�;I���Z���j�/#S��<�2����KPh��Y^�do>��:G���2����TO��6'6x~?aj
�Pt�M�qpC��Q_YB>7R��+ a��R����-c,�N���>��a�
g���Y�a���{�vk%�O�%�E&ŽZ��%�]�l[zO�+�+)i� m8!Ʉ_����u2
���	�ב�8���<�2��+=N�A��X|WM�zu������0Dvc)�~Tx0-���UT٘����7'�J��X�#͋��Ջ7>~�`�N�af=>�h�y~�L��ƞUQB죇�*o�a"�u�o�1z(!�b���u�Rq�۷�0��}�Ob��@�.�Hb"�F/�d_e������(�Q�d�&��E#�3'����jp'�M&SZ�_6�	�\��B$�X�k�� %ll�d�%hKw>���L� ��TҬf^���Z<f��޲����M�r�P��e	ි*��F��Ld����ߪ��Y�\P��}��77��.f�=���,�m��� ��~���`@{ߤ*s�0J�c|��I���[��0Rl}�)	��4�Aגm��nsi �����E.:��6�C�2��)m`q�6�\�W�\OmS�.v���@ �C�voj�*I���e|�6�H%8+;&�?%��<O?p	�NSw�]gnoK��kpl>p����ά������>N�]�eh�T���HG[ɕ��-;�
�k@:���	��Pb ���&P���>��3~�7ŉ!A.�N���ڧk���@�E:����z�9Z�R�6t��}E)���m%÷�
��c2Wn��5�u(��n�u\��n�H��=���	�l�%���iK�����i9*���u��K|K�������ӳau�،�Ϗ��K�Ӗ�㏈>J��H&��ѨgA=-	NTqoxLκ��0^���_餯�-c��e�\[ޑs ���#�5�����O{�����������e�Z�*��~�+��c�?��VX��I���Tc���WeI'o�AMlml/J&���B��0���� �vL�j���ĐD_������šJb:�;C�~��۲H����	�~���1Fɍ��O���S%�@V{8j6�N�g�v=\���W�y�`*l��҆��$y!��_¢A�&�IC�YS?��!�1L�a�O��>��I�a�
=��[����Z��j8r���o�w2���oZ>ߐB+dpoM������������Jf�J/�҄'��{M��G��'o��?9Y���_��Z�A�(�3��!���)�y`�r��.ˁ>�b������Ć?��w�ȩ����w�QI���HךO�B&��ǚMsLͿ�J%q�ZA������~ů�9"��$�痝龍�P�τJ�Z�hM�\���@�/�S���:��26i-���!�0{��3���5���[�����}�$BS���]�dng��&�-#�N�� 	���P�
���3�ٗX,��T��:����}��Xۋ*�+�i��ai�+�j��l���֪ӥ���@u3��?ߴ�3>V�5�����N�0`<)é4Ys��^��!/�����c#-�/"iՃ/Nӽ��!KV7�8��U���	�=��7�;�_���}B���]���@K�2�Z���同>�$`N�(s�2^��$�n!�Aӫ!�X��)�\ZE,���Eǚ����k�M��֡Y
2�:F�z��[������Ckw��]測� �֖�'��q��U_�Xڌ��R�EF�u���voH��|	@7`E�7�>�Z_�¡�LA+�H�__q4M�NPbS|-�2O�r�`�����,��tn&�k�P���ϊI%\����k)���~��{��O ?�$sQ���ptv�~���"�i���/&ބ�º$U8껮�S�~w�壳9��&-�,psq��G7b�U[�l�C6�"Y�U׷l�e���Z���ʡ'p�O��Z ��F$jm~����z<;`������va 5XXb�ǮigG�7�!VG�|���1�t<]�?�F�;n/dv��UO�Q�w�jE�~y��r�8���$y�=�6�h�pD6��h��զ����Z%"fO��@.��Z%�zbO[����f�a.��J���bM qj�h�S�4���8��� �=����kRS��KK
g�A��g��Ƙs��0��ع3ou�-cv�4v��w�OYl�����˔��u�5��I,%�.s��ݒhF �cʎ��k0�~�}n3���������N�M��҄���D� [��"1���/�S�pb�O��4���R���	�q:/�%�.�ۈ��Le���%K򥹗�m%p8h�@�"��}J(�.�W6����Cڵ�B��Fr$OSZv��,굻j]�Liy�R�PfAt�����m\���o�(r��¶��A{M����K�������?��B%��G@�=�{{"����҄S|��Jwң/�fHr@�{�ϷAM�6��͚�G���U��.
_��a��>^q����)��Ϗ{��]���}uc�W�y|��;�#-�F�Z����rh�O�K�ڴG�޺ʪ��3���Q��R��C��$f��p/��
����ud�Z@M���0��[�����
�Ⱦ�W%o��(��Tc����㡵�Ɩ�Rj�&mΧ�#)S6:��*�)'v�o���U���E��M���{�s2��Q��C&��f;!��Ǎ5���l�z�°�Q�	_�{���\i��A�B"��w`��-uG����!���K+j>��ض���$�����k��6�*>�����\4i��g�6O�,y�z�(�L��@[��%�hnv?e����flyf+��얥$!���OjE ����e��_����$É�,�{�^!�(-��Õ!��t� WF�(^5˷���K��j/9�P�7�|�x����}oĔp�5D�˧���^���_А#�,o�t��`��81�6�i��I�:(:�,���]i�5�JO��^"T�]��q��媘/ލ.��;��t��r���� �a%�3�H���2�AQS�%	
z���V�
��F��v|�ʞ�kҕ����#2�{���ΊC �j��obO�j�����&��6�� ,Qkqx\�c;�č	����p��x��NU�F����SsXo%��W�s𒌁4]���_N��)���:��V�_�Z�B�m��G�3��;��z$�����9I�3�l?�0��j�����vbdk��&W�Z�D��g!w;p$rJ��������C?"��A���9~�`���pOFxj�	*:����n��J����N�u$��f�9��������W�$�Qm^���}h/�(�
��-��.-�nCX�ދ��gL�? �C� ��� mQ�ObL���0ļ֐�>��i&&��]$(��R��1��@bᩀ���
�#Q��Y����AH�j4�]:��^��n��<�|�[�f�F��~)�h({��<Ό_��	�>�IF�ޮ9|�xo�x�g�~�z��,,�u��W���7���P�c�Йe/K_kM8(��N�ȓrJ)
��#�V�<2n����,��~n-������"��������!�:�CbDR.��*/]|cpSNd�����@T(��P��)BTX^�2��(7ڋCm�'���b���E�����e*����;�ܔ,D�p��K�;W$�C�Q9�!�-���bpV�pܢ�~Ɲ����?�pI��,`7��1n�[�L
�F��8�1r����>�����-��n3�}W �2���a[�V������#�V�r�%�.0Bㅃ��@D�dM|5$�fVxJS:��^�q����Hl]G�;g�� k�l��,-��I�t%2��>��Z܉�^���P@=h�>i�I7���2�]m��i�bMn4$[7���tw����~�����b��y�K~ү���*\°�爡R�[�*VM��*�޽�L*�VO��DE���H����8����8�֩P�3����u��>�98h]�}��9�p3ׁ�J
$d��7�y+����NՁ��1���s+I�A�!�B}�b�b%��<�zßE1�y��BOVθ��(���v�ǈ����I�o�ԓ9��4��M�90�4c^���>g\ʦ�k<�z̞�q`5�B1k�����W[���z�x\Ę�'�<wv*�M�ȼ31��z-�.L�~���)��b*�-q������<�~:u�Z6��pt�6d�]іe�V����g�#�%.�NKf�ҹ�k�NOq	�9���M+�.��u/8
�H'�����yK���<,��A*�a@N��X?X�G�"Kg��60�$�i_�f�Y
�6�Q��䍂�P`�9��®}Q��F���Y�!/c�xʕ��/���d+2+:x��'˹d	��q���^�����%MFr��]����"�#�X���*�P��açI�*i;��3M�k������+�y�B��e0dM�0���9*���'�Y:q��3b�B�r������!������,��?:{��ý��LU��.���"�u�~uӞ#�J��f��#8�҂�U\���p�k�S���l�xM7�(=�V�޲#��!2yG ��
WRj�N�B��j��W�ZjE�r�Ē�`j�_��-�q���=,�D�B�o�	�@u��L^7X��ҽ��0����ռ>X�l����c��gE�:���;���R�݌4��w��]:u��#�I}��l�W aJ���ܿ�-�N��^{�(���Vv��x��	#����;�t<�E%��ܛ��k�n:�����q���nd3H#�Fl؟��d;�fp�P0-}	j���#򧴦J:EE�6ī���+��"b�|⛟�P|9��s�g����B@��h�n�v ��n	,�=��M��ڟ���$����H��8��2DW�o0���-��E;R`	����<7Y8�I'59R��\�/���0�}�<��h�_q��y�-d�]��14�K������ϻ�X6��Ҟ�gi\�~�CN:�W���X�pNz'qԨ^/�\P��~�<�3n��*]O+�q�۽hͥ���Y/��H���@��,��2�kx(�'ev�V)P�-�r�֐��'���e�5�<�������9��ܡ�K#I�u �ւJ��W��!�����j��'F3L�Y��` �c�0	[kR�-{�W������_5��VF�wP�a^p�~�ȿi`Ւ�iJʤ/U:8��i�LG�j��1�K����[+R�%�J7}ڳ��X[���!�������O�J�d\R��>��j�
��q��#�1���ȯH�����y���\�B}�)\b�\�h�;nO^����4���K�I-����a̀���d����F�D�R>*M��p�h�hWH�{܌~9`�f���*P�p�6v�s��?�֝���B��x�\�S�	eL*�T�@����X�rw�\A�_�H䗒m�y-�ʮ�6`�}7+�[eK6�}��1�h��"M�T]R��Jl���P��@��	Ԁ���V��K~t��K�G�`Z��p%��o$ߎt�sN&��2�d�-B�}t8b�ޑ_�Ƴ�]������U��ьx`q��HF�.-���E,A,=)���0i��q�I��ħ�6�v�w��ȑrG��f6G�c�����"D�������#����\�n��Z�j^������/����)�? �D����cu�u�[D��֧d�pP;1�'����᥷l��h25�P
M�޴��A�2�<�����b�Y�0�	�� `��>߇�pϭ����u��: iL�ӨYu���uWy�XjXp(K�B��>��u�2|�C��l����`A�F�M'���C�T%҉��4]?�Hfb<jF�tA�RO5C�h8f�o�ӊ����Ĝb}=�	���X�k�G\�Q[�(�<�5~:�Q3ڍG��{h�G.���b�	���A;���-�:��=�~2hs;4�z��t�kJƶh�4d���.%��tU��O�m��,Ҁ�Sc�?4״��/�&�]�'x1�v�XTX�X�T����\�x9k��#!�M�������CưL@���W�u^��x�J�E��^Z4�j	���r2�vy�m�%Ƨ�\&�F�a�yfu�9Dq�_�i|\��R)j�1������7*A�A�0` #
0"��h���5�(��9���޹.^mL�N�:�Y�&�na�g�EV������j̠r�����b�~b��U/O�ьU����x�(/3>��ӷ���b]�=R��7!�xd*��4�SP�A<9�L��S��4.�TjS���~m����6&MB��i� da6I]��<����o']t�z*h���
tZԾ<����g9?U�Zo���aU�LB��،��e��	t������Rn�'�����"ec�Յ�b@Ov2F]ŵbgs��[��u�wP�c�~�)ѶE�5q���[�]���V#K��h0c���� ����,_ �aկp�p,�������N̵�x�,w��F��%��6�F��吠���#�����I��P�ԃ��5���f�Cl�ي�8������o�e?:NZ�T©/	 SJ��Ys@�^���|�>J	S�	��d�Ħ�_���N�l�vh"���?��7����L,�A����-J�h��ԋ��~a���b̦� ��Hc�����̲;Fv�� ��:�x�|���Yp�|~��e"�L�J��Sl~^��1�=H�6����9L�y�zZ�^�و����ݮHS2(
BǸ����*LB�3�`l�}�R��$���S��=��Ѓ2�d�����JNmk�/��8�X ��5�]�N!~'>��!�j��{Z��X�)���};��K�R����,3̴��n#��;�|���7t�;/_޳;B�d��b$H�$�2v׋�5`�I\�TO!�K[�zϨ��e�&��5,��ާ��c�(+Vӹ��ya�[��}���Ռŋ.U�Z(fD��o>��/;Sdv`�6?�>"Y��n��lt�2�Q85�՘Hw�b>��bݜR}꡵�#��{�J�����m��K��s���_������훡@�����sm��+d3��=~�J�I��3B`��6��vҩ�=���91%Gq<��m����RW:!�H�$� <oh��	0K.ls�H��0y#f34���*U_�IɊ�_L#�\��eɽ1ÒA}U!6��!U��d�U��ᆧ:�s��$����<ԚBTH��=��v��iBUQ������*�PI�W?������9�����}����-%�jXu�O�Ղ���(��X��z�7a�Y�,�۾�Fh�BwaF�	�6���*��,�W�Z��ۏ)�YP�,��~(&Ut�܂X��!4f��_�]��.C����DO�Sp�rӔ9���S0s��9$Rk6 B��R�6������a���dRm���ųʯ�e�������+kRr��D��f��s�n�)�_p��J���А��dLt���̬�i]��S�S�h�v�S��u���o����J�O�ّMc����!Q�2*��-��p^t��r��#ppz7o9��5�����8�^�ã.[a�ϩNp��8�v�-���)�F	rxq<���0���>��O��dȽl`[էm�ih�J�4�=�L���/R�Ii�C/)!X�0'�ի@�+�M�30+��cJ�T���$�0nr��%W�
̮:�yl�i��g%_��3_��M�vED`���'$�Lj&Tr���aH�p��[�%�4�+�����o�sL�a���a#
�������x_�4���g�^H2G�:�����ȸ����;�j�����wY�(�q���e�}p8�Ĉ�?�Q0sa�tb� �w������W�Y��#+��ӆ�^a���䣂G*��<�Y����g�>�� �Y�~�u�x���$���EM<bd-|1�c��l};�E[�m�FH:d�$3,%�]nW�`;�X��}>��8�G�#�nt�`�s*	w�~u7x(8_���S�܌��r �F4N��SlcL���e_	Q+wK��~+у�tI�7'���E�mEf��cЇ%�C)
�-�p��1�O��ԅ��U���Q�05u1MR/�5`��}/�����&����d6��n��o�����\P�����!oq,�_$E��	���I��iNt�727n����<]�A	��:¸ZB���������R��<���BϤ������*l��d[��:��@{�W?�d�Cd�fQ��2 �E��5֘y��	R�Zm{�a9�ݚR����r����s)IlV;���k�"�C�Ŀ������2yS�<���+�9ʌt���/
TAy�Ц�ˏ�_�4�������2��v� ���H��"��H���)��&I�w��@�P��{�ժ[�PK���ڂ b����|w0� �o�t�w����n�.??4	��L�l4q9��#�io��"�=,�����@��Z$�n^�p̒-.��Z;{E ���y2�c!ɢēt�U���;�7q=T@�{�ܜ5�]D�u�����ݍ�+��԰�r�/ꏨ'�y��ό� y�C��-���y��_������ק�9)|�5eL&���S��BW�rSD���������$^�K�U�ޞ��P�R��rN?�p~���8:�2N���\-(�)��b2��.�b�����ܥ�un2�6���݌�t��gx��]ʂ�/�'_�|��9+ف��@}���c�nR�6Q�/�̩�u���0�J9��Fx����'���g�0N�ՌH譶���0�XZYAD�=���:@����l�<�4�F����_V���~5�V�Sߒ�S��o,�W
�1� sc���ӗ���*Y���{K�Dw?Xi�	P�w�g��}0M���8�%7l]�����T��H�z��V��.�b,��6�sE���$~�����;p?��z�M���ֵ[ʋHaE�$�b�����׭���U���k�s�>D �i����u
��)����Y
ֽ���Fc(d�l�3Z���(Q�N�E���6�,�K�a�'�d�Ƶ�qS��l������K��!��Ĳ��8�k�d+A*1�^�A.x�
���G������悧�䚅�}���d�0�Ʒ�<r:h�A�:��)�&r�=����E�S-��S�����~`XY �7����JԶ:��w0�2k-T}���99���3�q3��W��<˚e����z��	2C0���킍�;8G�#	�Z_1�yRo`h�=��S@��T��&���
Oy/�������?�����~S���wd�jzR ���ׅA�	'���V�:��� 7~�7���e[c���^8�D��~�_�Xp���s8�`�x�H�$D��@�pt?o� ��x�r~�DK�"�M��/+�>�0�ȕXz�_����R��U0Ƙ�a���fpK���A�r{j��93�L��	o^��R�j��I[��\8������>�.:u�8�����r�ݿ�h6��"��g�e�$�YК
|O$LN&��'=J�\�jă���q
�V2�c���[%ɮ�����π{N�婈f���mh������=���-��r���*�J�bï*���� ���ނ� &�hXuUج����ZGH[�о������u�rg��x�YX(L6dB�C�:=Hi�m} ]^g?T�G)	�a��ݡ
�q��>���\BLM�Q����$a$2Zd�@��/��hB� ��4�C�OW�:�L\���%)�o�m�*jd�b9��l��%�2"���Z2v�"Ix�Y��{�ar0k
��2Y޻b��	��	��c���� ��< ��iA�ve-s���>k�����C�T[��M73��>TK�8�D�hJ��P�Ňo��-�I�P���������?�ZU��Lŕ'�v�2Å\"
q���djИ:���^��)ɤ_4����x�J�R��~f���}�q˃��������W7��y	Ƚ�񶎩�����2I�2*w"�oU bDR��#���L�64��+n�bb/s��H�Z;�M<�Q���i��!i-�7!}.
K�M5�upJmB��
E'��`�e/��ڥ%^�E-�*]�_tmB����ˤ�ޘcx-9PY(� u��꿎������4p�Jף�3��8~��Ӡ�(f�U�p�u���rry������� .\Oma�Ph31N�Dky]aF��I�\���<�D�b����7&C�����k"��|$�)�q����U�Q��7�s�.[?3n��5 �'U��A��x� ������y�[5�+M.E��mh�ȶ��r���Y�L3l�䘭Q����O�^k'�味sֺN��hZ�vX�ۚ�>lE�xs���hX ��/;�6!��jX��|�׆�X�d
���yG<����yKE�ȃ3С䠃S��(D�K{���ja���`�т!�VP4��g"d�{��=�$��c�/����n��D�G���B��C��2|%[y�g��i:H=t����UI��旁!�zƸ�m�0,�kro����5�-���hn:��t�$���^k?���a�/<`�Wʩ�%��٨�_��nX'
�X�'�ί��۔3� �
D�V叠�)�Ϳ3��D4��x0��A+��jD	�&��艥L$����s�%{cOV���k��o������(��E$�-����R�<2���O���A۞s�?�D7<��@!5�{�-)�R>&~CY�����GW�`�"/�S܍&�a-�1v$ԘnP0������,�y��?���a[��O��W���5�2.����z�,���C�%#�/A�AQ��s�Y,�v�f��?�K���# �x0}XW^	V���l�XYW`xgO��5�1�%�����4=��쵠~�C�:�FT��G2Gh`L�[�])0������xRf��|["�v+P&�����T6T��N��AX>70�&Da4 9Y%eeƖ�Y��kAw8%xy�9���ț��;i�n��,5F��LAa�l�V��Q(wGh��K�\��z�<ļ�����K�'�8��bBٮ�Ż��L�����J&��s�&U���[z먧�11�+��~����e������ �V�*$&���o�b��!�Z�x�@��7��E+�l�g��1�U1���Q_��H#p���Y�
߫2�
��_:��/���*���gΈ
�X��EN������m7�
��#nP��G:�8}�Λ�ɰs&=a���9-���
21�l�>����
'�l�KAt��K�P.*�~ 
��H,��������e1a'
r�u���r��E��*)�=e���NR�C��LǄ�OX"ul����0�&�j@k�(���çy{qW��Z����{��Y��+F�2�Zʽ�N��m��T*B@�h�D�C�vZJO�HZӕ���>h}��"���߻���a�<�|��s��@W���3��|��*u6���.���[k`,��X�S�Q� 1����"���iki@�1�ZJ)�����(r��c�pT{J�D.����]Q�b�,�6�e�x5����2��=p�t�i��9�T9�ī7g�Q��*pc�\N��D�$���$�[|�7)�Y0���iǚk��W�:xS�d}K�Q1C(}{��W�����y�R�:��E0��C~��A3�ʵ�B����ݧ��7R% ���1A>2�~�&@�֨��|����N��=��P[�ALR7����gʱT����,�9�s��25�`�_ܿ�,�ܙ]MM
͊uz���O'd��5�]�kj��&!��#о�|W�'��ߴV�.�H�fA$��:�́2�����G�Yf�ӭS,�; ���z*�	�����I�u�Q�Jf��BvS�����T��N6�j���I�&k��k���w�$�ˎc�~����������Y�(���� �+��,=�-$b�~���� ��.� quKR�ߙyA&O:h��ՄmmaU@~\�No�n���Yg|q�)Q����՜�-8����d�� �C��$e{�p}�Z�)�B{-���>3�w�|� f{�!QY���EU`�*� !ڴ�"�t ���q�s�;���(��T����8x�g����ت@���Ƙ��RKkdz-ɵ�������=$nۄ�,P�K���ۤ�кɐ��#�ZvR�m��HU�ѭ��d�n<b}��O�}��r�#l;J��rzNVH�Xt���2�Il�'WD����)�3�[/��)��$[�vd��^�����B�N�J�޿��Y�*� ���qT�-$�V��nd�_V)�q ��$���7���|��'�j`�wA���N���s5 ��1���V�kTS�Лp�2}�܋�D�f�f��v���²�p�{�vډY���w�d}'+��đc�F4���
�m�����"2��i	�Ʈ��1)�z?���Z5�a<�N{��h~�d�}m�W��WV)�∩�$��Rvj�5}*����P$/�<��q�"5��5�b�f��'��{�r'�)�n��B��N�K\b��T2���p�\�U��_�t�z�$}�KNrZ����G%�k��z�mG��t~�Yi؜� �.IH�n|��7|�� =(T����	h-�}�]��G��8�`ڐ+m�-�ѕ�^S��eꫧ_�F�  x�?��:_9;������[c��v4~���
|�+v��~h�J�{�]gfV��^���]Lw)5�!�w�F���&QL�5:�G�rd4j��`Ws%o�vʦ��)Ub^0�m�\�;�3���p���2^˿����
�,ɋᠻY�ٷ¨��S_3�C�zz�LąX���Y,����=��������� ���Q�h�Y6МѬj�@�AV��u���|1q�o`���	56�{�b��/�$��*���������./��R��p��}�G{��hI�8P1dg3 
E������(�C����)��-�IL�W+�@A���:S��F�;8���8f�q�"k��<Ԙ3��z�����s�Q:�������.�+�u�;�V��U�*5#R{:�Da��d[3�\�fѼ�9�O���c�!V�9�a�.�i*:�Zx5��B8�Q�6S���y�˅<z����sz�t9��]t�d���aP$3����t��{�+f��ׯb���O�a�ܢt	�"�½�o�|>k���UXƦ��
��:����e��x�H�"�]E_�S ���Ũ����V��X��DS��oj%S�Mɸ�5�L����|r�(�q�͡GD%�a�Y�<������]7ۖ_9�4H|���N��t;ro�'ЖƗ�֛сFH���-S�G���҇�9Pk	v������V�@1�2h:�/���D�J�og�>�-��R�]��=�O�$©���A�����Bi�k����u8lJ��.!|��)����5N&�sG��P�i�(�6� ��|gto���,��tC�1y�,�@n��# ��2>�<�'�3���d���S��:k�y���V��R����w�ő�;����u6?r�J����Q� !�VH�6���]���N�)+S�:���������O�i����sNP�H<u` 0WI�#<�707��|�qc/o*�-���$m4ܢB2��d���F�>�pv�lt���G]W4O!��5� ���{ւ>�7>���4�i`�)�yls-��?rp���c=��}�C���p� ��#t��� �*p/!���n`����݁���~�/al/�|q�0կ1�y,\�+OƝ��d���9�L`���K�>W�if�wc5��s�全q����Yp��ϛ9��;CG`�PT��U̛!�/�2f׾Ir6-��:�����!~�����`S��N�H��î	�l+���3_�`�g�x��Mb<n�[�x�u,[��o��=Y�kz�F��v�j;r�CJ~5�?�ltL���Iݫ0��K���)�+\^�_��J��<Ds�@z����H:q� ��4�Z�u�
Ks��4�G�/�ܾEs�
H���|e�,R6/�])�Fّ�K�x�r�_yR�z�j4,%��^�;G���I��{H���W���N����q0�*�S1������3����[vt�e&y�|"��0B�kҥ淋�.~���q�ymyf�z�둂�ν����k?��}R~<
�=�B2��[��ӧ=~�����Gg��%��J��clX�~r$G�n\zL���[���:�?�CD�jT���=�lf�j��<%�4�����
0ܤ>��/&��}T��1�]L��{:�s�g��ʾ�O�H���S�Λ��3�B���W�����OW��'�������L0R9+J��yx�YI�CK�d�jyZ�ZVl�i0 j�j�^�S7^L�Cp�ͬ�Q�貪P�µ>2��L)�L!�OƵ {����u�Y0b�n-��s���f�ݚ�{̓��#�a��龟�l�S�w4U��J�MtcW�7ҋ�0(�w=�=X��1�.:�jd��#����4�_D~X�nԂIٿ|�$��Z\2�̀g�+�4'�(KCŧ�!gP�U?�@A�H�'ZX�4W���G�ې4W˞Z����`m�G?��o������\F�B�p~uT9��������鉍�ģ�L�\�7�@5^���~W�oڎ������V��vU��ܲ���"97Ct\RD�
�fڏz��2+wӢ%���Ư�()h�"8ŋ��yc�����p;����$"|��"��ډ����aP��\j*��o��e%���ʔ���h"�JNp� �V�x��[B+�?�l�Z�����	 ����Bz��Q�}Du�� �{Z�F�������0��}�h���᡿�j���
�k���O�9�U�:27
��d��w��u��芭�t��,�@�P煘J��ߣm�傼�}4�{b�7DI&���,� #jT�u]��e5	���P.U ���qٸ�8��腲̑�4���˟�hL��pٮQ��uH�FT���)�cL?�`m�H�{�"��1#6J*}'�y���>����q�/��������O��+���7���lj+���L��j@�ȵ�X��u:�B�!��*�@G�N��έ�?S�����[�r���}����X�W����0~��BL�sv�T�t�Q�گ�N$"�.�����n���U8�1��Q `[�e.6Z����ז�~�	��«�&�v\����.�g%΂N� �����A��%�Pk��*#���*��v�Y$ri"�`B%�;yQ�\�-'X�����%V�r/��]z�4g��%��0k۪�H�)_Sro�,���޹��FzH�☙�W�D�ޥt�(`BH@֎���A&�9s�W�I��&���!c��5������wL�$��6u2��7
��4R;�>  �y��,��$[�u�T㻈�?�e}3��i6� Tf~��klW�:ko�-��>�^��nK���?J��J|8����#�s�f������|h����U-!�8(4����1DPIG�
D�J�0��gE�����E�0�5���l�Kh�H�8j���z�+������+�?z#�/����:����	J�$$���S�Hi�T2����#��I֟v���_AV਽=��2����,�T�V�P�kN���lk�%��X�k����s�/H�'��]�=�s[Tba5^��l��m�XQ�������1�1 i�Z� M�W�qL<���`V�ҳw���m^]33�G`�Lת3;�	�nݗ8�v��L��ȲH��bۈ2�ʁ�� 徉E�lU�$퇿����mM)�GGa`�VR��wS:�g���bc���V�&&�]�?��]X�\���n�889��=�dD�Ntg�~����ni9��&�<S�eH��8�Z�{��k���'�B�����6L� �-�U���g�`����W�Jr�@�X���(�s�	ģ�,J8i�t=�!e��T3#XUm��w�d[��I��c��yY=:7����Q�Q0`@�E���pUO���u����ٍ�<K��I��������?��:K�>M�<Z�v)�{��?�y�eW4�<.�����<{�OHq4�����ȡ�h�yW4*�Ջ�~����z����Z��S�r�p_���J)��8��c�i��?]�K($+� K�E*�2Ŀ��q�?���S�U�C�xd(5[����A`d8���i�at��h�S|���c��T	���3�_�q2��y0�}p�
m�w�aeO���,���TMl�a�#�>ިp��U�,�Ul�Y�6��-WL8%<=�X?By��x�ɲDr� ��*؛L��F��}:�<䬄G�>W�ǫ���H�hl��\5��J#`���8
��5�k��a����#P-�G��~���J�Ex�o�˴9�i����������q�Q7h��`��bu�O-���,]���{�����0Xm?w�c��>)(gh��1�b�����q�.��w�k��E �W����2��Q�N�%������G}��"��\Pn-�מ����qc�4��+M%YD��R�H�6�����@jZ5�4��aD�˽jǃm����ݟԻ!�ۋ%.�d���t��+3�i� T{`-룥z�Zt�א	"���g���u���4Q��s����@���}��iڜҊqD�
BU�<"Tf�c�i_-����\�R�S��2�����pK���Ni\=��4�9�b�o�Kl����ik$�i�|���:�c��&{{�ʒ�.���O�y�X�ib]^�y���ܻ�.V��DR���L��ߔ:�^p����	�7]����S���V��~�إ�h����s���jh�P1Y�c�~
A�YQh�NJR����Dna��3<K���ڳ�зz�_|�C� a��ф��)���dzA�NG�������G�Zӏ��k5�Bo��e���Kޛ?Cm�3�'�'I��p��}��D��R;g7&��}8�@\*ǒ@��Z��=`��K���^��hq|�1k�i`&� T�?K�AoH!���șq��7F~+�ҷ�"_2�J�15�8rv���l�,v�ƧԸ6�lso,��E+rz��	F�hR�:p��3 D��U����+>�y���C'Ԓ��P ��<��u�9	oυ�k"wHb	����k�eb����$�Ba�>�<�歳�<��P2~8R�D���}a4$tq���	Z�i����J`¬[E��&l[�
�4	��,�%.�i�ohť�4��������CC5y�~T]�����cL(!�i��"�4[��I� ��!� �3��^R�u��	)ؿXdh��΀n��n�{�[�yȡ�4I�e��Y�,�f3�Ho�
Lu=��&�x0����\���������j�m�����
�N�j�J��e35��\��+�2�Ϙ�,e�v{��$�KG@�p$6;f�vI�J�ש)-�%��d�)�8�xPi�����(`b��NdA�@o��9@��vT�ض��*_�c�}J}�\o:w-��h����{!6o�ׯ�����\Ʀ�)A��_�-W�[���1"V��N��҅�p,�0�5*�-ίLu� t~�/��uI�)ʵh��_L6� e��'���(��'3��{j^9�S1kntIJ�I��G(fވM�˳��$8��,x�:�Nޖ����繱&��A�G@CA�c_�\(������Lǻ�e��a�+�ns+7�|��@��xKG���{Z�#
�R���f�\�ܕ$\ip�`�8�Տ�`���y�6�&���%�%���e#�0
����J���\���=��'	kH�~�C�L��^2h-Y띡Q��$�UG<��$�ܵU����H<F��_������X��;��_�8�彐͌.J6�P�2[��f����y��?�o�p=�pݍA~��;�c�0f�	<*md�/���y�Lb�-�m��Dv��cS����ng"�(3?s����������q�.gz��E�t�m�@����M1*u�����$kl}�y�y�����8����&̾)w5����b4�=쇢JL�"��x8ݺ�etŌ7kK�o�,׫�( �Wgc���*�H���K5[�$z�Xzluu0���92�����7�s�|�9]�Q?+�Ю~3�")'"�.��V�O��J����0?��+��"FNw�3�8���Tͺ�pu�L��g>�!���h5O�ZS8�#�s$ѻ�R ��|�c���-�
��9]��8�4�^�râļ�2�J�ך�YV ��D�|X֯OF��ۡ������2����ߌ�g�N>�L���y���d>Tw+��R9�Q�;�*#���k�(���Cx�Z���$r���û/���[	�����~����>E6V����"M�W�;�fB���p�㈙8s�R`�g��$A����'���!`�V	^Qf�������`ԎF2��"3/���ϊI��Y�uo�n���k�{�X}7>��N�SMg�#�*�]�%�i��?��#Ҡ��̫�F������$t�#u2��d8�on[�cې�>�is~��Y��:�otd�B'AE"o�l�6ah��?q��l��{=���4ĊĀ�X�3���P�`�r6�-9�n/n4Ӳr5Y墆8W��Q!Y�u� }���gh�UI���_�}u��B��`�G��cEG����ߚ���[*i�ԅ��@}!0>k����l�E��^�5^�a��^�؄��h��g��?�x��eW��q"��o��ny�㫼p��r�i����`��,�Xћ��=�R�{���ŃUE�T#��Qf.�J�c���m�G�[�Ư��K4�AȂ��4��?��ް�������3��qE抏�)��^Fz��8�Ư��b3l)J�Fv�~��~&i�5(����gb6������0�J��Uj'yN��m��S��<�w��P��`_��IGԾ������^�8o<>�ds©:��+d�����?���C	"L�g=3��&������S��Y�y��{�4#��DmaV;_���Ib����G$&�`�	E�jsf˫<7&l��u.��r`�}N8��b͎s�OF�ͧ��Dkͯr�3��&Б��y�s����5�nc�7�cY˻���u0�Ö�O�&�ڽ�YϏ��V�c��q�u/��φML2ۻ_fh����Y,Ŷ������֨����աd��e����H��q ���xL��X�
gzk���d�{E��ʵ.X?�й���2s�4k�N&S�:��A ����>"���Sd�����K4�_fnN[��k\o�v--NO8�b��  �\G� JK���H)|h��#��C�!5*Ңf��j�$��Q��T%�Y)H��V���B+��rA����Uf���$9��r���o�?���wՊd��~}�Wz�WbN橩�?V?�𥌙��69	-�ӷ���(z7#��e��jS2ߒ�&�>�WIG�QL�<�<�EZ�*�D@Lm7��n3�y�������U{�YX�37���}P���R~�k`�/��iƘ�yR>e�Rj(�"��W㇧���Y;ʪj0����#u��忑��6Yߝ�������L�Ws�;r��� �?�lR$i@p��ڢ�T�W���>��[>N�Q֭>�eQ��ܡ�����C�f�+E��������$���pJH���i#+�n@T34�V&X��M�	V5�ͷjj⿰6�%	^k���#����bHD�����af��o�0�e���aQz�F���fsd�:G�~�L�h�L]	<3�2��D�q�a��*=�RM�f]H�+�$-״$ނ-��e����8s�qV��AIk�J�)���#�>�e��|~�t��P̐xge}��Җ���=��#BE�%_~�.��,�6���/z�ˡ ���i��@�b�h��n��#�Q�4�x�����v|��91�4��y�����"	;A�ӆ6߅e���[�����~e9�:�?�ם�VDe�QH��.:;��u��خ.4��?�T��M/!�>��YV^,���=!��ޘt������@��C�/�,R/>?D^"�Td��<w�7�>_s]��a�t��DJ�B}�!� �ϗp�O�ϼ��5z2�uf軁8��4WBz���}�����C��٬:���E��2��}�r�����K3�A�P�_H�R��Ì|��5�ו�0��ܱϳG���?�yR��G*�[u5UB�J�IR���{#s_��P)ɹ��ʿ�~�=�c��v�fn����l�^��q��s�lOz����� ժ���U�ҍi��f���z��![�k��K:j�,����Aز����o\�0%�d4��&F]8:��7����y���u�25��߁�9�D��,i�&6�g��q�'W�ϳ%��d�^��m�����a��L���K��b��������FMW}\��a���T��?kSF�bb�l�9ZQfD(����_�T0:�&h�K �7!�>��[��.4����S�Q���_�?:~�E��ν���>��F�<�75�������P=R�M?s�ߙN��;X�F�{/�j̃�~���n�*��He�Ԛv'ǍX��eI�1�k�Z�AY�L`���͢���'L�	g��cRｈ:$�>dx/������~ď{���%g�t��̨�&E>�Ѷ�cX��M@��_ND��E�����HlT���9-��?���K�l�φx0�@�k`2_G8N���K�$�#����{Z?�+e�%�3��J�C;ˋ��N��.�Zj�����:`=�|eQ�ᶉ<���m�k)�U3`�g��y'n.�B�"�?�{���T]*O��ѦW����j3���-
�I�͞B�e�w:���@�ާF����h>ڍ��k4��iqmU�-L����L��LZB�+��HjX�x�5���U�8��	���PJSh_��֟6�*b=�����x��;��wp�t�E�q�&���Zy���|H���gj��I�����3��v��֑Si��~ckvq=�_�r�jT��)�<]�z�^=���b�o8�S�rEXP�X���B�FM��]�sn1I�������4�ϝR�D�-4X�H�S���Mc��x�ٸZ�W��;�T�Ds���>^�⧬�_�fi ��ߴ�A�e�@sE�T]q�Q�a��?��a��-� ����էK��d��	~Ni��X�I�p�I;�Ϙ��A�n�b�1����i��o�Z3\��^T#�����Mpg�4m㜔��s�*���׸�5?�89˛�b�f?U�-��n�)�{)iI����<<���ǿ�?'\h���:��v4D]D��
��5 �9������hk��dH��P���a�ߨ̓�HM�\�_��,��p�}�����s8���g�>L�|T
5S���{?<�Ѵ�����ta�X\��qݦ����}K�7����g]S�0E�v�of�cN&jɷ��+� }Q:Yb�'��%n�Q�qԢ��m����]֏�, -��O�$�Ѱ$���������+2���V��M���dpa�N��{���CAN2��N��f�Z�8���@Ue��M1��A���nӓ�im
ƨ�䃧��ar��
�����?|��`�!�a��ԁh�!֌�=R�~�>��$�1�?ɵwR[S�ŏ�P�Q�<��En3���*�31rI���c�����{�_DH��ܹ��"��(ޠ����_Û��g1/����'�m��2��2�'^�����[x�E�k�^��X����;�H�I��&	u�RԳs�^��-�mj�j���0�^h�a"�]�v_F�+)�%A]�nCO�V���m����}X���L����3P$�qF��ý�����T���4�-[���ŀ��	�-�A��%�����"�6U�nr��]��=�/��M'���yc�K$[��k��󤦝� ��F��zȁP����_�ya�c�O�6�56�Cō���3�0)<�fc��Q�'=������(���ɐ襇~1d�b�8�*��	\�@a�����I?19�:g��>�����r�3�����'fڰ��*�z�����(�� ����e�3�Zc�v��� ۡx!�D��C�ҙ�ZG AR�mf��2m���)2�|$����Ʊ�ػ6��Ew�Y6s5^�`�t��D�*���B7�m( "����r��<��75�Ń��df�bP���(s|N,�6��� +�gI��͟��>�� �Z���=���U^8��喥��ˮ3�Ns}�޽4����V�R�1ʶ�:�Z�����,&�V��� �*+��o%�PS�U�W5 Xi�Wv�{���	J[�z���H8q����V��T%�u��J�(���j�x�!�&Z�m��h��fܥZ���Ux�9�E��Fo�1a�&���hd�J����g6Ƕ��H�����s���d�7L�*��j ��tn�����վw��Rf�g�&�~ZR��J�G�I�y��������F����*[�����w�$"����!^@�O�v�*^�׾��=PE�U� ���%�iu�eQ �.�sݑ.�r���-�J��L�$Y�W-�����{�\G̑�6�.uL�E�h5���/�ej�T|���a����Ĺ��Q��=�{�
ko:�����K`�IR�<b�r>���jӮa�,�Í-v��!�X��з��}e�A㷳����+��{� .P>�ě���c[g$�*�����_/�P�i��vn/y�`S������9��~�ψ%�
ְ�"a�J��Uݕ��C���"�+���	ġ{�����S@�ᄿ��e�b6���u�>�:�Va=n�`���KjY�O��#��B˦�����Aj{���?�ˌ�}�"=�AY'�A~�ݭ�O��P�a��K���!N.�$x��t5����+ 1�-l��[݈UD�[h����=����gA��gQ���o�e�w:��G&N����UيS_^��p5�Lr�0g;���:#*N|�8/ϼ�y�g�@W9�������*[�M�]?Q�6N/��Fވ��Q�~���'g�-��%*������R��+"X�CH�z��IXU2��xr�f{ܖ_?������m��c�בY��;D�n�"r��[���C���H���W�%�C����"�o�H�6��~�̈�	��K��M����+�)[!�%o:٘�M��^� 2>�*�!D��Q-��K�So�į��INׁ��Z���s�lH����3��O���Q�Tf.#�:��D�Q ���c�$o�)��h]�2��c��9b(�X�,����B{�a�`�T.�h�S�ܾy���X="��&�Zz|,��N���+���̝�5�iUqֆ�!�T\(�b�Ap�
��b�٤��,��ǚ���DN�O�ynEfC�@��c��@��4���d�}����%����5��E`(x�)��g.�k�(܄=f���8�ԇ������Qw|��a��X�xvg�렿D���YD���0L�؀�H��n��ۋ\�؎w�I�AE�L����*�YB7_�������7 �qQ��5sy���1��0M���W"QԂ���ט��������[~.�Ʊ��,ٮ&dx���p�b$�?,~b��g�ր+;�d6����H�U�|��=��9��̉N^���������������)��&/�~�W��j�g���H�)I�����gv�,-y�� �R�Ns7,(}s�,a�o��Y񆩩�l�?��,("F��}JL���t�N���-�$`���X��X��Ub�mS�3�f�V:E�a����/�E��c�$ �)7n�x���fE5~cL��75�B�,r�p��&%�<I��T�@�VwyZ�������K���?�m4���5��\�Z�P���靠d�rkC2Lٌ�O/Q�HR�	}�[J���$cV_�$P�*Q7�w'�%��I�{��2���&��_�� ��A#h�%��ۍ��4?�A�@7��gC_'~r,un'G"N� V��)ұ>�r���*����4�>WCih��T%WM<O����Ay�D��75x���_���4BxRl��A	_�H�N��JC)p�0v�?i�Q!'��ڪ܏Ta��,�5/�Z�@��4�N�(��i�R�d�ڲh�k�q����R��J-�ߊ�0����K�"O�ܹ	'��ݱuÝ���G���%��Bg�$E�HR�JR�:m��B������Z��Qcc��j�e���CZ4�?oѤU��U�Rb	hI��l�-ԙ�4#G�m7"?A�8��V�wd/B����wW �9�O������{l�X+�E�{ON",��#Lε��AŞ�٫kz!�Sg(}&ĕ}�u�yw�{�1-T$��x�(�^��QCkp4�uS��:k'��=��1v��i��d�!�%�;��R��2�0��9MǱ�W7�!�i�
oMf@;@�4p�a�`��bիC[T����U)~0L�y}���9d���h-2�∎�M /Le�&#R������])�Jޞ�a�Խv\A�_�n�k8p�=h�5!j|�	�����)e�]s�{��`�,Fś�5�������g��5��@Iɉw��ռy�l�R��<���mT];������^lL2�}�A��ʧ�\O8����.��;��50���H�Z�>��	b�	_?�F�g��E?�a�t�k�.�����ď���̋ �_��f_�n��eJK<5�4dϜSĎp�Cy��W��I��M={��7���i9.5�L�6����=�w /�ҋ�Йi��v��URN�ܱ���f���X�6���wĬ����?�k/���{���"T8gv��/8ĉ18_�
_� *0�R�����wM�R/���An�|oɩ��)su�!�|�{nX�!��ژCR�)�:�����;A���B�������9��o��?��6�����-���x�񧒝��o�#���&5�����kM�����@~]i��}�a����&��*��{;�"P���aQ��D�oþl7�ż�5f!L+�s�.Ic�:K"�v�/�G6I6Q�`���ڴ\E�d�y듫q*n��\V���З�ٕ�5�ݿ�<fvr�f�*�RGc�6�_��Bd}�~�!����}ni�0%�]B*[2�����b�_`�)nL٢n�����յ������ꡎG��$�"(;cA�H
}��W2c��� ��Zo�Ɣ�z� �J�����P����2a���Z��(�ٖ�0�>�^Uiqj�)gN���W�׏�ݓ�1�y�$��c���Pխ�f�������V�#%���I�kD�]�Ë����2�����Y�q�qW�R�p�j�=���|�[�~\Qm� ,ZR�<�X�>���^����d|��y�2�QaSR1a�q�ô*;���s_*)%Yɽ�E�L��i��!�x�꾪ne6 \�����4i[�3�9gۚ��*O����|;SJ�ui|�����m0(��s��7���&t���\&`o�d��AK���$�����y���zyd���(?s�(��
gp%V�ঙ���5'� �Ͷ��7h�]J_�,��Ш��L:¤T;`�F�䪠�MT\�X�K@J^��S��x�
3�k8Sv��_��Z�����G`$���P��"6U2	^����Y�:�̊L�n��bތ�����ڽ�i}Hx��yW���XGH��dӑy�X����h����Q�]���N/�U��-H�s��&����J�b/#���0</VW��L�0�,@��p�74~���]�֞)�VJ�~%�T��y4l�A���'iu�����w��C���o>��Vت3;ެ���[���W�Cfi��N�xk�LLO�&���j.�B�ѕb�J����+Pl��4Z�_�y=����@��Q?�xF=���y�C=C��/����tb�:t�'�V���!�@�E��c�3�N+.��9ցA�Z^+��p��d
���q���?4�ߌ�8E�0%'�_R�H����"Pzja���"F�ǹ:#�aIn�|� ��􆴻xQ��I�(�<�G��Αe &���p�͆�l�����}���z���>�ky#����&�Q��2��}������j��v_&8�4��2�!���.5�Q�ޛ5;M���^<L�������<�(,�`��8^�?���?�������;
n�~��A&�>����e�U $W��|���>:�N�'�L�,�k���#��L�2���k��|�Ì\��Ou��"H����G���}S �m���bsX��[����>���8�t>?�xw\F��0���E�8����,��ą��-�,B���$�+��	����2�-6�9�Ax�ߴ���M�o�O:Re/�IJRת=�(P��Kad٣B6�P�;:y�Z�y�&�6p-n�=P:f�;7��A�����R{ MեwH���-��P2���|H�;�@*~Q�Y����+Gf�{��I}3��:;�{� ˞��س�8��#�������zw� �g�E#�;紫���g����wı̾ѯ�{�55Y`�;��c��?�͉���#�eDAh�l��"����% �_-��^(�9ab��<�6̖c�bҋ��˗׋�\�/w0m88nBl�����l��rc �C2�u�� ��� <�9��~�	�^��.�U�zFRx]�j$�^0��ORԿ��QU�=��(��T�X8�o8mi;9l��y`F\�N҄6%������V:��V�#ģ.V���:D����ۘ�kd[�-�f�;@���K��n�J���U	g��p�i��-���1�%FE3J�B����~�>��m��Խ�*�P9O�D���:��͑'�)Er������$z���t��E��#��5cA�#�a>*��O�QZǵҼ�@�����U�S�%��9X{힫A��O��w��,t�n�{��]\�+k�ج�I&���'jy���RNd��x�.!o���؝K5Z2�7�^��%)�
t�2��j׈+�3���T���Q�:�3�#��Ǔ8�h�U�hw-�����ʸ;8�q��1�{5͎l��hY��v}�g�I
8�ԋd!�╇ϣ�4%#�Y���.�\�� ��D�rRS%����Q�R��%��M.R
��F�}3rpc��ҕ-��5��~�� ��^���-�B��[��yGޮ#' ]��/��t��hy_B�H��ËA��hO����Ĩ��p�	�b�,�n��� �	��r��j[[;ʇ=��O�o��?v�m@q����-V���z�#�7�U��{�
�?���B���7��jO��=xku@ҭ�O	Jׇr��2]�<�Kl�Ⳟ:�j㚇!W��"��,/�qj�G�Z;��ʑe.nւ�R�F0z_�תw&ݽLC��A�����vGy�w>ѿ�.�E<��$6r峠L��� Q��	J�q�q��Kõ~j&�#�/)썾��tx��!�_�ܼ��[�i>�Z*L���ٻ�0e$��`#v*Z�;��<��6���t��|�u
���d�7;P�?��J�̪�T+p����3�mS��eA���� irE�'p�7��v�q�3״��n{�:\��U[Z�0nW;45oȆ��6�%q0�VH�n�K�J�}���cj����~)�2u�Vo��s�͔��Y	�&T�}�^��%N{�_�(�&��OHM��W]�3GC�Jt{a�]CƝz���ٛq�Mxh�ZkQO�K���'*j&Btz��L���9�j�x,����~�HG�[��U�9�^24=ff��m��d
� ���_ �����Fe
�Čx�3vE��pmI�P
�Lk[V�KV�֎y �Oc�2�Ɠ�0ؠ��(��i���{����w�f0���~���5h�,���=��:�� ޗ�"������.{���`g΅�v�!rg�{?=����aV/�*�g�bgb_�
��ɕ�m����|�|���b؛`/���o(�Mw��z��$�[�|��Vn�%�i%���@~ȋC���jˑ�Q-��
�{�7�����]aхbyy��*W���,���-�Ku�5���@�i�+D��4��w}�n��-�]��{Z!�GuF^��� �@�_Q���L'�;k(���C�0�~�>1{;�9l��f�L�{y�����;I�-�m(z�4���i0"r=`�agԞ��Iۺӗ��i�X���VqȜ�p۳SC�Q�X�xX��bܼ
/FH��kQ�q��y
*]��)�Ǳ�`[K��T�V��ct����&&E�8B�M�zz�$>��)+��'������>�DY�4�2b6���B.~"3��G�9(����NE������d#{}��~�&b�؋��ޗ�g�[�N6��>^��y�\6˪gY�/O�J�w�@BH{����0�#Ҋ�V��p�H��g�:�����d�8bއ�~/�T�^B,<Q�GTV���zO�0@����0�����G ��H���m%�Y�|�F���E���e�Pd�]3�H4������`%�p��wO�C�P���9�.��;���"/6ٶ��V�Mݘ_� ��cI�@�Ո
��-%��Vk���;���陻�iA�YK#L�������޿��G�ԇ��~��k��,��� ��ʖ��R�s����Tͅ�moJ�hi���Q�[�����ֿ�Pi;e�U����@1!h���@�_����(�Fz�E��������"�ل�?�d�����i�i���7�p�L��=M�d�@_p&�MF6�3�Y��/�M��?�MFB[7~���u���`���	b���ա�a������޶�YեR9z�i�0�����v�g�G�����Ї��4^�:�p%7e5&9������L�sYF�������J�\B�c�FC#|T��_�i}�r9rمD�AMP�J�M�B�2b�������y�zc���kc{��'�zU/jq��c��詚/Ș���2�����
���x�#��d���]�]�OH1�z�}�6��o�En;z�8����U;zNsv���#V��דs�-Q������Cumd_�x�Z	�R��\�ǋ�F)�|�^�B����>E;g 7ɰ�ػ�z�R&���{�;������g��n������H��>���"Ͱ/�x@���/�9��^����@"
�����5WG�(�(DI���a�ڎ�pz��DQ.��|�3�p�����×��F�3��}���Y,�<���(� �k�.}�!��fO:���R�@����8O��i/�,�̆��� ��������*��Tѝ���N��ߩ��Z��dW�Ys�@�( �wڵ��,k��Bʱ,߈�QS�������l���z���poS�W��V��<�ss�z&�^4�&�a���ۙl�`E�%�+��U��̏IƉCZi�b���q?a%	���sc�&��B�8A�VB�ג�h�#��a)INo0���N@;�9T� ��T���UnA��K6q�$�a:ٜ����fǮP��$�a$^���\Z[��ڏ"���K��_]��8��:J��-u�L�^���O�	C��\#��Ac�lT�;89���%����v� �x׍�B�� $F�_�$Za�ծ���լn��,6�����ݭ�* �E'yO��ډ���VF��JaI��"��q���s�����Z��fv�/�������ќ��(�r���8D+��)�æ����j����c�A�i|{>�[[EԮ�)ob��uR�HU�SI��,�p���������-O֘�����i�'���6�;��H�Ye�<rY1�:�֠�N��b_�41���[kp���v|�k:�9Po�Ձ]�A?YQ �V���l�3*�)�OJV�QB%�X}�+OxEA#���`p�M.��� _To�g&\Jֈ��{��4'`P\C!�;�B�H�ay��a��O}C*6̋:YT7�0	o07�u�٨U1d��K|xn˷4�lܞǢ4���ŵ:^�e#����A���nW���+�a�@�%B���5wz��������� _*��~���E���J���a����Xy�ƛ�A��*s���=95|��J�Q|���4�f5����)J�9���&��{�'% ��m	o�1�G��e�J���p�x Tّ$/t� �u�p�҈i��~Ϩ�5�S�����Y���i̸��k(Oڈ�8~Ϡ���GqQFd�<�v�J�����~Ճ����Y�v��ob�R�LR�?}R����P9BJ�Os��V��|/E�*'��/����6���E�o|�w.��Q��M�F�:��ws�W����n�6���G�w��v�WL*ȣ���i栍b����"_=�Ht���,�4�n������Bk�Cq(P��Lʂ�6A� Ia,5��_V�2?��wW7L��tdhv�}�Q��;�-�8��-���l�6���>�_Lo(�}�X�խ	fg�ɗX^����1uW�2S�?���2�^a~3�&�N��~Me���tH@J������\@����+i�|��~D�ɪ����iSd]�4�Eݴ�)eE.,BO�ω�u�3<&����z:��&6��9w�0OR�۔ԭ̣묏�SZK��LMM&��!����+Y;2t�f.��*r��Y.��Rɚ�@G�X�^���B�k���R����P���A����9�[��7�n���C�n9�h�\��:-3 G���:yw^9
T.;�vT��T39��xՋ�gcX=��b%��Ď[�B"8�|��T}���D/ȣ���7�����]Q�"1t��[��$�8f_y��c����G0˛�j7-\���<��`����t+Ɗ���R�D#C(����`�"��D����0���&&�oD�s��;x��GAsY���?O�i�^ c�,�5�g�����,󆪄p�s����,մ�ֵ��wI��lwG�4�kR�{o+Au��t��@~,��_��^�k{n�}��k���(���G�}��A����5Zt��vv�i6�mY����@�ȣ!!�:�L��ۓ�۝�I��n�<�=7i�AQ,�?t��(��R��Lؚ:r@��1��e���ũ�p� � vS��!�'���J`�^W����}�@ @%l�(O#��?)a;�D�������
n\|�ͣ&�G1�d܊��?��d��B��������{[Mu#%��T��
��Y |�/�D0��o���5N���W��H#���E��#�`��n�U+��)�*�:�&-��iˡ8�b�Bi��K�x��/���Μ�:������y���d��\a S���g�V��eBZ>��~�����~�`msS�,S��l^����t��<CaJe��»��Ӱi�]���寢V駧�ʭ{P	�!�z1y *��t��y���EK��)��p��N���.���8X�NM7�KE��rV�l�ij��x)�t��ו��"���Pk�T�<�o����q���~��A�*��+���ՠ�sN���C|�q��C�@P ��:m�jӟ�}]D��z��P��)|?YW�n�:�=��=][���m*k�Pr�/�⒌bn�J�:7O�l��O�"�	2G2�V�7؊���G��6���RK]��Y��g{N̾Po���9r2o�NMmirY�z�)���a߬��}����[�P�����~���M����JeA����#G�O������C��?��~�<�B�^J�&�td$d{+���~O����@"Υ����F�&
	^�а����� ������`lx4r�K����[��R��P�������.���	/Yx*ϭ_]Z8qI�>�h0@��~���Z4׬��P�Z*F�J|D���a�Yt@A�sb��Z��uuO���L;[zT�W�s �zP��@&wv�-*��b���) ��`�|$���]�EHw3�^R��D?���XFE"3)[��+Dݭ{�"�Sw��z��\]�6vW�/�1�ۅ�-g y���p]����M� ����l����f��4�R�N�o\��8+8�Y�Ҩ��>���h��@5Fy8h�Zwe��W��`��7�i�!�K�?-��pD�)!��9|v�k�|�J�~�hwo����3��ۺj�Njd=�娪�c�G���g�[wӢZ�55k|5� rVٕ\h�����_����8g��S�3<::���'�s*g�23�+���05S�.�n��^W����~>�:u���Jm�W�`�u��Y�eLh��ϣ��-"�N��:��k��`]��x��o�ĳɬ�6����h~z!�V�)���)�T��NX�b���%'<q����uOO'��^S�*�0�gP�|�����f�*/X���)=_8~U��~�P�?D�,0�\��F��1�2W0[M2xv���$:p�7��g��.�g����q�_�ULFL	�/F0�hlƭD����'���=�Hs-u���`�ʒ]�eQ^1���?\5��ٝQ.���{����9׍��h���B�%���/!�e�9�GN���R?����t��y�gIw��g��-T�2�n���E�UF�*�ؘ���JU�g�E�-�-AG��J��=\�쓩�������@YBP��=[j���[�{$Hp0�L����j����2H��) M�Z)X����ڟ����>#�?�EJ�qK���𱩾-���@I�H���ߛ��s��ᴌBM��u�ۡ�p���H<1yAh��@�:�O�����I����C�Sq��v�N���ѹ�1���yש����R�Nx��6d�����ɺ@b��~���ԯ�O\3j����}��L[�'�2�^&?�rq����í\�66����B����4b|r�Z9:���gM�1ެ�cC��"���띹�O+�p`޼���'K��H��;��8��O��]�sM���cxv�LqD�Ơr�-�	�'GS�_J����Z�(#�X�q�s�Q�����p-1��7�і#L�<sejE�Q�-P�4��m�W�~�+6��X���1����Q�S��P�������5
�5ΟV��^3]�^-�J�J��zT�����4-���� �gnj�13�+�܄�[ʶp���8����	��3�. ~�(��
�PY�n���{o�؍+�ז֧�^T{�>��%T�T���G���ފ�<`+�[��2A��{��|�;b�OW
�MT���+���}A}tfb: ���t"�;�9�g�-�������=�,2b��/d3�ٽ�� l�e�2d|o�|��Xͬy��/O�r�U��>�_�̌�/��'���䪎/y#N�~8��l&)vN���Lą��c콆 �m�X1�v� ���W2�e^&n�lI	J�0+mi��Ȫ����P�!1!��y�C��쟴貘�#^��T��0Ȭ2��R�U��"�i���0��-<#�N��c�N� UnT;���-Y��G>lԍ0�������P��GÅ9���A�4'ٙp1�u�n�&�_Dn��RYAG_@�xǶ��Յ��׶�s�+��U_��с��������Pȡ�����L�`��=��ބ���@	݋�Y=�!�]�ݸ���	�k{���z'�W ���.�v\�|Gb��ݰJ1%�Q���'��K�P绍�;av1� �x��m�z�yfEGu��|��>�ZD�Х��=����
��tL�i2P���"Yh�"���3��d݋���_���P�ħ�4�G�$�zv���Ȱ{L���.zۦ�i��� ���!j�T:	Q2�7 �o
�G��	Z������3�����,�TY��|�!��JTZ�v�/����\�����{�H ��6�@$׎l�,|�F%�׽�tHj"F�n�󉋲���V��<���ʦ���ǎ��;��2��Vt��(ed:V{>�ڛ��e��^�@��%?pƍ��_n���v��Izw�%2��s=�MQ�ܡ}���l|<���p�7��R���)�ܯM|�<E�_���a,��G�(������`���D⺼D�:�;��y�����dY�S�p�Up�$�f2iN{b�#ു�1lB��d�)��	��F�Ȱ=U��=ys'MmvAפ��vLA<EQbB�dy���o��5RZ���M��{�����f�p�ҩ��j�'b�� �o
I�wA������n��� "���}DM�j@�%
LT.�=ߙ�QՌ>т����>jM*q�w/��i��3�4G���*�8��v��&��_�#(q���^������.����nP�eݳ�M��(�Y�q/��+��l���W�lq`l�U����vrE-��ql�ϵ�^�B�\�Z�2�8�FJ��>d]5�t�q��KT-o~m�4����\z��@�?axmxrB��E���?�5*�b��5NR�D�WT��b�զ��/N�'	Nl	*���L#�ή�*gFz)��w�_�0��(�����C'"��R3�I��q����>���L�5�9�K+{Ks������+X�i����]_p�axv�L��襱2�3`ʄ�k0�p���á��@�X��:���}`2��}�������1%,a�W��)0�F����C������Yh�	�5F�YB�
�ÄE�B���P
£y��?�K�
o/+�������$p�G��Zz��F?!J�A+m�4�A�tQz�o�<7���ШL��Ƒ��r� $��
�z��X�� ߼n��V�]I��8�/Ϳ4��G�\P+�$�8����$�7�U}*1O?�=��ג������
ˀ9�����`�$0���/WfT 5�U	��"��oJ�����[���@)v���_L�z�m�8"�UX'���Q��o���;�2�]�X����kJݕ5)uu�0�sp�f�vk�$웽�\�7�g�x<7�{�C}�~�`C��bd��Թ�lH� ��Z;���?���m���>=��~pښP�	�r^���z���#3�g1��a�s�x���/o�^��gQ�ʡ�#��Q�*���!L6[��tD6�e�^?y��{��֬I��D��3L~r5���&�;����g�J���-W���UqO������C�)Ab�|L�g��}�[  Eut���D쯳g�[8��v�����ۙB�m[�8\6��#�T���8�3�Ũ��|�=N��**|��b��X��ќ�������h /^�h�c˄A]�J�Rv)羅�*k�α'F��︀;�2?4��>�@F��I0��/*�\�Rk��IO�Cc�bi��Et��~
��!m�lp�a�_魐0�㙌�yY��4<�_���.�NX+��G��[Q̄\|�m�O�z���W�/�P-�
A/�a#��cNL�e�@Q9+�xn8S^�	�ND�JYE2v6o/����U�5w��)�߳�Z,��'���!p{�J$L��)���U�`T~�=�2j�.W�@�IMLgR��	Z��I�f��ڬM�����
�H�Iy*���Q�uT7�$���97&�O����N�PI7G
�k"�|�o�&�$�>#b������R}���֙vz1����*e�'W�݊���䆗9��]~g����a&�r��g��oh�JR�t1p��=X��IV��P���M������k?,�}�ܝ�T�{�*��8��B��OEW�Mo�~����a�t�r�ը9!��e\A����ו��LE��A%�kM�d��B��K����B������a�X��$)�-1�P���,P��4�'׷g̹8��Lw�L�?��K�1iќ���;;��(�]<d���mom;���8�<���B��0n���}(#���yL�Nre7ڛF0ɦ.�����@i\�e�P���d'�}��>=��k����n !�`���L���_R�p�̾���2�ث��F���Ӑo���悻�u�?�-�RD�����7b1��!O�X-_�	��(s�X9�8��߮���Ӛ���R�w{z'݉pDi�E�V���{�c�S�~�3�*RY#*����~;_���ۍ�;�	��c�ov\�7��+r�W���V��w�'`+�K�I]�X�v�GQ �M�~�����7}#*�IR;���)/o_�J�����T�au�_2�����S2��λ7���#�$���U�\mBFl��ue]#s;t�X���\�>Q9����jy$�W�:�uU��l�ռ�z� ���!�+{���D3C&J�����!�c��s���v�|��c��.3�.u�ݏG��&��������Q��C;v4� ���G�o[1spnޟ�XA������Ѝg;�8��Ύ�9�zN���v7��ggr�o�P�D�R��v�D���V�w���+4�1Bk�
[p �.G벊2CÐ�~�r��$���14����<�����{A�l�d�aȬ�;1i���Ҭ<�G���-�Ϛ�������QB�ʱ'�T]ܧ�D���Y�d���
�W�ԅ/�#���X��#���Kx����0����QTan�l���]CR~0G�w�p�Y��e������^��߼Q�����%<�Bg[WhM&��Ǳ�!G/"�ɻT�x��FQ��#������"������&�K]�Sn5��6�FXO-��)�{�b���� x�,}�W��R��F1���e+��i�h'˕�?x^��r�(����'[�s	(=�ٶ��O
x<���n�+ ��A��9�7&m>�����M5s�C���d̶5#�P����\�p��Yhݶ�t��ʤh��{�p�[�ɋ�D��6p�ӽ�Y�ꕶ�,d����3aw�^�ňɿֆ�]T����+��׋k�.����ZF+g=i��i�Qd���^�X�E &l]KT|���L���<��)��p��}Q;���&oo>e���{r��3��& ��J�Ӭ��Q`��?<�E�P]"��ۮ�u�	��d���ŷre�B�i�ʣ�v���D�=G�\^�M��Q3�������#���V�q͹��;s���d�eW�"��olL���3ZM��j�2NzWH)�������eq���?���ذ.��X��Y��N��МF�"ٱ�td�td�����rk`�Q�}��W���h���D�2^ڒ����;�k�J�����>>Hd�@9��Wx��g6�>�5mlM�.���Wοv��l1�DE0��΢��6��?u1̊j�j3^/*r7�� e3�����k\wp��~����DId��N����pH^�/����,|�7�B7�E���X	��d�H�uO�y��7��/	�	�
��c�|�C��P� ˽`�F�	�	��Jy@Q�q�x��V�jB�ޱ`'���������/	���a�m�u�뎢񓩤e�I�B���]������F�E5_N�\�D�D�S���J$!nQ�,��&�Q�a�����N	�e9zJ�1Æ����o֞��)(j�Һܤv�y��k����Yf_�ut*XW�c�"��w�,t�&��"6Fg��$_2���u����P*T��t�z�L?�9�D�hX�֙G���(�+�N3.G5?��`ؑ!pbC��C"N"�kTp G��f�)�����4�9M��ٻ�U-��t%�C��qD��� ���A왖/��� �}�nM��s����zL1�&����IP��?��^��+���F61�A�-rk��]q��\x�����z�%�#5\�A1��[�TǐJ�zcJR�)����ї�&�b`�C�N�kЭ�2*&dq��Oj�ڎ���{i�����V!Z���JE+�e���Gmx���R�H���W:E��FÆ��������[˳Rz��/I^�6����#WJ���k�*Xz"4T�+�DIL���"xv&�5��1n�m�6uD���p�RQG� �� ��q�VÝ)O�u#֤-��[e��ԂXl�He�ڊO��}R�ǆLCHh�W���g���u��9����쉉�u��~-��]P�_��rU,x͌�2�A2/���"v�n��� �#(��i	V%N���l�&�&l<&ɏ0�6\� .`�#����>�6m�*��zˀ�>~��>�sZ�:��$L�#��$�!�ë˲�G�h���L�GCB��XL�3�p��E���@�}�2��JMu)�,&.�����J���eݷ����?����ˈ>��}=q�:�s��gR�<J.и�m´檽z�6� ��jΉY�`ӏ��w�3/�������o�¾ս�M�7K���ퟅ�D�h�K@�I �%��!�$Hk震�0��h��uD&<rv_SD@8ܕfW麇'�٭�g��� t ˴��a��@��8���J���O)���+��o�(���&r�p�;ysd�A��5�a�5���L���<�oW����L��!�r���l�`b���|)�0�������(��/z�h;ѹ�k�n�ń��T�z/���,�� @m�h�qy��.-{0�^�YKҗ�⯖�>4�A��g���*��Nxr����Oe�����l�Á�ܷ���9)L��d��;��_T�	�`w��L�hGC�O�Q4�K�#*,\����cd�ci!t��)��?�7�R:��Ib��Tw~��S�	�sQ������1����hs���l� �S��ʳ����N]�,ZE�:��zT2�^��m>����p�dW�2��\E�l
Qg�3��r���Q����	��Q���AU��n�Y�y�8NP;X�/�=Bm@KU/�r�J�I��`p��#�@,Ay�Ń���v�NR��0�U�N��0M��yN_/�g����g_�ΝS�)�;�3p�d؛f�]=+	�殽p�3�m=�[ŷK1sVƤ3*lL#&C�d�Ln?ᦏ:(��A,7�$�&�?m��٤������8��U۩���q~'�䘞����ǡtZ�Gۗ�+NS�t+��u?V��		�|���5ӢB��+�d�m>��U�El� Ɣ����K%	�W�Û�C�
ྮ�#�W�T�Ϳ@x� tG��0;�,�k;rU��}s'@�~��f��?`}#��C�w�//���m�����
�[H�B،uK���Z�l��]#=�,���:(���uswX�Ⳅ�q���(P�!y�@?D�h�`�(�U����'M�q��W�`ڛ>��g_�2t�%<+3&pC����DP���y���[���ϟ9;�7�}j�Ah?�h���V�ҳ|�:�
�	�R�5��k?P����}���j�Z��< �M��D8iS�ܰZ86��t�T�N��a9}���i��~ڻ��WS��X�V?^N0l͢+� @{��r�Yuh�R�rBF��gc���0SL��劖=��^/ X�B�^�x��?o�7��T��C�{��U���MGO�5q4�!���Ez^l˱cŹ�$���u�����k��2����e����ޑ�L:Q�4�>���3�ҹ�^�KR��,0�Բ&h��ĝ �9��FAO��J��Z\�5P�>��}�U��w��L�ǊZ�*��S��'���ˠ{��ݪ�a�O@���i�L���Ru���o�6�{)��[-;y5�̗�(��e@��]��n��!Ԣ�ym��~]�H>�ٟߨ�i(kX����G[�wT��k�Mw�;K6����ӍEΞ��4�-��z ���l1����$bO>�(�������G���W_7U�ll8��/O#q���}}RĴ�v9]���� ;At�t� �2�����G�/U#3\�sd.����&<w�4R�v���S��o�.�6��P;�i.h/4��?����~3`��W$������G*
 ��H ˪+G��$~��n�Y}��͌�� W��l�w#�V�W����J}��<�:�XSA�w����V�?*�96����&AWI�E����(\B�|�� {s�u��?�IA�*NQ%�In����� qN(�_%1����iis��B��§�ϸ�k/�A�XN���ŉ���Ŵ�����A�O'(��"AՄt�;WJ`x�\Z���M�+��fP��ox,Z���~�5�W����8.b�g�<Ⱦ���f�w�=�;a�mYN�Z��߽��՘��ϭ��#]��-$�C�t���0�G�Z�w���S�*A��!W�V���)k-�:����da�o�I�5�̷wAa,��9I�?���8����p��H�ͺ@64Cd	
y�r��Ɛ������������Jme8ʾ������D,EX�����i��j	������	��b=yQgQX�w�ݞG�Nh��͓���u�]�5��*��Z��Ǖ
�W^�N��A���FW��1���[?7ӓ��JI�̴:J�O�B�$�B�����a(�2�<��I.!Ε\�^�]��l )9;_�����hX�+E�b lz��˼pP,�o���ȼ��Ѯ?^�w�J%�l�$��P|�P�g�x�뤷�=���8�{���	��W�ZEz��
���Ħ;s��ςeD�N�/��Uf|�'u������	X��u9��n�X����e�p���f!��v-�X���$��L/�I���������J�b��3���iz��9�1{�*]b��ȝ����p�ŚW�v�1������薆*���r���.zf�	2��kFȂ���������a#՗�K����)fm��������2W�u��i�PA�Wxn7���d��N�Ǧf��8AԳ�Z�8d)ƞT�6� u4�E���nr�%l�Q�;�6D����<��|��L�nS���+ �v�QD�B�a�7� �iGF�z��a*:�MS�,R��:k�KvX;AK��{�.Yy�S6"]K�]����Fl�6?B���&P�q4�'�Fvz��W��e!��9>	Z������>����ʨՉ���w�C���r~��0e[����.g�|Դy�
����\5���g�Cz�����7 ���w����O{�nO�!cZ�-L�<1�5iA�X���XPSd_��9L����Ίti =�d��15�{�7;i��R�W[X��vQ���KX������)'v�-}�=a,�-RM#�����P��q��g�4!7�S6�������؝Vk��@5W~U[�C`��Dc��{��plS��
m���)JRDI=y�
��;�nk�ә!�Te4�����.b
��f�?d�DC��l]u��8l7?sJ�X��G�)p��Q������aH�(J�X������q����U�8**æ����jh�9�a�N3̣O�t���<5�y��*�$���Qx��=�5�W3�G�5�B�w1x�K3/;�<��'�G��x���7[L�Q��#��)�O(H���l���Vة��Φ������d���fk�$���,�Xp����]8*�QɺJ '�jV�����go�>����ߢ'��] �_;)i��)p�Ve&*0�U��&-��/�q^��xw��v]HZ2���9'���߆�����n����Ţ�y8,S��G���r���$&g��S�>�3q�[�Q���%����J����m��56�h0R��ru�exu���	���x�B���ҽ^�wX~��3�K�
���@�~/*���U�Kަlɬ&{��� ��#��L�lv-*\������?]`d,m?䮔���ıp�[�p4������9�Um
��Z��-;�lcQ�q�)�#��	�~o6r�;��C;�c��e�Y�|�Z�g�e�:ؙ�� �'����<���hy\�R���~�c��S#�ʦ����)��ԔXG����A�j�["0���z��.� �2��j8�ʑ54*���N� ���0�ϲh[�(4�[�F���K���i@$� �EĤ.Yo����<���_V�hYK����A�}�\� ��!#[#*�T3=��s?��l�N���N]N3�"eyğj�J�U�~�k����<���V�>%�����}��`�bG"�H&���Mw	Ӳ��ּ���իH������b��#h�p,���U��^�@���^2%az�;ƌ�єB��@v��g͞�N�v��W�04@׈�j�Yyg#B�Z��%1���\��W�n�NY���U�p)Ϭ��/�]9o�w�1S��J��t}J8��;ic��|�P��
�w�]i����^09j����l��F˴Dh�h��� ����=�9qm#ͣ����M�x�ĤO����]~?`�������A��fQ	3u�
}�6��qQ����톴�����3@��)�/@*s�V"�P�>:�@�+4M���̓
T�u
��;�ӷ\�A�be#�Cevl���j:2n�w��8�P1�/F_E-jn��Jp���0:7�<1�Cց�ʰ�����O�\sr���2[˸�����X���;�����m1�{�K�oTYc1	�= ot�{Q�ݹ�����rrW�/��Q3<EoAu�氽Q��&|�E��sO�v mn�P>Wq��N(�Y�@��lMi�����س�	�@�r�Pgu�:�9�v��*9��?#m�@r��4�_,d��~�.�o��ff��9l���Z��� �}�2��ֲ����"�~T�Y�����V]̡s��Yz.0S@&N��Ns|B<ͧ����N�}Dpl*���B�L�ecZ�=&�v�^���Lls���F�JA'��N��)���V�E����V�ee�LroZ��{��M�_��Ua"�Cڹ�iG��h�p`T�ȶ�>x���ak7y����!�Ѷ�������Z�^��`������dn�	��	V��:2�2;��}�|�Yv����*�p%x)t�:�IڈLZ����cb�7@��R�.�)�m��W�RG6�_ ��A�>��Ȕ��������8���)а`��^!�6=%s����0u�zvwT�Y|z�G3�
��q���xĭ�t��dm�ĥ(⺃le_�������r�ڨf�i�iհq�Z2�]J]�����Q/ ,s�~3&��󘗷o�jT'�L�8�����#A�{,p�����# }�+�h�o�igWk7l�/���,�#�@�zO;#�և��AY��Ҹ��*����PY����O��>�@9Эg����R~&�@�ݾ)�?�R�lyk���f������p�]�,�u���6���L� ����:�?ϊ�s�D��GS�����WH��F��P��s�q�/���5�p-�s'��$%0q[����q'#��ԯ��������E��X��8�lQ�����H��j�-D�|��~�L�X��`�	<�L�om%�I�#,� 0R /ê�&4
k@�qr�`LC>['��Za�է���ـ�����o��n!w���������.|�>�RҔ!<�����յu
���篨��~�=���rƍY��Vf�-]Ǻ�����x�)��2�Ƅ��p�����Q*���h�Ω����em�.���܋j�� �%"���a������cR{��ʻ΄ �̳��,,� q#���"�d���$�sWia]�YO��� %a׵��hv䡅��9v��0����o@c����4�w'����S���á@�m�qM�	��N�,8)�j��&�#��n�T�.�Dmꍨ {J@O�وW#�Y�qQ�n�[�u<v�G#x���ԞуK�&`�4� Th�ǒ7����>�wU2��x��<K�p}����G�U�Xcu� 8O��КDq�Ox���*�{ ��,(źTQM0�=�`^|�Y�{�z��9y0Ŋ{�߅^T�_��ͯdC%#�g�4e{f?��$ʣ��g��sݫcJ���$&��K�T婐!��}�Ds�K2���l�+kP���D�Q���t5	8�;�Y���SSk�V�@���0�ox���3��]�+��)4�:�i���oZ���S7tS��V�f�.�7�ʴ}��A���<�%�!j�x��F;�fVB�+W:�
:���lk �l�P�����˂7g�q�0���-bN���[��b8}x(�EHs��1	�����`D�D(������4��f^�� o��Ƶ8bO�wN�3"����r�$���J�#v�e�\ϙW8׎�u���}M��<j���~��#4ž���_�)3=�r�1����)�E �����x�-�$C��k�d����񏀚G
n-7�����W���UO�v���U���X��4���+�$�M��P��]/ijh�u�8��dpC�ֵFt�D��]5��Age���s3y���:�J�'���j��Т�qѠ<G�����~�5?
�FXA����h�P�{�ԑL7ּr$��8}'S�@,���="<�볬3v����!Xg���o0)m���C��Oq�4'��D3ݐ�0`������ڌ'c�g�\��F��z�m?���͡��x��c�mYq��*E��
�"_�.�)d���{�o����Y�A���1���x�yaq4��ح?rvfڽ�%��s��S_kR
�7�g���Ӻ���r��2�T�:Q�DX=)�-�SL+,��`���}�=�%)����H�@xdRxvE�3,8��:��P�-�NvukG�Hޙ�A_�"k6L}���<�Ɵ��Q�^.7ȴ���{M���	!}��D6������s�N`ltȭJ`�7S�����̍+n��"��ܐ�L��$�X����y���D���n��}���ͨ�ۦ*����y"@ֆЏ�( ���	�~\��w�hc��k���F�a�eU�֊�Ӭ�"0�/��I������ A��3�� ��abK���d�o$M��]Dm[���4"@��3@�f�$_B�_���n��#��Ur�u�BU�W����`�%��%^�!��F��{�=�(�ē���I�N�yK�(�]�Fm׈��%	�#ڢ����Ɇ+Ů0J�G$S?Ty�M��- �%��ʚ��Y�%�u��O��n�����|6Ɛθ�R"S��[1��g4Rp��m:NǫL�Nl�Y־L� ��}�w����gW,N�^x54�f�D�ϰ%�Tُ�����-|�\}�[��(4�K��$O�(�����\G��%K����܅��j����\� ���t{�r�_!���1x|*�	�	��6�qT��(I��z�AK��S ��ͺ(`�����$­�Y� �������6��9�8:��}g� !IPF�5�C⒓' �j!�|�)澠Ћ>��Ug�����O�{ �mK�9Rb��8-�����?�sj�X�ߌ�ܡ�8����Nm�Z�c�V"��Ξ	ȸ�N{#��fg�/w�Kݍ��^�D���<ǘ�S�/�)��U4��֦�����Y�$Cj��H��RZ�k��v�-�t%�^Z�k@|N|��m�a-4�%9(Ax�8/ڲA����D1u�1
��M:`V�j�<�gG�:�6�;Xdލ�3nX��	h�����OЂ��`74��|@C� /qUf��5���'4٠S���kʰ!PX���m����a���C�P�ځ����@1a{=�-�X{��A�ҁ�#���A�|}ѽ����s�5�&j��[��
ܭ���xF5Y���iC��Aݢk�J�&�Z�v�^�c1�i�����\N�0��6'�
���Jxm�պE���ֱ�y
S�tc�`;�`_�H
����;諬v��R�;dNK�5QP��� h�?�35�4�ʈ�D�p�0QHV7yh�'/M�<����?':둓+`�,S:�v�i!+���ٹΠƃfDK YZ�^�5��FJ���me8*F���e�ەG������6�����1���YO:�U��+:��8�^�%i����=�H��D5�O%oN���D���4���8F����N�POy���p(�&`�f�E|�Q���Z��]j=�=Iwr>���zyat`��O@��bH������Ҝ�Ǟ�me �C���r_�����=X�1�m0��~�'.�#���i2�l�?a��~��H}]�TA�{{��a���f)C�`���YgD�9(fŃI�˺�s��+v��d�<#�=ٱït���eZ׿�bN�u����!�\���J�z���nKsI�[���>�G�WB�#�}�������w�f�ƾ(k@$6=���֨���8�3��=�+��YN�M!�G$�v "��O�,ML�Z��[��_�\5
�����5��=�Z��C�I��>q�y�^[��G)�D��3�����X�H�}��7�~!*<���V�)�Ս�Hm���$$���\G�c,d���|�v=r�����,�g�V��v��]��9�l9��Q��:�(K����B��E%v��-
Q� ��1Q�������:�E�� �H��umG�ZPA�Gl�^�p��m�&k����m�![=�q������h����
}c���.���樭U����T�j�.Q����8]����l�����l܍B�F�̓Rj@�����;&�Iu٭�(yҿ)����.E�$o���~6�D��	��R�zE��F<�����˵�?K1#Q=��ݼӤ�U��*|*ۄ�vz�-��w�m���7��iZk�n��~yj�~�\`z�I,�#�($��i�r#b��ܿ�;� ��\��+�T}I�R8��	1�e��pq����VG��%tQ�FV3�ina}�v|80h��yU`�=�Z�J˅�O��JkY��X�x�a�y�뉖�ĳ#j&8�4B��>S����H��ohG����m�WT{����ռ�~-����ԧ��vǪ����˵h=�吏B0����I��zҗ5�[��gȰ�R oպK=�lx6��t�O�be;؝%�8B���H=ne�
ͤ&�WNr7����E#�Cn�!m?���L[�R�Q�u�uH�4%?f�����^�h_�꣚�k���� `2S�f�m�è��+�YĢ�$'s@�>��U��&����)�P�K�z�4K��`Mt4o�M��n�N���69r�%�|)�������퇭�MHI�;j��/�v'� �i��jj؈�߅ �����`%"�5%/��ɟ-k��-��Ѝ�y���n���W�X�\x���Lnr�|�J�o��K4bƩp^l5qc�"�	F�|��&,��o���Q�f��.e���?�F�����S��a4���_drO?o��D�/�gj�KZ����-��)6��Xz���e�;F��<c��m�Ԅ�Q�`����� w�G�6%0ί��c�T�??k¸�����.��u2#�������,�a���)���~0�φL�/���-k*^1FM����)1�4z�Ǻ���!����9�1@*:�B�V6~�ev�@�K��a"� �	#�S�r�(�+ݲ�Ʃn� 7|�~�8���5K�}/@AF�8� >I�BDc5ϥzݡy{���4�mX�\��f؇�+������u0�� ����e���	贳�S6��r�k��"��U��r���Z|�=�Z�#��+��a�P� �A�ߗ{*�=|��gF�g���8�:��Ք�K�휽�����m�]����^M�!3v6J�8�c�K\f16���y4bXЌ��yK������D?1[Վ���ꡑ+=�Z��c�t1�"EX�I��������XHbcZ�İ�R��|M�7w6��ALmbm�`"��g8�#I���q�%�������0�����R%�,���%�z81�-��$[1M0,i,;�\�d>jJ�+ܑ�ɡ��u��D�&�Yr��y�Dq���7�PO\ݎ�,�z�?U��Ȓ�%�<�|d����ȕ�&�exs�B��&����L�qf_���k�`��j�+~[�7�|��N��sZP�/���]��q�Rk2d Ʋ���1\���rf��+|�J�e�2�i'n�3ٺ��z-84���yk>��4'�����mo�Jo�+k����"C���X����(�v�.�J��8,�
<��m�yt|bTյZ�5�(O���Q�^զ����"ə*�T�C�9\k�&�*<hD	ug؊�䫞���> ������587�M���ݤ�+�*�o,��#ɉUϭ]q���~kR�o�d��}W�����6���_���D�η���l���N�t�0Q������$�*����ʺ��ھ���i����ڌM�F����sR��`��+�	HWxh�2pn��~����v�Ԃֶ�� �w�/��^�G���M]!�ձ�Ή�4aU3�F6[����hs�RԼ"]�7N.��p��q�W�.�4��L3W�o�#�������¡��+��o�>f����+���A=�3��i��\,m�]NG��M}�x*��Cw�0xwGn��8Df��'e�[w'�Mi��R1�k`�`�&p�]��8a�+���b*�`���&��4���^�Zӂ@�GU\O����%������ ��66	������Tb�6�(�_0g�~����b�2��&k�mSl�y�B��O3��Dj�2=_�����*��=�M�e[�?a�zɣG�h��3��t�����<&���x�@
�#��%+nd�ʖ�4�0B�ùLn�V�Ե��T��~�Oٺ�8�=J=Z�4y�s��
���B��)u{���~�$����CG	�M<�W���0�T��d�m#V�'$���QuP������	�F"�����\��r]��IU���;��q~t/��#��]�s#�����c�6�˔!�
[�	6y�j����"r[����9gl8��r)M�����	%g�L{�U+IE�vk�%Ѳ��D@�.�P��#O۞�_�2]�	��Jy+������$g�>�W��i[��7ɫ:l�%�n9S��cd	;N��S`�s�A�pf6�
�%�񚜽h��<��ݥ3���rR>���I37t\�A�7�VY�뾔y��z?�T�&�%t����pnY�=�zm����y=��~�򓿀 l۟��2���`�<-^}7��!?��m33�-~Ʌ�\qU��r?�ɑgX�0梛�1?ӭ���.y3���s~�g��g��cޗ��,	�-�t^ߍN������ݝ�������e�U{�Q#>뒥���\�]I6�GSx�e�9EK�@L��[r�7�qJ��h����Dתi�����v���g�-u���0C&����|�I)@!.C�.񛺺��n�� !A�H�6���S[%��`��D��_�v���_�<+�>[�Pw]��h�^�B��Γ�i��L�N�c/��f��_��4�f.O��g�f>r(���zA5�*�Ϲ������e����[�,@c�ܥ���]wAj����F���ϡ�7Չ^��kbbN�����������t���h�܋y�wU�a�>�F9�
~�R!�z8�϶��;i���e]�Z��lT�ٷ�;[�t�z����,��a��\x���(PEߔ����\T�:Մ��Y+�^�p/Ԙ�;���װ�kr���ؼ.��_=h��/_���	ׅ2�yaATw~�
aW��2&�m�¢�g�a4K7lM�H.3�|w[�)r�L�-)�]	?�%M�b��n���	��F��R���u�z�ʐ���C�t\UJr�K�/��:�^	>#�c����d��P�U�''pW�Ϲ���`/�4	W	n=�KZ<T�euq��CI�����!f��^��)�k���7�'���K�9�̽����d�YD2$��:3+�P�30hA9��J8t�3i����.{�r�],��f ���B_�6\��"�LA\Z����l�����hǮG��������b/q�1����PI��h���}��a��Z���E1F�Y�+#�F<3�Z�آR�Gp�P���#ׇNX�Ӫ/�a�
��%8���z�,�, � q�f��R6f���l�X�S��Xl0�d��/��ZQ4K��UԌ�1!~�5��,.��JZ��;�	��<d��iϸ�N	�[G��Ul�U�F��F3�1�sI�i=n��	_���1��,8^�C<Iϕ ����2�&[��0��`q���c���E'0�4�b[�È��/�D"��c1�G��"�y��b�S5�>�"�]�ؚC?�����f|e����hRYgʯ�<��W�nT��$ړN�iq��pҀ�[W3���#��'ŶW8��je�?ĺ��;M���&N�A�>m�ǉ3Z��ƕ�LzzϮ:Iau60�(�Q�m_O-ɥ�<�����١J�D���|�(��+)���x/��f��U䏂KwGc�~Tb��V�������bG0\uO����8��MǞ��g��Q�"�Ŵ��mN�z�>X+&�9¿��l��&��d1�(Lp��./Ve��w�5��]�N�������V�@��FN�mz|q�K�/֚�>��/xH�� �ۏ��B�}�`�ƚ��q;���y�1��Ӟ��(��d|�:C���H3c��<� i��l~Ոn�yS��z����֥���̷@n�sH�:���۾/e��eH��o�� �.77��)�;��o��*�@��_b��_��6XPJ��Zuj8���'�v��Y +�_S��2C���mlJ'�!\F࿱��h���^=�=���m{�.%eյ��OMQC�`}�&mE8�����:�1�����ܤ%�ӻ퉋��ߙ�r�2�)�!ST�~	�a�)�K��ZlpB"��.\z��ߵ?��;�%ِ�}����Zx���^x���-�k(W�2�Y	�"?�M���D+=@J��x�����`�nI7�D���&�C�☑..{v�A�JS��d����>:-��d^Ǧr@��n�Q��^T�߀���K*c�.kr���-����s��B�
=ˬ�D/y��Fɨ�d�b����-��jr��� �9�cI&�)����ݝ?���F8��n�o^�(�_�/�>��c�����փW��hq,����ll��G�;�.��$.�R}V���j����"�B�kT�~ڋf����yy'�#Ν�o�6�mC�^ALԯ�?mv�����3��w�I %���{�A�7�7�q������t���;�≫��fI�p��tH���}�\ğ(�[�'X�$����rw�r��v 8���$��,�/]����e����E�j�� ��J�[��O�ѦN��e��I�+�4�_Q��E�P-�Nr�U�j��ᱻ�Fba��'�a�c���kr��6Vw۾��^10U�y��I�ߒ�2҈,��~nd0���e�ƸL�����a��o׼���~�s�����D���6�.SD`� cD��S�0&=�`\� �Ua s���LB\1����0��C2��c���+�T�`���Pg�u�j�?��"����~b觇*�,�z����3���1_~Y
�v�64MYJN�֫��R{FJ^0�gefu���J�8	0�s��� ��-IEH@�nR�:�qߚQ�����Z$�)<�xs�Zn8��	��!C�ʍ��̬�W`���k��|��=I婝�c����@��!*�����������1h��'RIj�'�&�.5��Z)3���VY<�v�����z���_�/ʇ&/=C��6�������RR�'�����Φ��Wh�3��5��>��/or`���ؿw�,ʴ_��h���M�$g+�WBu.S[j]�E޸آ��_������bfO*��y�b	d���S[���c���T���X�p���:H�D
�b��NgHf�Z_ׯes/������"~Ԧ'������x}Ӓ�8/���2ϩk��X6 �?�X23m�.r7柔�����!vaP�/�V��+%C^���yoL��}����~�O�z_=�u�[ ��+9a��!����y�'{01?n�����'vh��fL�b@)k���h袴@�1���u����7 >5�,r�e{�m~�2(Ly���7H�������R6���8Z� yq`�h �A�_f��<��˃��/��"4������5�H��j�ai(
�������b���IC�xdw!��V5xM��0sU��y�j&o������9�t�#I7��a&���rnF5f�}�"<M�u ]j*k�~�/F��u���(\�.���Ym��p4�{T�d�V��,l$�A!d0S������)��"��eâ�����<����IȮ��[�<�r�r��k�b����:��+1�n��>0�ˮ�p:��@�i���B��L�pg|^�#]x�4����v�
�c[]1FsJ,��K�pQPd�辎�?��2�h�I1����?r�C)�^� j�U�w�i�C�����<������UWVI���q/4n�&�pլT�l-ו[{�a� �i�S",E$�1	��×��ķV��5�����L�<}��M3�����lj�tP_���pOT�[bL,2����n��15�$����-�t�Kh�P�au������=�D�ʒJ�E12�-om��D�y��y���B�+߫�?!"���b �ͱ�A<���)z��qW��%[�Z���ǖdm��������~N���U����-��H��v�1�
�����̽���"�e~R�6j�84^���-����(�w����5���åʥTh�4��d:
���3��s*���0��^p�Q`����Z��)V�h�P��U %� �B��\HӶk���p7��A�T��X3Sfvvj�y��%C*�tXr���O������	�I��VL�:Y�>�7φ׫IJ���NHC���B���Xc��7�8�r�M��.}���0/��&�����8Q�[�MC5/u��i��C�B�����h��;�e�\��.#�2�@�"߁3f�$Ef�����:�1US#�m�5O�o����\�KV��W���E:N�we@�ͭ�?٪���C�z�u�Z�jV*��G�.�֋8�9.u%Y��n�V��Z�C_�Q�d>�g�Rѯ��"F�������}�oV"crt���$�paR	�֊IKM;͛"Ѩ���������C����K�<�&9'���yr�-�#�!i�h��\u�R	a�	Ml�r�#6�V[���Wc�g]~�<|Y�tR8�"�{�Y����l �	�વҿ�sv��*L��ݩ� ���?�+S�Dl� r|9H��6-�dK�["��0>-�|���$�����u��B��W���H��䷇4Ğy�~!����������v>X��i>��XdĂ��z�m	�V��~5������U�8TYXX�=�M ių��;��e�fS�Q4�)2޲��z,��T\\&{�}@�����hi���$y��Q��Ѝ~fL��Z�Ax�P�(�߱ʸeM���2��Y�{��<�V2׋��7��+����2�mO2a}J	:J� �R�{�X��jQ�hS�P�1�o>�D�O��t\�: kt#]�v%aD�
Ϡ',��0�T>Օ������+��к �N�e����@Vr�%����3���&����V;>�aPh=а�eP�we?����^-�	A�Y1�����%��j5�j��K�t�;<�8h�z%�Wv��A&[����_H9���˯�"���b����R�4�S <j�{��KF_��:U�6wh�o�j�<C�N1m��M��У��O�{1K�h� +�w��@��/*���zhu�)V^:����F| Z�J�5i���03��&L���C����	o"��.I]i(7R��}�U&���K��w��8l]Ta��Sf�b1��o
S��3t�IR�k�6]���#�/��{g��#N���_E#�J:8�>7ɹ c }vsȭ{y�WGJ71��A����.J+�;W'N��t����(
���,8���O
[e�md�z�aU�8���1�@r��l�������.��v�>1��y���AV�K	Ry� ]ǋޅ�ϴX��Ა�X�*H�j%|��yޭn�q�F��.�z�>i�wN�`��y[�}x����r��$87Y,�ܒ+H���u��c�''H�o��uK�?�C_���%�r�DJ���>r��\�����(۴�~i�8v��
H2'l5��~���E�.�5��:B�[jE1��$'�6Eʁ �=���!�]Rzd�Oh�u\�p���&[��xg��w(̖|��ltSbȧ���o̷��4�G�ۤ;���,\�R���U.|·���9��>4�.ި�ʥL���P>��:��wk;�U*�P�^=a��i��a7>��L	m	�v����c��h�D�%�4�K�Wdr���ܾ���V(7��d[��q5�N�~��kI�k�L>����v'v�+/ki	7�)@������}ȓ)R�e��8h�a�����^P.����~�-�㠧2���� ���߻�6��\^��t�P�¥,̛��|㻿��d��
�X#R닆'��|؍�37�R��QR�`��ܛO�wX�e�z��	�d\�S� ��)X���;���	�}�����j#�!��3�2la_���g���B�oq)��
G��t~;d����9oD�gp+��}�2�(h~�#�gM�V��/3���a�����W*�qQ�j����Ձ{�X�!a/�
��n��Y�X�I��̑�����\^¬��=bkH���Ll��q�	G�S2U�˸A=�@b��Nx1W�����gŬ4ⱹ��:��T�
R�g��G�����P9�xe,r#V1�U"�ꍟ	����Uф&���N�>��]���R�-n�!�����c�|V�I�p%�$C��VR3�Cq�F�$��c/+��ʞw*��#ql��F�4�?)��~���_c�}��bQ�J�<�ԍ{��95X(�ȯ�<�xd	�5���^�;=���_b��r�K�<��?�O�EҖ�<��OS�]`dz���'��'^�+�T3y�ʳ|7�?�b�~��Z��ѳf�T�X�y��Q��I�Zًf�O���j��^UΦ��aNؐbԽuC���,�X����': Ӎ�:d�PIc5-�<�fe���O��ٗȆ�6�����>�@d��&^J�Т�-�$"���u�؂�\O��5t�#m�������mƱ��w��x�*�S�
.5�� ����FV���֏�p��:��l:S�'
��gȰ<��zI[�Z�����+���׈R���ʪ|t�;݆����� �;��{���3w&���cF�\�D$�x�:�f��E���e�Z����t]9�r�=�d'}X���mz��Xz�_�t�No8���qт�$(���d��Iq��/xs	���0����ʿg���j�,��w��b�Uo�1/w�.��q���iG����
M�msi��b��y>A?���P�����	wM�}�ڽ��
�w�<�Tw�FA���K�Ŵ�
qb	���/��s:%��'�fw�'-�)���	-��g�"�!�r��DH�R�f�a�a�c�a�F�^�h\r}��yZ�}J,c����Eq�ו�d>�D�7'ξϰh����@t�k���j��#��W�����)��!G���X��9IUn:��\ݓ5*"��u�f�>�0��r)�m3��@��Oi�Ҝ���T�(m��=˹<@����<L�b{i��S�'�7-�51�R��f�+�*���ރ��p�����N��5&L��E���ٶb�-�CQEwܭ_���\q���Ae���xZh�4�nPn�z��ն��3
i�����^ �3q�s�ol�8#j�E����oc��a$���w��a���T��`cp6gy=½`�A����b�q��lV�F�Eؤ�_�Y��>��@?1���k$�ʫ�Zvu�+'A��3���T�@�9X3
�0���G䂏[7w	9m��k2"D,@R�d+׌I_�,�l������a~�Ss��s���XEOʨ�����n��F3����b-��� ����Cp���`W�_�ʂ�(G��H�oU�q�T�=¥��t�P�,I)`�d�0��
��h���'d�ˮ�$,�錶>�Qc<h4q�é���f�h�h��#LcFոZݰ��\���;�S��p��ƿ~:]���v:������-]�=B�b���Q�ED�o���0(���C��ík�#���'Gnye����ƹ�����q��8�dL��������'��VC�ێ!M�R{��u�1%AeB�'.�&4�-!A�
�|�1�7�t-\�P�|��ΫS���l�L��O����##�V�O�W��J*��4T�c��w�!�2�)�勤����,�]6>��N�����Tjm�fb���sN9a4Ew�=��#qr[Psd�`��r�ᡊ&�i��I��ŭ���G\�D�O2�$F��޶-w��纨��u��!/1������ٖ�
(��H�ov�̇{�a$���0R�Qn5��̐o'���$�ܐ�Dz�M	��O!�LV��ՠ\�,���kf���k�S-�n�7̚������%X��^�^}���^-��1�O#j`���+q0B��.ΚH$�蝸�d��By��&�h�i��S���	�*�Z.ᛗ�ľ$��gM���/5sga"z�}��Ն�|i��鶡xDa����D���[N%`��iATc$���Av.��0<�'>^ʐ����i�6����,Qj�G��k��X��*�Y�up�3��YZ���+��u��>��Xl&X)B0�6��ҭD�l�����u��9� ���/z�а�KcL��ڶaD�!�P�9
��W�ˇ��F))D��]2�dt{.���7����I�5}<=�{�������My��B��x�PH��&�|BR��cHsS+��ϻ�B\��v��ʔ�X��y^y�<��Y�=����*��:Kz�� �����;����T߆ia4<��F�Z��	���PM9E�B�+��t5{�F����f9[�N@���_��؄J�V1Z�n>/���W�U*���ϸdܭ��&�!��i��7�����n�Q8��!��F
,�dUjio�����7W�1��g�M���K���vz k>������W��0n����}ˏ�����`@��g�R	/Jo� 0])���]>��� ����ŎT��Q5�𢘨v/dȮ1�0\L�A��1	l���Z�Sϣ�����s�*D�����Ӣ'�β]uJ�Q=[۴��`s��2_�,\8gMS˭�0]铭ZA8Y�J��A����2*3������;7��0��y���,}{/Ϳ� ��'��=9>�iM�IO����Z�+��I�b"� B�R�H�>��}��5�X��S�Zmd��g���n��Ȅ=�oo��q�[�Ⱦ��`q�}~|���K�r~�m�mH4���Ԡ�RXL���� n�����c��[��~,B��-�����]� ���O	�]���t��t��D���0"��1�������;.W��� [�T�[�[�F<oH1�]�A�bw���)��4݄�?ԪV�� �ψ[m,j~9�)�,&���͑��Ύy���}�U&���[w��u��wˊ�B��^�sP�s�w�ґŏG<�V��:����v^�\t��@����c��|����ТB�eu)��]N��;�������v|ﶨe�?׭�$���6�DK��U9��)Ƥ��
�W�~+�KH�Vg:V���S)4/9z����j38{i���rF!Jo����H�����v�A_O���N�0���>��5 �P�L��?`���~ ���Q}щ��Ń!`�?��򲊆K�E�rn���k3Yf�,�OQc������U�.�h+����a�v��A�Z���9���;�yE=�q���lI�7�!���Yls��QQ�*O)�d_W?���[�����ވWJVB��������>1�W�o� q�n�(�4�%$���),O,����O��{��������hވ��qw�s�E��W��,��E����#zar��{a!s�FƬ�by>/�tZ��L�j'j�����B�yY&�@�V(�fv�w�5{�y�\ah�� �e��kٱ�i'�Ύo�f��~�Ib�A6F�.�[4�^���2j�s�s���G�1P���V�@K���[CFE���
D�����Y:s�9�h�;ιa��Mݢ)b7�fMڶ��{��1�~���-n�5Q���F���1�s��;pK�W�4��$^�t:�!���G;Jړ��/�S���re�<.J1�GSQvy�L[	�*�o|�3�Y���^����U�Īe2�64�l�� �~���Q�#u813$�1z�D^Kr�������i�<w&9�%Ћ��=�U��Z�_2�=��>������e|��{A��ŚP���ü�����]��۩=�]n��o���TwV���ɿ�\��!�ݱ��j��4D�-u�sc� |�M�ׂ�5((S�Y��8C�fvTn�Cc�T�$lGe!\���Y}RXSE�獥�Q����~	�$�F�ovS�wN�(�T���7`ЎnjC�v��4*���9�CkR��t���Xn���)�A��^�4�DY[�s��e����(,��j�w����Eu��>V�d6�H�f"ˮ���S�\�!�k����E�=�7��Q^�#М�������l���Q�؈�R7@���0���Ȗ7���2n���v\ʹu���G�bP����KA=ו*��4vy�ݖ�p:��;5�:�8{R���6骭�0�+,�<���'�;�VԦ�.9���;�/6�҂;�J�V�IR�
Q�<�I��M�
FA���>�6�É����m�SJ��Pc��L�`dSY�:e7 ��xs>��m9��1�K�����+�s��)�@5M���}�d��Ef�$�"J��5^]�Yf=��0ƞB�������s�1z��Q˳��°�$��&tfrh6�e6XU� �7�\	��M�8R�S�y}�Jt��l8����W�f�q��f	*RΤ��3���^Bߐ]�:��Bi����|U�����u5y�;|D4��~RKR#�l!&����!�������m+R1�O��0W��]�o���Y�A@գ:끌�[��֢���W6���j�y�d����`Cر�8�χ�$ ���Rn�A"-P]����
a���(���0�x�7�i}����i���l^֞����t�k/�483�N��:�侐.��d��XT��"ҝ:�n��y�j'ɛ�����0���2v(v� 8�eש:*��V���k�%?e���^4>̭��1��G��4 �pn���_�M�Eǭ7�p8~�5�NQ& *K�־)�!/�d���1|h ��N?�ˡ��J�_f���j�~$�j�����_�y��͜p�L {1X�S�yvJ��-��*l՞vCx1����`�I@���d.9��3W#��4��Rp���B4���Ă����nS�8�X��A�@����iiTy�ZB�FU	NL�<�*�V�����~��Bq���>���:�s~�CAu`����&j5�u���s�/���g_Jm�!�xz��N_��l0�H��b:`%���믥iF���#�l_8˗Ժ{ޛ@���oLV��&�t�H�#��)T���!��x�x
���s
���)�� ���m��6xLH��{��!F�iL����Eq*��ki�ќ��%��A
��lP�o�G;��M�Qq)3�ɥ���5a�6�d��n�ios�YŖ�j���ᡔ���+h����q��XR\�;�s}���Êjo���`�}t^�w�}/2F���n�i\vl1:�JWe����l�ﻛ-F,"�� ��#]Z�P��g���3s锶ݭ�g�-���*]��0)����Q��H��������L`��ڱ��
 '����Z�i����6��R/W��l��V��f��+�;I@�r�� �$y��bڲ\Ky3-���L�h�5�W���S�?W��r�Ctxp�S�Wˡ粧s�Ȏ'�%DO6����[؈�\�S,��f�/���� zE�2��w$7�� �\�kǴۛ���XD+8�� ���dfvc��r�۴MMW#�P����c���kYRjuc����H��:�Wh��C�5�s*�l������X��QE�-g�p�@Q������T�����α:aU4(B�53��_D�����NX<j� [T�i)�7�VFK��%B�F���O���V���g[�1vtE e��;9I
۶〔��&�䱊u��&�h�����:)m�C#�^~�?d4(-$� ���E�JgkF^CoP%z���jIǻ�$9����Jrm��YD-@2/t�{�G��Z&ޑ�D��T1��z��:�YM�L��0ğ}y$o�,~)]��ZTg���͜�"ŗ�A�+��������K9K�aXg� CQe6��(al9ے]�kM��r4P�ި��j��rHG�d+Kg�&~d��9��}��M<˄SE���D�k4t�\��x�@j2�x�+�A����?*6�Sw�/0�	���SEnYM
���'��ye
u}�� 
����He1S��1\�p�K� �w
�F+��~�\�=i�½ZҚAx�K��ҺygT�Ep)�اd�g� ͵>�u�i��ˀ� �� �Һ�)]k��C��/��ư.3Dr�k�iq0�?� ���c2��e���lc���="�F��:�����. �\�u��稠��b�F ��;/!7{��[,�����ZHףgN�}-:�W<��q�5�� ��+I����
�=b�y����7�~"����Z<��� ���ђ-݋�D���a�u�Y�[x�ӲL������̊%C��� ���[�6D�"�׉x��+���^�5P�5�qP���ŕu�X@��3�&�Y̾��N�p�̥����wR��Epu{Ă���{��VG��9�O��>{�ͅ�>t������1e�Af(���0o�LȊ��tM-�����ԭ�Q��#ZiK��=���Q��X�r}$�*q}(?�zc����G`,����ݘ����M ꑓ��Wal�,�nߒ�����m��;CC�IK�Ӎ��//b?��]}�O�����i����*w��GG����#�48��0��@�>f��GWJ #+�ȓp�a�1���}��ϕW!I�'٪���)�<gy�#��x�o��S;V�*���Ec��ڠ�����77�d:�=P���8��-��:�O2/��r�ez?��53\I�3���DĔ�q(ޫ�1�y�I&J��м���o��c���(��O���DH���p�H�f��et�(���N����uS2B�<p��ꪾ�;��W��P���s�_����C@��2��(��?X���&RF|Y x�)SF�T�k��}>a�vŐS��6!��%5n7�?^a�j����;z�
�4X"�N���ζ�q0�I���Q��l�R"�n6��`�P���z4(�#�nUr��f�?k��3du)��{
S��?[�yr8�g�b$�~.�O#�����YW緙c�>���J�qs�������v�p��/#.3�㳗S�`M⃅�,�J�6|A#��eb0�����zV^W%�T�nAr��jS��A�V|ӱR����Z��G��n�Y��F<��4��5��1��*���G@�K���~���_Ƈ�]QE��3+���&d����l��37�0{�\�3�F�u?������&5(����2�2HR$��D�C���.���5�Sw�?���9�9c
s���:һ�Ek��X|��7�faY�%��.ڤ��Ɩ?��z ��a8�.�N~�:��_�y���ט�^N���qX��5෣�$\ݲ��d푕F�����gn���p0��f_TǨbhl������*V�����޺�gy�@��	
���k���?��^���%Z����!֠3��W�m�����2*��朱�Ș�� D)�z�њ�U���LH�?C2�U���d&��S-�=#(�L���k�U`��$�ޜK�)�ndy[?#�S	��0���|���Qf����&P�ۊt��.�Ψ���>��E����(�&�Qn8����ɰ�������`N�G���ӣ�o�AX�`IO�Ɖ�iD�o��K�秊�1h���%�z	Et��bO�\$�'k�a��	ipg~EK-eJÀ-;�	�Ikv�E�?K�:�O����څL'�&͕D�i����JY��Dw
"���`-�r�eb*��F�HhIW�;��f]Rc��dQ�p������l���/dĲ��OT?(��{�C0}yB�;�Eaz>���%>��=��+&փ�\�
n�KH{R���#?��v.t�{��U����I��NX�'�*b*0),O/�R�QE�c�M:�;Y�$_m���e�D�1T����^a|�ښi��r�7��#����~����X3r�&Vl�'�xz�א:cEz�����]��Uh6�,yS���?r�r�ת�ޏ���������4n��g;�?���ǆ�-^!�*��}�T��,fy�L�)+[���c�e���iO(ۯ�g�W����D/FB��4| J�F�{Ū�E�H%�c�p��f"V� ��,�g��)#��|8T�7�P��
O�E+݄H���\�AN�
��r�T�C�yV��U��O����$T��Ez���$��/jF��{(��ӽM���$��ZZ�-�Jv,�������E�Pĕ�s��إX�ᵵ��F�$�� (�� gȹVK$������9�� ��*0��(��h��+�?��ST� ���*��W��O���a[҃��l�.���P�ʇ�¬���9-�̅u04�}[}�jRB�-��g5�R���.X,�(xb��G�J~]#Bl4�J���v�v�΃�]�UC�y_(�����p�g�i�Y��7[��9h��M��\�=�L=#���M�`?�SF�vWլ�b��V��P�%��v�����~��4�˛�-��'5�e�Y�=!�Z�i�9pOi������3�D<>y<�pZ�x��I�c?���� p�e́L�l��$�w_ln�#��d��7�H�;X�UE�~�S�<���� o�DN��n� �~�Ť7/?��.}�d�U0F�K��M+�+"��M�^���ױLbS�5�^���Ӓ-dH�lCj��q�/�~t�����N���Fa�P:�C.��8����nhm�����Pmk�A��!%ۉg��hW~W�M��,w�Q��~C�طg�q�����s������<"x-�^pT1,Sa�]H1$�6\q��7@�N��Ćd~ડ��QY�nGaڍ^Cn�:Ԫ���#�i΄4m��FdQR���P����=�����0�L�g�u`�r̿��I�z>4���.�pN���Jt^�m�J���S�u�k
eD�yL���C���KS��p/RM��n[}�oU����z��;�_��v��ٓN�	-�b�dI�h����3�Ʃ��[e̺��.��0��a�1����Wz�8�<���4^?�U::������Ym������:{mѵl�qt���8��gĳ�
�5HU�8���F"�8�ܳ��;��6b3�L��)?0�W�&�֣]�z�\�¤�	.�9�cǾ���*����
߆��0<%9���}�y��6���D���؍�b}4Q��Zt|��4�$��k�A��՝	J�)�Sk���u�Ep4��S�|�=�y���<�Vu����N�L�2�rm_�HK8J�8�GZ�JYn�l툛�m��a���ۡ��ͫϡ�I:MզWey�8Ps�� �Sq��Q�f�jւt��nG7B�y��v�7��;��*G�b�&Ps��U0Xd�q۩+��9�"Y�_��nE���7�t��C$o��J�Ǒ�'C�?{�T����p�3]§��~��_�M��S�����^ )4��N�4�d�%��x��z�.ް�
Z$mbz��{�ae���c�-!�}��#v�4`����*Q�E���~ݪ�w\j�F�5��A}4���~v6]�i3�����#u�b�=ї�#��:�����Aj�~F�C�~��`H[�D��jx�EPC;a��z��/!uB6Sv� e��?�FT�����ώ$�qc�e#�Q�К�Sv�s�#��t(A�q��z�z�]�[���?���B���߂�8Έ���c]	U�|���j�A��
^	s7����Ǧ���lF���N.l]��I������R��z��JY�����Z��G��8�)B�T�_y`��g@�v�ӻ%af�Tp�ei� �T�o�:�h�0,Ga&1�M��?��N��;�����.{��M�zC�%�e�[�O��V=�/K)�>���R��:t�<a��\���rvm�m`���8v�[��o�
��W����RP���������[wW�='��j>�� #���� ���7��M�8:�w/Q��|�t� ��1�k]������\}�iT�A���9">'Qhל=��ޕ�;0��XO�C��g���%y�����i���[-'b�g�|Ē!���Z�o/lR�#��9qS�s�����*��r� ��l�"���S#ߕ��ْ�t2���z$.S�_�1д�A(����m���Wٶ'=�%�!i�
E�`wT���C�hreI�����	�+Ca�	:��a����) ��d\'7��2�hρ�$$�z�P���0�� 7��އ�M�����|:y�����΋ֻg����?j��h�%���9%�O����cO��N7W{��dsb��/0�e�mR"T%�0�ZHՂԔ����Π
��h�n����SH��z�<o�ܠߞ�����+kܱ�?�c��6쪌�i6W�C3���6�z��u�����9U�0w�	0��ỿj��-~�R��0}=�a��C���N���G����P��n�;ة`㶋��[%L0�ڰ�A���_Lά���z{����}׻�BZ���>�2I��S����>lRۈ7�5u-S!%���X"5�#t���;�~�S���a(Y|����g�kCF�RӗS�<���[t�Kb3�1�*�B�x����y:�wʰ��&��u�9!K�N�*~�����\/m�B���?��i�ߧф9�6&�^���\�_�qht[�#�+:�������i��Z�"�0JD]'
b(n�t�FNT3',������^D�I��"�	*Uj�njb���u{�vԾxT�T9AQ���*>О�#ͦ(���r��˵�g*Peͮ�|�F�D�w���5kг�ǈ�����t���Cg�0��!��,M�`� O��+�9����z�W�;������p�l�S�N}~GϖQA!�V�B&re�C��2�W��s���D �}!8_�!>�q����k�ܭ�{U3V�Ѧ��^�7)��=��eq-d�w!k��^�h����X�8h��Lh��5�2#��]d	x�2a՗Q3T��Pҭ����M�u����=����v0.qgI/�y���Bޜ+(�8<�0���IP{��%�p2�L�����?��mE{�.��Xa�Iݬm��,�%���vn��a��LJ�nG�FC����]�L�����*�Ԉ#,�4��t�}&8j&�Ek�^��������:]�sP�h�Y��c�����Q�-+$��-"�d\�΁�(�L�"�S��Em<�Q3]�~�;�Jߒ����!�����*<~�~�Ze(yv�%.6`\�M'0��5�E���R�AL�z�v��y�c'�O�_/k�4\`!�*�5��H%�r��'>�����E7����t�*T��糲3���Z�S�瑱�И@R/��ӌSK[���ξ���Ðы,FW*�P�S�Q&�}эk�a�gM�?���Ib����v6��_����Z�x�F=F\>�.P���6��Zm;]���C#���Z�~�����@����wb�(Zql=�e�&�!�RC��N����*
�`�ω{�8s�f��h迎 ��*�ja-9AvG����9e�~��ɶt�N]��]���Ȅ�MP�g�e�qV��a$?��cuET�����(ێE�i��$�B��%w��E�������q������Ʋ��Lx;�I|^b"���[��%��b���[�y@���L��	�o�u����4>�A�AB?j�Q3-��C�
��Emr�m�m�zn�T�b�~#���|���$g�9d����HCO����/���FX[��X���t���۞)��0*��7�<[1�O�WWN�������G�����s0x��+�pآ�"w�R!)
��;x�|��?���%�[XaO]��9C�0�����|P�3�^}��G�+,��Y/Z�_�����kTQu�C�t'}�Z��7���1׭߸�Ev�O�g}�Xi��K2��ӷ ,p���Z�&���i]��?7d�:�
�pL�t&I�ϛ����,V�ΰ�#�|���Q���Bڅ��E�M]��$Ju��"��;Y���=Qrh���F	�^|2U���ZZ{��+����ѕ��5�|�jr���TC��Q��گ������\��j�Л��~��N�`���t[��:;��1��F�%mzh�W�j@^���M�|9՝!�6#����
�1?���	��U`Ϫ�#��z>�cx�|��3ܼ�@c�eZB;e�k�BWj	�:�J�r4܀�ֽ-�����=<`��x-/��Wr�*E��'�z�?���P+�l���Q$�z��v�y�ұN�����h�"!���d���5����V�<�ƥ?�do�I�HlW��)�lD��L>Dz����D<�w����N�8Ƚ�
�[VQ+��[�^}q?�)�L��6[�$S�"�,��)|�y�	�|�uP��m���� Ѳ�D���һK�st�b�Ҕ���2St�N�����O����,x����3��PΨ����D�Pb�L5����YM�w6��+#{�JRF�ǣ4��aP��@���o�̓kL����Zó�oܕ+ �J�6X��|a�&o��u+��Y�͐��S�q_��A��4��v=7P��f�ř/�D�f�t�Me�7&���h �,�zPZ����o���_��6unuu(N�U���u��}>^�N5%��p�Ň
���m�͞�/w��A�3�Eu;����ݧ�����P!��ؿ42וE�����/<�޲(���)�����H�4Ǭ�=���bho�*Hl�>�_��\ �B�V��ǉ�2�ɨ�}�ǭw��0����S��K��.P���v���K�!K}���N�P�)y<�Ԭ��
��f5���!�g��zO7�b�Us,Q��}�d����������b��x� $�z�<��x:��l��A��nd�
F뚆�5}��O!�"~oמW������۲U�;���$�2%LN�[%+G��y>��r���$5h����D:<����o��l�,4Yأ�����6v͎{̗	�>��_�e):�Tɻ=.�uDn����t��_����:�P����"�1N��;��j�e�.��x<�0L��� ��[,<�UH�����:��k0��14~�R趘C�F��B���"T����l�g>#UG���Z�)��|ju����y�^�<��u����>��ӣ�-����� ��CK�x��͡_7�Nd�kZL��e���+�6e�G[˼B^
��/1��ڃ��jq҆����H:�m�N�=F.I�>���s���%P(�=O�'��i}��LF]�udo.�"���;�R;����{���.�ul�^���K"��a�O�����G�
�\"��{�9j
��m��<c=w�y����.^�gu��s��� ���m�����P_����P�)euW4<T$�_��#��Ѹٮ[�� �K�ܹջ�[A��i�H�y#Fa;G �/�������|p��r!ѱ��g�9F���j�Fǀ�@����Ni)��Z�#�L���k=۟5Qt4�X�ؠ�쟽�h��S�l/o@�
Bh������������9���\#`
Y���Q��S=Ʋ[��o�g�Iٛ��Y�0^/Z7�؏1
B���r�i4nCH}s`��u�C3��V{�7�f��R�d�"6��1���!S�!�[2��Hoe�7:���$�������P�7@�)�k�ܝ�� ����f���l�_����n�ua�0�ʫN͜'J��C������u����olQ��r��.�9�o����n�*f�۸����ڃA}�yK|'�Qx��'�)�S)u2��dV`�����*�@���1de� f��@�@��M'pY�[�>��͘P��&9������T0.�������ϥ������E�;+��Tl�OZM��wU\@�]w):z�I�F��w�3�Ho|sz��9o�jM(>�Ϣ�Jĵ��PWn�-Q�N+�Qӊm�?TY'C�3�Fs�V�Q#1G��{?ьe����d@r��J6�!y������3p�M�X�(M�;�)�M�h���k.�I$��#0aC�;��U�$P�f��O�n=���W����D��������b,��a����F���Ho�Ә���U�n�k���KQ>�n�Ȟk��t��Sr����O���#��Jb2%�+b��ElR�֍Vm�"T�J��6BL��$axc�����������y(�V�RL@�Vs/Z�{��9���}I�<9 �I���,�@�&NRV������`D/��>R��T��7�:K���U[�G�D���T��@��V�cBB�y����y\;��w�(�˃�Wr�9�����Gx��q�xR��3���а���6��6�����O "�#�>���f]�{�(�ji�r`���f~y��M�2U#8��bk�!�d��&l����PQ^�� I=��y�q���ϼs
�[��>���[?'Y�B�x.�fj.��
���]��� �{�� |��73�BӪ�=����K��X�T�ݡ }����V��%��K���ɟ;}��4#��c�4���+5��SCL��G�XI�����`��&�� 0U��:��Ƥ9�Q�e�j�d]��qo�e�c���@�C�w���P����WsqB(%�)ρ�7g�7D(����yayJ��-�����&��K;������;V���������s)�E�좤S9��h�W�4�F{̱0��i�x�.���{b�B��q>n����uh��f{R���唏��T�7�R�H�����s�\ {^ԏ�A�Ay��Ί��N��Jo\�>�ő\�"��+f�w��2� N��7$�'�\� -�5��ʣ��H�;=$J�@�,�ң]��&����jOOc5pI��Q��¿ö�4WHAk��j8��8�=���]��v�q
��.Y\?�pB��l�٤N�V"��>l������q:J�:�ER�]�:�-B�  �9���ŎE�c�,㕆(�ԋ�U@�h��7VxS���&)��l_�O�.�b�*�$n"W��[	�à*��s��c$�~�p�b���ٯFtņ4Ev�8R#��⫫�d���G�J�;%���5
�=2�:j�&R���Lxcx^Gn�g�&��ee*���#���W��B,PI��TDA� �([��R|Ɛ�';�{���|�mz���V�Kl/h��^�Ļ8��-�hxg�̙!�\$�8�j2@:�ɕ��-�1��ݞ>.��@%��E�٘���!m|��L,�	ʐ��
?A��ͥ/�P�!Z���n9�4,�Ftd�p�`6Nz��`e%\JmO������QNG�<�=��p1M���:uaAa��ͫ���=ēo}��nG#G��B�5I�բU���A��ؑ��1��!��}6�,��.ACo�cf�>c��ӛ:u�W72q7tf�m�l���v~zG(��l*�� ,H�&;i!O�Z��h��Y�����f(��Q1r�`/�6��緭��V2?������M^���
g�y:�I&_�>�W]�n[��oT�-�T�G 俍��qH~W0����8��u���L��ȤĹ���]U��1�-`��J�%�_[.ћH�?�yg��gH�"j5:�[t����4�v�)�zq�b���o���-c�B�7~��_	�Y*�|� �5���+�dۀd &o�m@x*���i�O!�MƀnKY���<o�#Y*��S�$nR ���C�yDtm���=6 �$L\�Q�����K1�f>p kT	������.t2�8��VX�Tr+SdQa ���֗+bk>s\�w�Y�E(�M�$,���#��;Y!����S��)ր)��W1������#�<�T�ŕ�B�e�	�ks�a�n���EN`64Ϸ�`�N�zQ�4^F7����7�Q�[��	8�X쉰����_��-�H{]#,�%���b	D�����I�K^�nJ���W!j��.D/�z�JP���T�>�@�S������a�0:+��m��QS��`�:�C����	}�E�=���چU�^O�8����_8P��=?�4~ׯ�N�l�s��"��GF�8�}�x���6Ǧ@Թp��߭B�-�cE���"��d�S잝�@r�v1�eA��[���_�S3�A��:�u�^L�DEt�G�Н�a��o��?{V���;P��W��&��*����,|�Y��a���i��i���d5���7w��P'�Hh��ύ��c4�hQ�g=B���3ީ<4��躆8�ƢsQ��?��F�����ˡf���M%�L�6�/]s..�E뤸���Z� ;�&�aSkk�3i����5e?Yv(�3�R|!���oI�/ڒv����V�b#<��u�J8"&��ӡŚcw%���V��O���m$?d0=�먨A1(1p�S�u���o�9]��"'����-�A_O����d�����|h���=oM�B�vv��Ft$�2
�����	oP0W[ ��{|�d		쌵���D��G2�:��Fr1�AN%_�_.N|��ʘ@�©�@d�Kv����Z��W�gT%��H<�0�YX�'�#U��}��n�3yF�G;��?����B��"G�f�W<�ro�~h���#���ȑ�����N��<��5�L�~S#��u�2�	0�Dc|���î�ze��}?����mh@T��vbk�4���C���>C��> c�0�ٓ�a�^#�F��?��Va�v�
.4f�ȋ���Cށ��X�g�6XaG�@�(1�:�v���� XbF('�i�c�Â���֘[�;���[9;AFl�ؤ�<k�
 }���W���X �>:#7\Q�b��u�{ne�\�9Fd���?v�����B�a��4`)��?�V����x�DF�=��_��{leʹ�����)���mD��m(���\u�!ɟῡvHX�?|j6��3?�7�N�q#Q'E�����-P����1��S����g�dש��]%#�y2�X:W�f��X)�,G�aD<TF��������|��xK�ʋ<9�F�ʱ�W�\�3����q�Ѫv'��ΈƘΐ�q��=F���c֑��pL�7��o�GoE�m�`�/��ҭ�Z6F��yޕ�����l���ͤ�K����7�~"��E�\�"W8Wm���w�C>Z)War4����.�W�ݿ��\���6=6 �o�آ�/�b:'��\�u�R-�¹5sRB�@�xR����Æ+���2��F��s���!@�YaX��L�:H�M�״"���3r�.����zngr�1Nk��r�$�t�5�%�)�2k]��N���U�o��9�	��
t���R������S��۱���a��Kz�+� �p��v.'5�p`#�´o�2J����(�M�C�;���\c����0���]R|�$�#e�k`�(0V�r����2�(��1K���n=~F<�QGhP�*�-�V�O �z.?%�F�R����?������&B���V��Fw���p�N���Њi�H�U��`n�n�C�=���da\�Z��^�0* `!&�~�󝚑�9.�B�H�"���$�d�1�C�q������<q��0՜�'G�B��'�-�ϔ_��.#��ᖇ�����n�Z9�8�r�\�(�+�GU.FxZ���p�\e��=t����{q5D�D۬L3�%|��_|I|�I��W���5����xQ}Rj&9�����#-�.g��;D9���U mY9&��Ű ���&�#m�e�S�0f�uh�	�Ũ�d8�$��{�>���{IK|C��YM~ѓQ�ǤI���1�b�D���~��!DX����Z�Ч��V�#�
�}
�Ƙdw�0���$rȌ?.P����ݾPq�׋�/��yM�2Q{c�3Q*�>y��X�^�<0lp����$�=V8o��l%Ⓤ�]-�5�����|{+S������hq:`K��#Qp9�I8���Q�����C�G�}Z�0a�CxzB�_G����Q��˖�3x�y�#�	�U����a�a�h6����Jxq��?��զ�?��� �#7��1��vS�s�op�s�L`�Y�`:0d��Z�\P�~���
\ۙ�5Y����, Bd��%I�2��e� ھk��:��42'n���Q�S�w�8R=�$ ����Ol� ��S*�d#7O�L/�t��8��R����������R�	���/7�	D%���$��J�>�!D<{�����\wӜDA�ɟ�������=��a��w���2V�&��]L�����$(꾕��J�9 )���,(����j�J��^[�n�X�.}�Q� 7v�<����ȑ�� ���E�H1�l�}D���L�^�
�����l�3��uF�fE�H�̞�:�����3��*��%ڟ壹��	1I&��g2�`��]��U8pډ��4�`q�u��l�0��5��N )�B?�]��p�z���Q���^4���-�@/���ʯPc�KiΒz!eyh U��R�Rz��[@G�5k&��mE�� n�;i�*�"lL���_�]�+��{�h��-�yf!Zb��'=q6=�R�_qW� �:��8i�3} 2�E���8�4)Id�b%
����pB{Ѯ�bq�ٗW�/�\��ݪ���wBbm�]�/�e�Aw��aM�Zx��U�p��HF�*(�O0>A�_�&�q�-+ԸPSPP���v�f��H��R.���5ir��1�1�!�bZ�e&>|��CP�+R�%ǅ�H�����~��K��F���JWR췩C��<����PK��U��ܼ�l�ЩM���>b���TJx\��$���m�l1�OWX~G�K-�'ed��v��҈�`�q�\k�$i��Vǅ����t�5�j��WO�0���,��m�����P�^��o�B�p"iǍ�
Y�7����2�E������^b����uv�J>�BN��c�I����
U�~?�����aJ
�x�\�#6v�F�.��FP�瘨��f��z:<d��^��:�E��9�v E 詈#7�ި+����'4��}<����:Kf�ďA/��ٯ@u���S��#���o�P��>iW�¢�s,�ſp�uf�&�D=L6²�����|'�8k��v9e����ʿ��Uh��v��U����GV{O�\l!��~Z�1��؇�_̓Ĥ��ㆻp��2�l�z�N!���Dͪ��-��+	 ����+Um	z,M�Aٍ �3~�-����(S&��<	�-:6�_/�f⾽��0�o�Н��2���0�k���CU5�'f��3`
�ȣ��)�`����gN�	���<�De���J6*�;u���ڐ�[��8��˙O��l-'�BPm�y1\�⚝��tN�؍�{��-��)�@k���J�^�|@����`3�p��ނ��'����A�O]��ۛ԰�(y鸼�5��]�j��@��:���*t������r���	CO�E�sܬ7���*��_~�ɲK��i�c��|�UFL��y1�+�5d�o�̰��tLiׁ 6�G>0��8~Lm�RH�o�9ch����!J���:��!e�n�L�ؤ�ײ^�n�c{����"�c5�7�i���@��9���N��гJ�5�-m�CCi�P�r����I?H�B�8�r�r���\c;:�U�[ZԱ݋�K�?~��.�W?����dE']4�}.`̂��o�x�ظ��˹�ƴ�uy�'P*c*������MD朰U�z7�*�J����&$m��j�n)ݨ���!S���l�����]yX3�۠�Z�E���Cs����I' �]C����:�,V�.��������B�\s��j�c( ��
��9�c҇r;ya��d_���-�z�7�]5g<Z���? ���O���8�ٞ$e���$�+H
��2�
�V�
�\�uL^��.�y}��Es%:���
;&��d锳~��`�@�7�/������<�0�FwS)rL��*I��GB�̠��g5�H�c�|/(=s�2ŭ����W��[�m�!��=w�瞀,�R뵩P��Q�g@��J��<ϔi\L>N�=�Ip��>�)5��ܷ�x>]�#a3��-.�*�������*kL��7�x�cMYKڢp�*�9��*֝����G|37����NP�H�^1���ԩ��I�Y�.�J]�X����P�q�)�R����WÒ��h�P.�\��6�p'"�J��N �xK_��x�m�{��R�LT)"<��,��(.P>K�m/:�n�W�v��K	���@��B�e��R�c�K����4�RWJ{B=��2!�s���W�b�����>%zs<�����{���'�!�J�Y
��s m�k��',��\K�A(�o�d0h����B�̨#����Kk���h�Đ�q��A��A�j�(�w��n�1�Y:��R`�H��f���?��/7R�@�\� �3�����liXC��ە��J��[\�٢sf7��Z�{T�ZK�2.��b�S~��t����mA?-5n�<��+:�T�����	�e�ی�WC��=y}�=n6j�A�foP�:�I�g
3���jK���V�NɂWl��K�=6������P���`aG��R��nܓ��6�$\�hB�C�%�!]�N���V~�%u��wM�i�8WG�<+Pc]A.������F�u�9�NF�@�iV���;P?��7�=µ�����˕�>�
�%��� ]�(���YEE����a8z��FegN����#
�����Z-tnhe���ʃ��$}(��±@��:�əb˓6�JG��, \�������)������*Ma6J���ki!�w�t#��"�!o����I�F�,%�E8Y7-�j߬kZ$�;��W(�ޓI�c�<�|C�1WR�r^��M��H�/������͒�á��]��<#D�+5��������&{�=Y[4}V��D���u*����z��p����x��j������~�uGp%�F�x���;����TNG����`��Mt���5!ٸ�B��g�@�C#a�o������E+2�,��v��SF�[����}��~.�jM��Q�&3S�#�c���-� �)��-��z��V�k>Ϸ�H���M�Y�:Y[�����2�-M���T�'�Ԩ��f#I��c_�eċ�|y%��I�:p�$��\��Τ��A�,���9�p�y����p�Q���}�5��MA�I�u��. �88l3��(�����/�"�rCp��א�l�C���	�T6�?k������es�z���_��cU���i杷]�g$�v?[@j�>"���y�Ua�s���%�h����R�C���}.�U���D��I�lI_{h���x.��;ԩy����K��s�!�oj1�����H%{��*b�����6��tfi��&p�������,G[������S�K?Y��9 �EsK�[�Ԥ@�A*�̓?ßJ�9mb�!�ܨ�4^��*R'�����h��+u��N*�g��w���dD|�<b��� �q4]��}J�\b�@�4���.Y"ɢ��Ȥ�ij��S0yw�e���8Ffv=��E?׸=��p�K�[W�PB����̗܆���J��y��8F��۰�Bn�T%̠���kz{i��&ѯc�ǸzD	åA�7X�d�vHT�Lp�Ӿ]�x�]�q!Y���"��'��<����׬�`�Ɠ�Ѽ��X��Sl �0�K�؎�����L�)�Sɀ���3�P�,��~Zg{
�9��p���;�ŚN�ECe,�����>��sh��T�T=�*�dloA�4�h�,�&R���3�	F�9�hT�$ɪ�s߱���p��3yc��l^�L�a�Ql�+>���x�ě�:�0/'����J,U�P������9�����[��l��)�����0L� z�AU�'�1�O���X�b���(t_�(_����ã��yܲJ��ą�M��G�A�+O'�	|� ��$*6z[m~����u�6�q'_(c������ň����,�8Ҳv�8�qc�)�rl+qH] K�/�c�9]�qַ+�M��*��V���c��e�"�s1�2��#�K̦��g�����;(�����N�59+�?��m��R�R�3A�Y�ҾM��p=����9 �oj�o�2�X�w��;g�aѱ �!"uX�.<yx�E'1A� �ͤ-2�]��x�<�H��*�)x�����50��ڵM�����	��� ~��M��r;������5���|�ģ���m�MW��8�xE�<��}���nw����<� ���Ӹ?Ɯ|���ApP��U���xde���Y�Q�I� ���hq0q	��)6�_V3�S\��@F2x߭��6��{����
�X��ED���"r�L��ي� �oX<���_p�L�_����f�����}y�:�:X���T&x���QQ�\\�Q���sު�4��_�}�4gÛ�qr&�ƛf��m��� J��#�;�#õ.J6�k�T��a��%�z
ȵ��SC�Z�MRD�2fZ��+�b�^� ԝ���'*��8s�/r�W��A�����~�eA��
��ckm�γ�V��s��11�����'�x�����?�hQ��ܠ2�K�.w��0c���+��{��m�VV���$JP��إ���3�ؿ��m���Ѽ�_$���$��)Aν�Ao��-���4��n��C�"X�ע �ܵ&�A����
Z;�G�6Y℻��t�"���S}�5a@�HJ66��V��,���?�������\��˞�:� Z��/B��U�̺V�NsOP��W�x�G�]�����G�ܦ���Tvx&�ߓd�7j�30@��n��j�@��`����"-v1V��[���6]6��EP�U|
T�������}�@֏�t�����)�&%���
=TVИ�g�e���g��q��hf1TU�C�<^I�ꎈo�(�Py�'U�����Fb�������>����mOyTSx�ފo�����U�Lq��ܭ�69[k�`y�����佚��$I���ϲ���t� ���h�ޱ/��Q:��|�tʔ���:ą�����/V�����y'��50�j�4�̬�$|[^�Zhv^��� ������ҟj�q�d��{S���ͦ.�,/
i�?�>Z��.Z=/���;�:�w�����5/����(k�r��Z>%��"�=�	3�G�����j|�Z ]0|����'C�F"�����Koq�*XB�q�F�iI`��[�邯Ð�I�-�V0��L�ןD����:�|��A�׀O�.����x�6?���t���3�#���}Xs/��FU80�ޟ7��	��I~9�!sɃ�j��pl�U[��	Ҏ��3���kv�ˮ���(���fp̓n*��K���u�r�ޣaN|��^V�Q��gw�]������#�ٯ �w���2K�gr~v�NҠ��8(�E�x�a�_���\'���g K&w>���#w1�D �̄�p��j?=���ȋ7a�̏���h�T�=�WQ�l�/!(���\���v�74��e��B�2+afWM�<^�_Þ*��5��$bg��� TJ(%���;�C2J�@A��0��C]�:=Y�jg��hʷ�Iq�/b���6	~m[�#��Ez�v��{�6
�������r&��
��f�
6��eo��!:M./b�v^GIe����<u����M���,���R�����G�3�a�R�%ߚ�)���aO���`� �r�����BWxhߧI�ܭv�V���n�l��Q����Z �P/�1���,~ ��z譙R�k�]��lF�
]ƀꯎ��^��P��W����qc��q��9g�oQ�����j�������Fk5���M�<}�VW���Vָ|��:���TsJ`a?>3�����7��\�����<;��U'���_� �3�M.��\Ԍ���+�����9�&5EJ`�h<�*=Wrb^Y�;�w;�����Vj5T�����`U��f"I��e���<h`$?��a��g���x��q%c5�����(KU �K���$��&�7܇�6O�A�>����"��	p�B��-	6ŉyvN��ђ�����d�$�z�*�����`�A�)AKM�̹|�?�ۅ�7����Ge���K�X���H��](5.q��N�e�o�㵈?�]�i�Fcx��%�E��SM�\��8L�����>��V�j|RЩ��7)�94.q�T�+�0�l���O��	o��� �ڼ��vC�F�:�Z��{2t�Qw��ˊ�T DPM��Y3׼!'�?�e��"B��X�s�M�Y���ZK��y��CZ��#�����yhb��>��:8����:�r��� �!���=�!nAJ*��WBtD(*iݱ�yøX���pU�����=����8},Y��n���}��ț,���;E���١9�ýnհ0���5���a��&��Y�����apQ�\k|�S�̶ ��<3?�<a�\,�;P$�J7fy���P8w)l�2�<�R�͓��:w+mpj��/p�o`<�D�@������)gr�,@n�A<��m���7u|mϷ7�."'f�O���9f?��sE�8$�
|�M*��I��ϋ�-�Pi�6��E��e�1"�}�.\}���u����l�E������,_ê �^�7B^U�/�E�^�*���Wj���!Z�|> LV�bh\G(������p �p=F��_��r�i F�Ǯ5���ا�h�#}Dс�,�2c6�bV�
��/2۟:e��N-h�ȶMչ���#�1���c� �sŧ�8NaW��(=�!<Sd��;��!��}n�w�$<�D��;$B�X^]����YK���K}6�~�qK6M��Q��q�Չqg�w%b	2�|�^���@�NE�.����n������a�1�#���A{5}�����u��=�׵��w�O%U!V4u��,0��͖ى��:a���.
�=��u?Ւl�G�ztᰲG���kf���1��dԋwt�`e����ߍ6��ފN[�;�ϋn�yz3��R�	p�FwB�-���&4�:8�A>����o�j������GH#s2S<kp��XSg����d\Ůo�|�S�
U6�G��)����{�&O��k��Q>�x̉g�^����j����� �uq��H�:��lh<�`��u=���[%��"�K�>~�v<���C#�>k ťZ���=9�Q�c�@�&ql�eݳ쇆�Zt���Eh�X(�V,��ϝa��D��s$�C W ��[l8���2@Le`��׿�)V>��lR
l��Z32F��w�*�,�t=d�o�L� ���@k�&�U���|L
ϻA��Yk;"b���!�h	�sqv�}���!b��ݙ%<JP��w��i*��8K���4���F�xU�E�/��c�@n���ycE�i�D�5|����'1��3��4��`��3f�{�H*!�Gդp>$�KAD�{�3Kt�Y��7I�Y�'[r7��n��2V���u�����Y��`5�����W�'U�n��U����6b�s,��K����j��mBo�y� 4��=E߹�.�{9�hh~�T|v�#����
�P+�����p��x@? �-)�+Y�9*��~`T�1i��B+h���v��iXk��Ч #;ãP�[�ⷋd 2V[�[�/$y<�:J+�J0,~�o���3-�����]�9�=,��\������o�ڇ6Zh�xj�[猙l~$�꿀v�su�M�o�n���^%�@�V�B���O�]>g�[���X)�]�X�g�t��"h��N<oa������{sGx���="�&��(�
R:L�%׏�o��CC3�thE���]��-k��{tñ;B�g��\0�&+E�!	q�yGK�cO*yM%�9����R�X⩻]VL��#�=�����ʽU�C�^���YA�7O�B/�X$��.�|����7�����������pXi|����7���kS��r����g��5^�Ɣ��F}.��q��<�2Հ����;���o$y} <����	����r�[J���br���U57PtE�����Z��E�&��0�h� L�↣j׍x�+�Ĺ���O�g� �k�� �:��(f��B
R˰��Nd�����#�o�ךʳ����q�Di�[E��M�߲ �Y��j��˯i]�h~g���L�ƫ��s���r���퇂��m:m�IәS"^�����t%�
D�X�Fm=�����pٖ�k��u��E:5�w�Q-��������A�+D�e:[�;J����he���<��<1�]�ߺ���?+<R��J@/AG����(�ݧ���o��Le�o8W#�/�>b��-]��-.��9Ut��j�[}�3�-?iT\��l�P�rzD�f��(^�!���r��C��fK��O��}��V��d��ԩg�/F�L���;D��+f�l�:��\�����O�t�H�`�ϋF|�D���j©z�c˼W�Ίp�Z�eM:<]' e��7L�R&�K��Y*]�P�X�t��V,��4(b!�U��b�CG�vР5ݫ�O�4��<\�Y�M�N�R�K�~�>6��,�	L��t8r��]���������g�hC�C���X3�D��{���ES/Dj`�|���v�	���--V��o�M3^/�\�S�J��'+9������7w˜��	Ɩd=�c,�H&��tq��sG��;�#,fxN�bH�b�gQd�P}���^e �zh(P�:�.��X��G�?P��e��/`*��&��KT�e�{�Z�=�U8�7Z?��aa�RQ0&�1*�T��p���ރ5�G!>�S����G�)�+��1���5��>i}]�,mX��ӵ0'o*���Y*��Nn`�t�ۀ
�	2@�!+Ln�?��c.f����-��g#.Q���C���8�n�X42,��N���+�e�������o�e?�C$:�#����?鍂�UOE�/�oӂ�8�s���_:r�k��P�
��Ly��N�`DtZ�ߐ�cM��c|�n<z��p�����{� ��}J*�SL�����Y�4]�,��R�ϟ��!c!K�`.���u�
n$}f�*H1r�w���A�݂�9Q��,�0�DF2�800�x�yJ�bݩ��y���Z,t��m����ZZ���%�Lh���*�~��,\�!0���T�R'i��lPK0Z1]dI��U�,��eVG�^3��n�B���l��F��a����.hlH$� 1��Q��s!Y����Ìv?���-Ju�x�Ѯ���;u�G�B������$����� y��|>SP
U�����|�Ư��Nw۹��r�h�I6��ɝ���X���=~��r�лw�����߾�W��+'��TbhN+@;�}F���2����@�-@�$=��`����K�|��`ӡ��t p�q�L�Q�K>��՝Rh�ri�#&
� _`P$�L�ry{O"O���[��z����>�x���I�W�u
*c�a������f���t���q�A���ٚ䳱C�;۴D�IX�$��öYJߋuЗ�#rj��BָZ{��$@E��,NK�8MBB�!?����on��3L��ϓ���e�2W/r��zl6 $�w7���P�땖0��~
���4�m����;E�B�X�|Avm��v��G��l�n�	�fO�yydGp�}*;o}k�MV�H=�+��D���_���Yڲ*#t��R��Cчѵ�ꔨ��ś?#d�_�g$+��fk�5X+6��Ne�f�f�i��{�	Vd��������+�Dؼ&����§����:.���ѕ�'�0N���=_Ը�xن���Ӥ��I��W�4�w�_R0�NW�,��e�����|=�	�Tg�T�Mc\�il@�Z�+�Cr��}�K1-��� �/��C�^h�"!����ƚq��SB���lW��ԘM��B�4	�v�g䣜MTd����"��S���md���g��{���V�Z�Ҭ�XGm�f5��ݨ�y9��e Ue��i����I��^��a�M�V����AM���4#��e���^���Ń	K��s*<~�}w�����r�|	�^w2B|X[F-�Д��65�T��7�o��}ZR����vW�Wi/!�2A�U~]��"oKM�*Ni��v�:x!�,�U�umA�"!r���O��*@�\����r�>4f�dϩ�����wX�Ϻ�}fp���+�TG�߇E6�u��j�i���cP��/�ݿM�W���l�T�� Y�7h��h2�2�ʞm��*
Mwܨ����������������сi��+�/o*$x4����ė�-ia�q7���l�n��Рh.�`Xh��!��~5�$!i�zߎʎ������~D(q��dQ��~�q�Z�U�!����QbaM�uɱ5���j�r����i<I`�%q)n����ۚP�w�Mq!��	Ǜ�{*%SF�l�K4d�N�S�e�3: Ǹ���@,(��>_���p�p�v��1e� ����
3��q�ܕ�u�!���s,z���۠�m�ծ�V0�8r>f��K�(Ď��9Kqr�r}�R8��^S����f�Qޖ���S�])���ލ�J!]��Г�ǫ0I.MBU�_ܸ���5̕�=����>�-��]�l��5���#rB�@��:䙎�+��ԞGƉJ'<=K>��gK�nG�<����mU��jP#����~�ze���c�Y�x�:��I��e���82��,��aq��O���NC�'�t���h�����[r"��S�g:'unL��-����ݡ֠
ۼ-qD����;)��?��s�K8�L�o}�ݹ+�wTo��ƪ���@M���nm)�Q�`N�@֯��t��~�?Hp��؋Kcqr������w6��6���śY�{q�+����~X�y�-5��3��4�~
�IM����Kb���#�Mˡ7�Z"ަ5�+k��Y�@ǿ����2�8,}���Y�_#�{籘�^%��ױ
��������+y�c��f��M�i���0�H 036��ԟ���D�n�ͅ� �W�s�/nX]�Y�,�D&b
��B�
�aH��~_�{s�>����'�{fk�K/fx��wT�N��I[9o�ݮ�D�������@)]��q����pԟC`4K'F�Poa��m���8�<�XD
tZL'T ���t��z�,�_�f�ؙV�͸���Z�<�nʷ��!��[�ww��%W���)��Lx���:�^�(�e��>�Gr��T="�P�j�5I�zCf;3�<�+�GJ'�Yθqoj�>�99HN{���,W�2�M*$t��  � �Bzg؀ �\t!��Y�N�DT�ƭ�Z��${��S�L�_H]�����{�
'X���&g���4��
��,v��B�ނ���ْ����ǵf➳&�����z$�zW�X�PƂMq:#���2V�r�=+�nU4�Q|,��nҭ������W��lJk����{"6�ִ�k������ٲWc!�=8qJAA���{�b���E�K
�
g���xɊ������á��11�Z,+�����!��6ڮ�Q��x���_�u�ڄ�h�������R�=��Lp$���7CS�T�'�,�"Z�
��8�|���5����f�N[����7��ֿo�@`iQ����<g������{�tK[M3��!����eL��`5�n��l������]��;֦��+�@B�C|A��Jf���ڤ��V/)Vju���j�h��.Q���E�	�2O"�����,)P�[7*��5�����s��c.�l'/����r��2)F�G��M\�\���2���i�����{L�����yhE)��mK��-�ۇ
k����*��ó�]@�HT[����.q���n�P�����5KY���>+�u#z�R� n�0���0��MAmް��b�U&+�zo$$^$Hax�eS�Cn�:�+�{����EV1��煤������g�C�m�����޷�a�q}�s����)�$���1V��m3{����@��~�X+�a��n���g�F �-?������XhC�n��� cR7������{~/��<}�>̷('W��ܼ+�WX��s�&c���z`L߬�֝/�?z��-�+�X�v ר����q��y���u�|��;D���%�(n�Ar�K]���I*���b��!$��ڶ�-F�������� ��E��58��V_�̒r��$$� ��`�Q��;4g�<n?=׭��G�m�p�[�3R׍�S1�D>(��Є�Ey�U2>V`՜\�f	�p�v$Fl���������2��7��/l}}fl�ܒǅ�H�,����!�U�y~����b8i�S|M�xAv>��´ ӎ砫:+����e,��=)�c�w�^��y��O�D����}���g����feE��E���}���٠���S��@����[���od=  MDX��� �(��޻[��m�-T[���q\`5�	"
pv�;��F��|�	Ku[B��DĖ��#����u0m(�l禋\y�NɈ4�u��h��+���/���|�d�6!牛��J��i�{�����0>��E�ւ���g�ע���N�W����|�rH�*d�k�>�Z"4�t��nx�_�C����#M���}F�
gNEj�Ĭ=�xx�7����?&7��g�����vӄ�_=����=l���jEh�e��MDl蔸�/�g��D�2��Ҷ�Z��}�I�eKA!���d��'#���Ow@�o��SN7��?ml�vb�a�[/�f�����ޥf�A{���"kBbtwc��ш�wO���q�+���mo-�f3H�l?�Um�!ȵL���|�T��<}YF0p8:mD t�0�܆^'e��,����7 |j]UC#*q;
��3)�����%LË�Oy7�Igc��5�G�=�Y��%�Hԃ���,�H��P%�v���R�+���0����Eɠ�M��@����Z��0�ރϫ폡�R2��Y���8K�:���Қ�VWqbP��ut�'���=�û�m0bpk/��U����R�]���U$V_��;�Z堀��C=����(��$B]ZE��Ԏ��~+�s7�����nr��F&�W�qS��q���ǫȪ�	�(C�)�Q��kAvv������d��AME��j�����l�檗f��d�kȆ�,F��lk?�HPu��¢�~:�6�Z�W��|i��)`�T�(�/]5�b|�Js�A�1{�t��(5Ǫ��5����ޔ�}��wl^�������~��*]�q��jT&Z���7�	�'mjw�s)ꩥ����T�(���b�͂pܠ[����W$G&�/H��q�~#}g
��� T�K�t�m�y��WV�C�������>�
<�����On)�:h�sn��^�Y�Wb�(2tk���v���>��
����������Ƈa'��X���,>&ݨ�d�,�EB�A�7��X���� 	�0t���XM�D�Iv���1c�hQ�/�9k@�Wo G�2����l��PG��E{4�39��q���h|,7���c�l$ִ�]x-@I�F�5	"p��@D$!�Vߥv��ͱ��y��RlOĮf��6�����(n��&������X=�������D�1��6y�x�(KXsM�Xp�QzD7�k��|-f����c{Di=x��~i<�-�-]���9��(�D K�'wx����ldp��vVo��Gy�;&+��ǽ��ٮQ:�<��Ud9l#�Bc|4=�K]|�q���J��䰪*� �p��i3��7�z�\�Nv��6�M+���gD�@3j «*,��'/_�Ƨ���[�s��2f����G9�+!�{��1}�o�{a�ܳ{b]�#,1r��K��(�Y�� *��z�	����<R��,+�+I��@����8.��D�3��׻Ӥ���c�0G���D� �%�"�Ζ�sd_h�6�%"�;����k_�>;��o�{��X��'���6�m�	L�Jw������.��[	z�=R�"�8R���[�N���a`�?M�|A��H���D�HnVf]�������uc!��?巖�lL���s�I��ga�������9���W|`d��H��<['��X���h�{Q�t�Ӥ��^�\��X�e�Eڌ��� nv��������ܤ|�G�!e�M,Ώܺ�N|#��cU� ��r��u���!���d��	�:"����Mx�7	��<�b�� M�S�$ �}�D��Q��}�ϋ��)}g~��D��a�ay���20�b-K�K��+��bt���G!v��PZ��8`U�W�g����&�jú!���S�e>���>�������Bz�Y���C���ٵ��Ԙ5=*��3���űl�����?�v���̳�5y��ܙ�P�U�mV_�?Wȣd� ��;@�{�)��{߈3��`��Q�%[Љw�R0@6��R�X��R��g-�,U��H���W�N��t`����#b��I�F�)��w�(�m�1F�'�F
0К��>�\X��g�t�B��ZO�K�ed�u �������&����RJt&D�������Qm�����e}n������24�=8;t8x�%�?)H�Z��� �w-'�c�G�Y9���Zpz�P��"��߫�D�a;H��es��=Md~�Zp�I?��4��ٕtmOM�����B���XP��������;7x��8/r��0ɦ���+5�BVÉ$�l"+��]?�P|V;`�xW�PD�ax� fA��iM��\,����T��6����H��)S�@1E+%���3q�_$�� ��)n$��Zڅ�.�k��^��00��R�Vp8�B����}w�<�8�b�`��$��*'j�3T�g^�*o����<	���)���9؄�D�d_{��pn��~R;8��Q��w�$������4�\B�Q<qb�ҭFd�i�S��D�Eo57k�F>��ނ�^�}�E�e����Q��b������z_v��8F́ ��wK��4��Y򰲝�:S�� r���P�50�$���h9@jb ?�g���}RH��qy6f׹xN����7!E�F����9�	p}D��j!������;��Ժ?_7B��X�:��m��Ҭ�]��xM��ė,�T30nv�׿Ʀ�<q VO��iؔ�G�^�LoGn���M�7�̱�E�Y��
C�=��E��x��w$���8� ���1��o�3:ܶ-0H	!l������/�Qf�r�N��Y�JL�v��+����ȫ�%�t@��5����<�9jG k��娣�0��cP�bZN���g=�vb_��P��#ُEg��K���;(�qބ�a��䔶��H�܅���$�s'��>@\Yz�He���5�����)�+K�`����&�ϢE=�1���5�O��>�o��R���eE�맔��d\��*5���X���g��32�0��H���W��1#p�O�(�r��؅�����8����:и��y�Fռ4���>��[�Cꮮ�֝�S���(3b�v%����A���R1���$HG|p�v���S���I%�m��ĭ����B��~�c=��]p�q�k�z]� YR�~�`��H�f�&jȃ.#��[��4��t�p"��od����c��_��wFZx��ZK��\�D7q��'�J�E\b,�J�1�J>r���.�OM��+��Z�h�?�=��;׺_j��徒?i�I~ȝ�)��a�3h������P��X� 䄲�Ѝn�61l�@���X�x7�T0�x:�]��#d�H�SÕ���-m����((A٩�ެ0q<�{�Yr�+�T	�j��%j��U���ڛ��l�fZR~�8,�V����	��X�~�{p$wRw���g^Ǣ�_�\�@f��C�u\G�Q��ri���)b���FP�A��z�=
���CkZ�#��,��n���c��!D4�������K�jSpy� vw7I�	�"�+������À#�V�B�ܟ\_�b�s��+T4�w.ty@���mƪ�s���l6P�%b��T��r�J���?HC7�����P�#	��4'&R���M��.�wK�
A����נ}H�u���΍�,sӂ��-��bܓP�kl��2u��/�FV}���Q��9@9�,�Uk��9^J%G���E�����N�Il:kP[�Hn�YvE'�F�b��rת���iH�eYّ�aS��j����߸X��E&4�@-����Ҙ��-��Ѧ¾_�[����y�&�Ny���*i����N�PqI�<N�W���i�Ȓ�8�̕�M��O��b�3㧏i qs��A{bXP�o�nCٲ�)寊8�����g?��v's�}��*[&F�%�d,l��F�B�g*��K�y�)p�aR�c�?:�ɜ�T�!Tj��o�E��>H�:)d���Z�E빬
�!�y��C�#+���;��@����]τ���Y��w<K�'nV���:� �{���0V�+�����o5��ঊ�BɘAz[;pƈ��\�{�guG����!�v8S�2Q��@��j0	�EaLy!��:
��b�괚>0q��+\�:$�_s�r�im�����y���<�	�4G���=<��D�;��e�7���x�F_�)�`c�A��I��8��Q�"(>{�|(��kU���R/�\�D�V�ɀ�6�tADS�]��=��!X7ǢaA�ˏ�n�-��9k5�v�ŹK���Z�!��z���T��n���Ж�^�gh���.\�0������SM��2H꒺
3�Q�f�:rC��\�L�?�
PǿKٛ��O�R�(`GW���<A�Q���Tm�r�*wS f�g�(>]��ˣf�Nj=�Ē�5�P�2���-��d����ME߾Ķ�����q�|@�i�U�C.Ȯ;j� 95V:T�O�>L� �$�����ݍK[���$H�C���d�C��&�m�C��9�(�I,��߉Epz[7��{���<1��H���&-�5e�9(�C�/i��M����X¨��LZF?8�5���|(��Il庹�� �� �4�T&��ܒ�3s�)+:f����+�<t�NQ���(��1�`&���3���ŕ"Є���Wϻ�dZxa6ɋ wp�*Ȭy}�*�Iy�ځ����:"��@v�.<󐙻��.x�0�F�����P}M���P(|�_�
�&U���������g�W�䭇�#�Է�K�*W����k�d� ��#�R�Z��n�UvŹ��2���S����i���Z�0���W�#������o	�uk֣���Dt|qґ�?�ԥ�Z�������
l�[ߟ���6K4@�\N�g���� ��Q�� �`/S5�*,08�OBXnr$P����?a��gOՖ|>���D���2����ţ9����Z�zծ�m�8j�V ��ɦ����ۃ�&j�(1�p�B/\Լ���P7����k*z���s�hR�u*f�o�#VH8v�"�Ź���jku�,����p���̤�kg��A�:xE�yp��|*�CN �pu(���v�T<��o�F(��] J�~��[��h�#`��׸�3��A&:��6C� ��G"��;�
�����z�~F�8.���Sg?�X[�9f�	�\�}�����"���K!Qv�bj{�m^0���m��[| ��6�1t�x���KS��N�ס�ހ角�;�#oC,d1��b��]�.�����pDL�(�Zx���󋂪��h�����4Z�>=�AV���e�UF�Rd4O�muwƀ�l�	���K}�Z��ʃV	%�>��1Ӥ���hkY��j����ߧ���ۗB���H��RĂiޅ?��aFŸ�����%��O��!Юxz�іBa츭�xu�oM�<��C��o�wâtU�u�p��S����QGg)6iN��®��wS.B�4$���!���ő��Cu�8T��3�!��:�|��l��Wd� �4G)s� ��4`jco]�(��Z=}zPG��E���?�X��\��ID�$T�oA�����Da���V����FY�8 πIe+�Pha��E�URZq���@%Rr���ʥ����t�� ���b�y�#12���f�V]�����\zo!�ҥ�5��دU:�&�ܫ�.�q1�6��������X����q*�>���d��W�i�A��L�D�̉Yxbo�*ս�Xؚ�Lva�y�'�P�ZI'��I=V�xu"C���Ӱ!+<�̇$k�s!�Rܖ���V���*C�p�mvW�Y�牂��W�,��} Ћu���:ö����3{-v�W16"�0"�K�h���h�LǬԽ�,_h���/�	����:�E6�����$��]݀����w��v�u�uc�K���H�.#��r�G����O��i��#]���R�6V�p� y`����C� �j�Kc�\P�Y�
��Uz9g��b���+���:m�3h���Ii�-�>�?s,-��w����ln�n\?C�����:��}�n��t.�DiK'����(�`a�kug\/rc�VE�@�tƩ��}�D�cq�?�1��^��7��CX������'Ɣ��Ӂ�Zcph�*�B -�E�vt{���� %��q��cR�#����k��W����wYp��Vh���5�2�=\�� �7�%�[<3w�ȩ��C�AS�ae厃1P >�}�q�ގ-w���h(�bF+��!��_��/���~ʹ�}��+�(����@:Qŵ���a%2Ĺg��Y'G�ӥ�4l�%�����\��#<#�9-q���N��@�T�Rцp��9���H��nπif�:V�Xw"�fhd�;q"={�PF��u8	^ߢn<�P����-�T������զk�@=b4�N���������$mͲ���t	?�Q���E��=��N��ٔg�B�A4%DH�5l���w�$�'��x�pmI T���Adyw[��h�g��<~z#1�6N�΢�1�F<3a���3�����!̜@L��!Qz�W)�k���]�Ƴ+u@ZP�0���S��R�������D4�%�hm��ٷ���N1�j� ����vsO�j3��`G���gIu����|�^��wOR
>�OGD�)����>TeX��bS���Z���� �t����D����73�gg~�S*���Ndxd�a"��XD�U\g�A��F!�BT��8	�h��2]�Kϗ�B���?��ڏ�4�S����L��Ϋ�{?Br���	V��u���a��@����o�˂G8^y�4��H�Xɰ������L�0;ˮ�"��̦d��D�T�cC�, _�h�T�Җ�L��JLe-7.=�_p�^V)Oڬ����<�Lz�(L���K�i���FnF;`��G7���ǯ-��߮��ķ7E�t��ڧ����t][��qi�8UW���Ǖ��P�C�R��Ii�d ��=26چ��P5���Y	z�+�t�Q�uG<�l�׵Z)9�|��Ѫ�]�v	�\<�*���2}����(ǒ���W��)F��E�<_�D�z*k�����)a�}�Nh�[�r���ٺ}���26(�6$H��ܴx�iܢ�&����`^u��߳�����nmt�Jm��+���Ͱb�j3ȵɿRf�d�B�"e�.���~Nq��c U�G�Bҧ�d�4A��"�Y�d%]���X�2�/��pz�_����PVh�#����Z-�2��tm%�RQi$�9��
SJ��;?��s�}���vńE�Bޝ\$�!�iN���휬�G� ��ySÂ7�Wx�T�n����]��Д��ҞPH�a��?�5pSv�E�txt��I��~���_C��L�}㩯O�<��foB8#�������ݲ��߫�Ǎy+ ��ˉ��*�Yw���[n���3�L�U[�oO�Z���!��Ea6zؘ�&�"��u�2��
��T"~���I���Q�X�x0�g�h*�,74�����&�7�hZK�[64 \�ݎ �Ww.��]{&h����e�B�F�BV��*Jr��3=lk�o�cȲ��]Z��_c�������$8�X_L ���ϔ��e|d@V��Eh��tc2�SK�
u�~O�:P�:dn"�������
��O��I�#�-��rhw�qMCo���K�o�+Wue���V����/�0M��O�
q��}���|��#���s�&���
"ͪ�����D���q2�Fi�{��^9���R[SG��=�?��R�MM3#�����y	��=�H���j��#�v��Hk�$�c��)»׳0��|��5�Y9�0�jz��^\�̙U ͺے��f	��#Z���H��5m�����F��⒡�����i
[�����r�\�i,ZE��t|�`���n��\&
�rK5~'c�`?�q��չ����D�lKt�g��)٪���h�h���Xt̮�l�6|G��u�s�1i��ap�㾏8N���ki԰K�/��^E����*[�r���T���+%C�����~��X��[=�X%��Bo-��8�8Ǘ���5�!�F�$�
Ѡ����?�T�H���I�Ǳ.�$���IJo�Vp�6_��1�Ua���ql`��5h�0ms��?(%�T=��a�.<mu{�Y���n g[�F���`[��?u����Ў|��	J�q�~q&.=wXZ�,H��cxo.�M��vx}9sc���_R�+���C^�4�nc�\d<8�y�#ǒ����f��;���er��eC�Ƭ��T ʁs�0fVW46U�?��&FK1�\��eg�(.���������3n͇ ���
�y��0�]���&�SjaTn��Q��B�����8�>�Mi$MB���B��ufW�/wU�o��/w_�8�J�G�A��'�xD��ů0�!�e�^�R�z�Uݠ�=�����^�4�-��e��s�����"kfŏ$�<�~�(��\gDy�to��{mK�1"�{�z�Fj�Nz�},�~��Pj×#k�6~���E��>�ZfS���T��4CqNkQ��4�h�B]��r��<�7��
�P�&����N&�Axd�1Q�\<h�� �y�TYc>��F;	�Д�0��t�-�¦������%�;߀���A����ٓ�{zFQ�5d�ga��fs�0|׏�'� 2�D�|&~&��۠X�A��jBgqss��@#��89�n�N� kX�������Fvl'�����+25�[?9~󯠑6̿^
�?�%9�D�ޤ���Q���w�F�p4��J߶�l�R����Ҳ}��>|����	�B��������	P�
���A�?]�k.��jO�N\�ǋ�o
8,8v,�ɂ���X��!��%�ק���ث����l�ʹ:W���0	�ބҫ����e�Z��I
�H��J����]��p~?�<
BZt��t������&g�#��	I���»��E�"D�De����ʑZ�������m���Ѐ�j~:$�P�@ �<�AS�p�[X0v	�x2IÀ#5NiF�N'��}մ�)��lX��$ʸ|�@FԮ'����e��&�Yc�U�Z�䶔����\XNF����i����Ц��̖����X�/�=��T����_�1CKF�'�)m�gܮ>5Hi�yy��"*�w��i��z\ҁ���@xq	<8.�=�'�|�ݾT�D�@��P�$�0�O"b�$���u����KP�HX-�S��$Q�A�����9K�V�>7�����?~�����J6�d�����
�.x�5�fr�S��	��$R�4���6-.]�脓�"k�Xk3{쏴L����f
hq���k�N�܇��@��a��jƴl�A�� T���m�#�ЎL���r;ҹQj>�1�W��sc�s�Y�`=���f%@����1S���m��s����H刦�|[�0t�v�!�����A�����\���U^�{c t��`L���Y�-�y�w@Ȫ��@�'����|}�z|��ha��n�8ncx��W4�4n|���!V��΄���	V0m$�{���4�qs���
Э�\�^���+�W7k��מ���Vר��1Ո3:Қ(�l�q;��ud�틊�g�Ũ�D���~���������e�ӓ��1V9�9�/{x�oq���@�X�w]\{� ��r�Kq���d�FI�m��K< x����tغ�#��DȈ��@洯��T�g��l���a�x�g�^�p�u������%Q�+�'M��N�<`I�:�Ѱd��aX7��s�Er�=������9��?�A
�m��A`Ѳ]83D������l'Fa��C���S��η(+�N�-A�̀!�c*H��|�6�7a)ĩ�qA��d��J�n��g�$,����aŦ�4qHB�.� �6�KC}5Rԣ��q}2$���?f.�*wX	#B_���ݐX�����{@j�w�.����F�E��$8���J�ݪ������&}��Ѐ��[}D�y��VN�Z�[E)�ޛHm�=���%�(㡧ӄ��Ry)z��',���\B�����fg�Y�Ü���Ü��z�M���P�}�Ѭ-,��Y���9��P>�[M&sѽ���� �gO�E3��R�-[��JE�U���3n�z>(w�X^[[y&��/C�-Ϙc�1������[�K������I���vĕ�9}�?X���0a��$TC`�Eb;EK�Ш�V$C��z9��겪�K��&��J%�"�ׇ�V�~Q��BXIC��I�%a*놀�特�C����2�2MP�i��~�@�E���ȁ/;� K���d3���U�@mޢ,��qM�rc%���U�mYEFޒ�a��}�C@Z���_	��n{�_u.�O�c *� a=e&�����	i���>;�h�4�z�r[����B���#�{p��\��O�Tۛ/�9��X#2ְ���v�l;..b`/�.H���z��g��m�)�w_�1��D�#�l�N����c�l:qm|;hx;�R�)��L�-������ Ҏ�G_�c�+>S��W�i�gy}����t���(n_@M�	P�q�;��`0��hęI��{1s@p�v�� ����N��;ݦi]Lb�����@�C��NK�5��o��s�#E�'N�� � �ۍ�������'����X���p�d�G���)Q�!�  ��n��eM��l|v<��@�C|�8��Co���:��Kw�Z��|�W�]�g�����K�[c4~el�V�ۓ�����G�>jt��ӣ�HK��Œ��ts��Gg��O#�^/z�k�?�[M�OAB����V� �%ᘚ]�݅:�|�$��zE�� �FxC���j������n�`�Q�ښ5V�O��_]:[�LpV�po����i$};�GX�EP�|>��DW�ɜuZ�Oye�1����P�(�����.�+�7N��y��ꇢ�q��/�J����D,��tش�0������W녧��<�����6�]����N]ذ��Lv���}�6~�~|)XU-��uK\��u�\�Ep���|琅�R��ߎ_���X��+ "����2Bd�FͪWGH�O&%U�|�`B�I��[����/�t���Qݶ����;Z�9.9��v��sV��A���;U�N��L1z���1�����C��Ƃ�?���m]���eRH���7��	3pQX���%��2Խi��̗�cj��8c�K����T9���k�g�qY�:*7���\I��pɡp��9�����"�����v����V��Uň�;9�,}f�n��Q�a���̉�-Q�>��QDh��+�G!��O
Ӆ���oP�h�G�Ϗ��b��O3�'�25��오B[i�������O�X��t��$P2,�>� ��*�Q���A6v��+WDi���b�,7��s�ٟ	�O�i]:!CY>��;�����A)����Ȫ"����\��f"��;�	d������|?y�G���k6��?!J頯l�,�.�b��^	bzK��t)M�G"{��ƹ��V®zI��ʄmw ��lx��&�|����+Kal|}�nf\��������Vi?������M�����_:�мЮ�s�6<p1�������v"L@�Ho�Ք�\I\�J������ʫ��Ș1r��PaEU��2>�Qݬ=2���1F��n��J".�8}�vA�ՅYu���>}���
�����R�,��ߟ�ר�m��$�uqw�_��.��B	$�I��m���	o��|�e�a��?�"���;g���M�
��Ɓ�}���|��"ػ5/���y�oiQ����[���A��r�;ux#	oBE\��� O��>p1E(:
�ml�H�b3��Y�|�.�w�Z��.�	D��ޡ.96E�
_n�y{��]��MG.�iW�4̒X��kC_]��>3X..c(�d��e�v塰%=�9��������؆먓kR~q���8$'������q-�� �����W��3y����.^�d�:��=
6׼;������1n�$��H��uo�/�K]�:*d���?!1tب2T����������&�L�I M�`��
R����~ �"�4�)u��D�H�O@rW�u>)6f7Z0�ŌxD�J�� W9f�ZyR�;`�'9�l��쎘Ao�V,~���e�����#�O1��1��bm��^`<7�DZ��k\:)�4~�/����Ud	�'���H����AU���A��g��W��'���@nfߛ�r)�@?�ۘ`�j�I_��Q�fA�%�ۛ3
����9-�3ë�z~�m
nW5������SM�e�:@���A�)�K���-�N�4yGO�uE$��!ͯ��
Ė�gQb��Zk���5ڞ��]G��U�����o�E�u�\��5�JxCK��+�O�և>!�4�����ĺ?ȬP-��+ DT\���\�Jnn\#75�K�s����:l,Ǝ{;�D��ڄ)**�޵�vՔ��w�^	;�I.���W��cg�x��W <=r�d���tZ���-$-w}�BpID��^Q���vk�3Sw�0sB�F�'c�q�fQd��U���e�QD�����Eȸ�Ey�@rB/}/�?;��S��_�o�իZFLf�>�H~��xy��H��t2����;���Ό-�	�#ʟ;@Y��時o��C��<��Ƒ(����|EI��1�w�!�hɪoqQ��-��s���Jv����a�9����{C}�y�0�#�{�����c8}X��ҿ���n�����$!�ҁm� �K!�Ǣes;ҹ�~�!DQUW�Sb��6FsTIj �Ԕz�;9�$3���hVk��O���*(ZҟA�4�yL��s�n4�D�ք�7R�B��?!��:k*{�U����O/��k�Ҹ�����G�YcH ��$pg�٩�5���ʤ}�����d����>�� ʈT;����)��2G�mXd|D<��55��/_��gE�����k���.<���ߩ�v�B�������/sMq.��#JM�Y2��-(Kх`������L/AYk"l�ImX���M����w1�:t�(�6Q[_��_�A+��T\^sh�@�_ͯe��]9���=�=9��:�����x��n1C7h�������T��q�U(K��p����%h�5V�'�y_L���q�8S˿��B?6F��j�!Y[�N�9Q�7*е䃵dN`?�V������@��v�'m>��r�?��^��y�{g9���r�V4	 �7$��v�I)����G=���� 肬�Y3�;�H�v���J��^'t������z�v���n������qF߇-�z�EY�* �	aiJ3D���1]�8Ie�醿y����t��N��ӊj�^��2�S�Y��C_[u(6�c}cku�i'4�ow'�7�/�^OP�S\/r���К�����H�E��׫��{�Q�q���#����*��s��S0��>5?9��H˫�'�GF����j�ݞ���oLQ��-|i+�_�Pr��@�}1{$v�-�[/z�����ۚ ��/��q�׸'5N����HEO#��kl��D�$�-R� Ұ�T��˷���ܲ��7��0�i����-���?am����2���+�?���rtF;q��8���U0׷����=b�%�=� �����,AceSJ�X�(} �:c$6歓AyP{����v�t��Z�����yG��Ҟ܇'�:!��A�4;�v�A��V����M����˞H�[���B���N�����;g�Jx�lC�It�UXX�t���@�Me�&<���x�)#��H�b3�"6m��3G�w�A�=i3%�R�>�s|�*��
+|y�f�Q
�]���6���N:�P�SSFˑy[�n��A���t+"7	����Jh���s��5�6�\4k��O���@63`��Plm�P�c�0Ρ�y�a��#��:����8��G�P�z�|yON�h���.��_�\	��	Hѥg킦�b�&3��B�%�4��Ժ���v��L��)�f쓃��僄;q&�J�Mq�?�,H4͂V�BA�K��"*eux3�""s;��  wޔM�=�p�H�:�]%�H��4����?:4B�ݣ��)�Y%�B�GmUe*���a	��@�Crb��p��LKP�಴�4�!f#_�s��0�XsX���I���s� K�"0��t�M�Ҕ���B��
�jֹz|Ŋ�F�|<�m�X_U���@�q:o`��2x��t�V鹓o�U��Jl9,hg�UE���͊��#B���}����x,��N���@Z��!��1S�%��w���v�b-����������L����;���IL��S7�8re��B��_P�T\It�d��b�@s�oC���(ur�3��g��5�fr����]��m
�h9K@��֠G��ʔ�1pD�T�a!�it�t��{]�������vH?{=�~Z�n~[pn@��d�����������뮰�՞M�� ��	\�H[��3ʠ���m��Õ*!�.��&��t*��.1���J�_4�i���I�� ��S��*������o�7�C��I7$�Ǫ1>�<�c��Ӈ蝊 �=Ŏ��I���~�Ǻ�&�&��n���t�_#.ۖPc��|v��+�1n���HD��� �|���2Dh��X�Z`�/
�Gk��6s`�hn�n�sR���B��N���oE�B��'<n���L"d4����ح}D�~�[���Do��:_�<Ϩ��u�Q��ƨS3ᰪI�e��;�Q\f0Զ
 z��U�z��}`mA�/I�R��3��>����#~jd~+�q�'�0y&Ǡ*|w��0�
�Cl���kN�8�hR\����f,��f�u�@�Ň1)�L	��n�UBj�����2�)�!E��!�x6��W[�Qd$�����Qv	��	���Y�S��n?`�`��c�"䔍��K�6f�B@�������B�6B����(��6��Pifg�mId�vʆ|'#����ca�Ox��0,G�e��~[.��B�2���ҘQ�D�4�.���Ԣ-@%�.vu&��|�҇0��<���H��y��^l	�Ēn�s0��W�)l1��?aPp攬��'����$��)S>���9���(����n�\^�C����Y��&������"��'Ya�0cqe��U6
٢oY�i��k�[Dc�ǽ��,�)��b2�Zէ~P��'y�L ,�ي�_*K���;����9m�}��eHD�[P�fX��� }`�>�	Q����nZD�
�!�N/�]�-yމX��:���$���me��W1��L�I��>s#wBf/��G,}r9�RG�u�Rk�#J^:�v:���:���㲰z{:�}7�pP0�W-�� ��jbzо�6�@�Gu��2ZUd�x~j<E�-h���^�X�{+u�z�곦e�1����$�i|���Mv��n��b�Y�H��a{Q�W�J��j܇/�|��ޕt�[�պi��AqX�P��A�h���jAȰH��\3;��ު{D{��ja �g��f6����t��v�G���ja���-M1���G-�tٛ:ɫl��Qǜ~�􆞨N�X�1�����h'XI���)/�w�A	��Ѳ���	?���&�bev�a�ZR�� ����4��5�P��9�^+�W_G�؂�h��Y@�K3���n���.��z�g���&�?�M�e�6�͈ЧR'���o�dZd�0~J�N�qsn�A[�:D��>\Z3�'�j/p� 1���7u�cep�/���mY-���Lܽ4��P��pg����D+�eMY�?k�����RԑT�-�*8�kN<�)�b9�����b�\�-1ԉ�J
�\B�YI�e�����#g��k�[���X4�9�hp�v�+6���@hM��5>�ST��xb"iuFK�#;*�ORUL\�>|�-TS�Y�J��� �p=��v��~��4;%>�������ZA~��@�SM�^��S�7��O�'sj4Ĕ��pe����,=�r�K����,	:v�*z�<�̴^Ʋ�d��d�V�����D��M��Pa���˟W3�O��S�f�{��9�Ɖf$���$̽�"٠�d@;7@�9��r���[z�۱<0�
���`�9Z���Ť(�6��U �<[�o��*��|lzO��H.�4Y���mn9y�~�A�s�]�u��ܛ��
9��-����RK����`�#�GZ^V��?���R��t��4�=�]֊1�uJj�@P�T^r�K:�#
���~Mf���RJ=A���ʍ�ORQ����g
��Gr�\p��*��M��.gMMҋ@=A���G�>��X��neM�׋����%f�6B��؀���K��C_p��OKA4�M9JZ/͜<`!,�$o�\F�二���F�=�Ŝ��HڿgO��,\\�+��k6���p`5���Fp��7����7�L��"������ՠ��z $(�����dЉ�0�	8��յT�@E���E��'��N�������)%�ײ�k�V�[�E�a��i.�]��+/��|W�{#��A�i�Hq
[�� S�<%ݯ�Ѯ��W�[)�a�BhT��nȀT٢��D9-�^]V�	)f/2�d�!���rٲ� ��D���I��zkz�>�q����胂6�(�泫�L5��11m2h~-��[��q���|E��q�����]R����w>L׽B# �F��LP����
*�&J{�O0��׷�Jʞ�~��!�j�^�5>��s� ԢD�Ђ/�v
�!w���#�K1æ#I��$@�
Ψײ+��H��zc�˷����S!�O؟�l��xݲ�����f�9{x�T	Դ��j��M�i��K:�CY}^'+�����.�?��2e�`'4������)f�@ɓ*m��N�Y8я(ڷ����|\Q���^}��db��@��U� `mZ�r�/���zf�*���1O0�@�(�X'�+kmh�ֳ�3�5��� �A�Y+/sQ�b�P�i�R��<SHT�5g����D��+�k�6�I�K�x��[wKμ[���T�3d�d�UY���䘷��!�z�E(I��=�{B���lG�POb���\�K�+�Xut��� �0�Ԭ,�0�S��	0��1�ϔ���f�#J^��Y`�&B�Ip���C�G"����΄���Sϸ�A�y��R���g�'k<��+���1�/�Tb-�䷤sfF��d���&���Ɇ,g�n�?�'U���6��h�DVG�7�f��1�2���.(�	��$z�a�G�����wYx�o�ʂA�ע���_�jⶵ���O��XO��Gv�oPO����m)����6�����6�-`�<"�ʐ�=����|���;�>�w�
��	V�Uhz(f���Q����'��4U�0���D�wM�3i��klc?�E`,�i�	v!��U�&��0.���.L�Q5,�47ݞ��W��胒媡0J���j/m�����}�,z!87��g�T�w(BݔlJ�ݻ���k�%V�ܶ�B���\�XY�3�V�a��7������_!�B��7j'#+:u��R,�� �(i�&��f�o�'�.�|@Ε�e�����(g0,����9�GK�A�N� �7=�7F��1���4��w|���@��
t4+��-qs����0TJ �p��F��q:����	�
��y���}�T!�]p�th��|���)��k.��{Fp��sw���m��:u�s_R~�(n����B��k�����eŀ�"Y�.�2��p���2�c�����['fIߝJ$����?)u�e��j17���?��Rr:p]�Nn�Ʊ�2@0�'	��W�	�����vԞ�F�)�&ZU�f]�
�ЀZx{3ֱ������)���_cB���iנ���d�L#�����w�u���R�
����E�L7J�,ĵu ���T����E�-�ʐ�8����[���FM�)��S0��K�)!aC��������яYuB�嶯t�	��fP7ب���{�a�"wV��4���՚$7���o��6nUڳ���=.��n�����H�i`^��LN�����۝澑��5�Ng�`�ʠ��2�V8t�%��l
�+����_�Ĥo����.)�$�s&�B�¬ ��zx��g��6����6���f���NY��K�כ���z��RZ��+E�At9J��1U�H/7`�<d]c�'�uҋ�q�6�з��
;甤-���&pr����7xZ%+�.����\*1���+[��PnM���	b7z;S-�{���L��fI_��n�{��̗w�#����5�J�����B>�a�e�6\|$KY�N������E,ȢP�s� ��؅�O���9����A����ק�<4����ċ�:xW��"��y{m���a�Kӹ8$#�s'~9��ϱ��֫��_V���t^�x�w�~��x#�-J�@X�>�q"4�E*�\8lc�De�=:�׏2�l�O�)�4��Y��!!�9f�1H�Lٕc ��Tf}ǁ�-*�kY�v���$��|�twzx��A���'��ZY�=�F�h�Dq����v��Du��f�էl���#l"�K�!)�e�m3w�&.
��	�JI��h�c��q���
���$�7H|���f�N�4Mв��6�̇��9o?��W��`v{����j;�5o!��d�7���bgM173���W�*a~Aː����C����elG�'h��'��nY"��ߓ[W¡:�[�6Ԧ��7sa�D���0=&�6}�G��毵�th�Fn�H��6�J�tWG�#�|��Τ���>�
�Wb?�)�?y�p�>`e�x��Ǧu��~�x`w��|��Q���Y�5 ��5��0��)�1�����a�(z5�	70a���=�p��^t��<���AF�4n�`>$�ʓr]_�PT�4}{@�(�e���L4�%)�.���Ĥ���b��fGZMp�������Pv�L�	�8w���h+LI�:�Vo�(������V{�zSY�	*
i�'(���s�ag*g�~��<qm{*�D�yD.�	���S�������T ���{x��^�16���]���T�}gi~S���$Q��������Tb7qhE(~WJk4�������B:_�~�'�٩�CfloQ������2����Y��j�	]�/�:T/���uU�~Ew��y~A?�Pm�M̈́�"$v���9��X��k�j��Z�C����sp��s �x��&l��S`Ne�fA]s˙�2X��t�Z`��Ҿ�r��=�'� ՜���d�Kv*�ܟ��9�U��Lf�nJ1k3�ie�U�f��	��
@D��\Wܰ���d:Aa �F+��wSX�,|7�����PC���~��E��8Q��v"d���(4&,|n�U��q:�xL�����Q��K����:�}C���D)����,�83�-l���$���)<R�x��hTB�zn�2-q�M�=\置����<ݬ�o�5(gQ�ss���Q�}0��ddFv�_�EG��t��L2)���|�5?����5M1p�ّ$�W�*bF)u�6�`�ѝ6�+���E.a���Uj�����/.��ve��g�
j�i�dF����Hؙ��j�
;Ĵ�!Pʴ������"Nn�S�
X��k)�Pr�K���ok鬴����f�"�!�1|���P�Z+g]�H��3�����̀o�˃>9r��I�Π�h@�c~S)��>�59M�t]@(�s�.P�<��4AX�tX<_�΢-���ԧ�X���o�1h��f�{ɫD���d$�ʖ�{�pm(`�n&heZ�A�]���h�Qq��]JG��00��{�������|h	I��r,[�9zΣ�OSށs.����+��B�Z	��W�I52�$�#�~�`�	�K�a��~��ǭ!j�6zpD`�r̴ �Jǭ�OX�~�Gc���<o��*�J����b�!�mM��3c����Vo��Ld�o�����I�B��Bܷ�]}�b+��r����C���,n�BB����������ō^�/���'ZFܰ�n�������$}�R��`��E,U��>�����u��X�PK���^)��ZR����t��������ֿ�?�\xK�2�T�E��P��S�}���:��� ��0�<�R��A]�D��!9q�(��m�Y��*4��˒�|?�턷d����3�!)���T=l��*����C��E�a&���e�53����ѕ���,a�--�ｏ&Ի��Q��ɒ�af#�8$�q�z��:Y�� j�&֓U��S�t��[u�r���h�թ��6��f��;Z�`q����)�C�(�"��sW��=��& �G��V��f~Z���oK�Уn��aq�Ԛ>v������/}�E�������9q���w?��38է6�śa��we�m	���%an�j�{mb��d0.֔@�X������2F�~h�I�e~��U\��Ƈ��E�o��ʒ��qn����̄��2>F�^+L$�V��J�1��2����Ts��Yda�m���J��,j�<��+p:%
�aR>�����k�uo+�BrJk��b��9qQ6�0q.p�>1Sc��n$ъ1.eU�Tp���0I��k�-B�ƨ6F�M��2ʞ�U�1�L��pݽ#w��QI�~ǉGr��)����cC"�Fⱁ~�M�k���C9�%�4!�}�1���ô�b��灸e�+e�ne��4�h�)B$+&�8n,��pP`'�ru��lH���ܢ�ӟπ)�Ise��RZ�,���k���6˂N&���Wg� S�A믙��d�������4w�n���K�����.�l7�h�S�h������|rP��YԀ�v����u��(�kG��Z2W��ۃ7��>{"������O�ӷ ZJ��@sR��p1���L������{ԣ�Iر��l���!����)��>?�=5nQ���������}o�����ĵy_z�Y �G����s�?���6r�{
�n��D�2YE3��Z�A�M��L��4��}3�t�:�`�ߐ�XkI���uZ�yO�[bL%{`�����8ԉZ4`���R�nN�Q�I��n%7e�J	�z�N��:�hH��F�O��y���.�����7���RG  ̸�W\�%�NQP!������P3f��>���{P���\1bZh��������S2O�k��>jVs�x�-����FФ>Bl*h�5Xa?���1��O�P���͋}�3&$镗�J��-��-���K�4�E�K�=��yV��cd7n��ih���Ý��d�pp�����T+qo�Gv�W�J�5�r�}��	������*��_�6܌8���_�H�xM��;��Lh82XTG�'X�,��
Y�sG�J��cB}4�H���	�Y�e��� ��M�|�߅��#n_���w�U��'�E���̵f:E�Dmrv�[O����m��G���l-��.�,�S�����E�pi�֖�[0y��tc�[�-��S�U���%�X�,pd!��y�C-5˪������ǁ~�d�L���(� ��2 �9�1�$j�Z� ��yΐ���}WqH��6���=��(*�1I���Qe.�q�k`��L��{�.x{6cs�0�SM �9у��F��i{ь����fh�*�ք*�����/��^�P���/I�ŝ�O���j�1|;�b��rI�AZ�Z�u�Q�X���L��x��X��`�e�jL�_Sɣ�4&�@�c/��"6��pjܘ8��ԷJ@�O��R���W��Ptf_�ݚ�������<VAI'�؈>�:_�XÜ��/�W�3yQ�N�Gj��;�v���Z���EY��ulv��j~�PM�>�6R������o��ke,��R��ϊ,� ���^�c�{��VԎ�*�TC�������DO��!Vn;�J�T/�֊�$�,2��-l#V���^%�`���)�J+}��ʅ�ņ#�Z������?�X�(��A�`^����E�VI\�4�su�e�ǳ^�_�B���"0����}��ʡiO��!�`���A�V9�m��M��8�`�S�n�t-�.6��y�0�y��s�F�3��ph	�_r���&�ٿ�uy��m7�s��Q��j��VFO���e،���{�K"�1@�5���h<��Uu����@
-"��r�X�x_�;�mV���P�	k�֦��÷a�� !��y9��Sl
�y6j�aqv9>$�so�d�[m��J^���Y%͂�j]s�h�益�F�;�׋8��|�M�ՖOL����[��D�� P	��	ݦ_k�۹I�/�h�xW��1&�9��|m�i�������}~x��hO���n��#zg���hc&!p>�;�V���<5o�B��=�T�Oe-��9V����iL��
N�B���SS<g����+�uD:8~ཀྵ��t��+��[X۞q��
t!��줴�`�iM�~�H}��� Nh�4����g�t~��y!���}��+��2�Z���Q�形������pP������Ӎ�s��5J�mp�Հ��b����TP�y��:(�Ga���8�j�T�%E�hv����ڱX�r:�w���i�-Y�/}�g���p�Wؤ���Siz�p1ًQ���}?��;��J�/�Hk4��L���z���7�'�ҩ��΄)F�
�RqX��3��]Ғw�;��rx���11��[a==��T��Uy�G�GN��uH} �{�îI���`����4��;[`��;��#��j,�YW�P�����y�jNm2�����b�F���D������E?�OV����bQ��2>����wZ�I%��r��?L't�Л'�"u��&��RA.-tβ��f�u��v^Li���Zx�jyZ�
��eR��i�u9y�9+�����`��ئOPQ~!x)L㞄]�����mC�߲��P�^���You8�);�1ͺ�߽C>�˓Sjl*���f�݇�Ŵ���E!ʣ���6�<q�Olyz�9]8�\�*�U���{^Γ�Q�eVQ�����5���}=�0u4��V^mzo')�߉�9΋R���\��8���ns`�ST�R�
<����4v�&��Wߴ PӉP�F��|n~1?�����(�W�־��X�S9�28��Hgz_��D��W:��D�yq���5֫'�*�]h���/K�)^<�@6�]Ҫ�i�I�`[� '���ʷ?�m��ߟ�=�u���[ps�Xݞ�{�;A�.�}*K�)��̽��X�y�9�P�s�f��.[nwԿ�y�,����󽛪xo�*�N-���=%�	Z���ɩ�N!᱀�U%�}�h��Y��$l^*�W�0T�*.6k:�In�g����//W�����L:X��=���YK�6�ҥ̐��	g3_;h�U�&����K��$B��<���B`�d��1>��K����*�l�{o@�d��g̼O�V��;2�ӫ���GC+sp�<��{����9�x&��͍��Ց�2r
v���g�k[ʎy���ZL����^.��{ �hb1���&4����?�;{Q-��mh�љK���ϯ���(×z2��R];B����,r�x���v�]��aMIC|%�7�{�����7�Q��a������hru͎^��,�x$!ݢ ڄ����Ɔ>Py!�E�Rr 5A�'O^4 z@�H�9j(�`$S�]���v���!�<y�U�[�97v�wb�����v#��L�׆uL������i�p�y���nRbdJ槎��|V�q�Y�����/E3yJ���zk6����B͈;z֖����,���mT�YgL��6X�N�"���c�/��;���Ԡm��A��/72���%:��K6���yFb�B���Ա��sNҸ� C�Gn����dm?��x�'tq4���:F<dwG!���}!|�A)d�}bc�t�Wm�+�����є�~�h������C�)�"���J���i�g�Ƥ���DV@�lEp�}�& �K�� v��e�����(k�)��"���J�2W�B�	���<��>�GwT��}�]��tHߞ���d#�YZ���<�vT�"��:<��x��C���kJѽ�xFtHIM�h6p+��Z���;r��F˭�$V�{�8��gj� �Iu��QR�"�����
jk��8��du��Đ�_�h
�\�����$��;���f������P�����xԄ���,\dZ� ��k���?��p��w�M��#��Ie��荜n�z3r�$��4��a�a���� ��<�H�ER���)x���n؉�[���ěwz��Y	�%L`.u�ц�x���.�U('��rpE�	�S/�lԱ�ж�������P/r�.�ک��`�̈`��YIM��]ڊ�8Q� ��9��QVq�S�[�&:�w�<#a��uc�Of�*q���\p@�s,J6��U|&H��|x�`qxg�=s0=�����|��U�+��� �f�>�ZI��|@u-������	���r/�Or�������%�S���T�C^�Q����Ö��a^�FN�V�9M�pƊ�L��;Yl���G�:AA-	�$�����{�@q����Th��	�g�n��k0�Q��VR�e���,����C�n���|&�����A����ZcE[��J5�.݈U?����(�s���+L��[�jJ	���m��KĜș������x�v/�Ϫ�YY�Crj�3\���;�:���2<젊�9�)��/1�މ��)Ò�f�e���2���኎�> k?����-J�I��P�lڨ.p�|��}��2]��Τ><b3�Q�l�]�~��H�ɖ�Y���!�4-�$�a�j�r�M�b��q�r��n`���V�<���*�-2jK�{���i�90��JU�$t�f��Y�s��O�����*���(�E�.��i,�}�㒅����qq����IXC��Jc�Y�S��&�D�M�O횁c��<��૤H�9s��P-�4ȎB �^\�i>�UUa�t7W�=|Rl=(YI`װ�+��4e�����h�LBb����ǲ��t���~q_* IhQE8��m�+ޟҖ]���,�#��b�'���ĶM��|`C4�͟�{��A��FL�c�G�e��b"�M��#aX���AL[AcY\3�5�[n�?D���a@,6P0�O��s�:b�g��#���
&h-(���7���r��8c=O�zXv�@K(Qs�- �.�Ǹ;,�
�CX�	�6�~R�^=�J/���L �O[zf+��������ʛv�!�O���{�\4`�P14�uj+?��f��sr�*�^tϻD����o1�P�@�z�s���(��К������זq����%��V�=�F��:��,.����#�w=�赑1�8Q�D.yB��#�9|�0m��o���S������8�%��%�0
�����:h���2zP�+��nεG̿�魙��������^�҈�Jv���*�]�!"ᗟM'�YQ��Z҄�Y��K�&�vO��AQh9��&*_+��z�|�{6�D��Wٓ���.!S�]i	�xX�L�s����K�o����&N���$2�^~[��Q���͗ߠ��?�E���{�g��*��!�Yn�'YV����A�Q����#5Wp����%����u��I�:����ӛ<RA�mK�'	�0��h�G�46�f��S�Ŧ����[+^-O�N(>��I��ᵩ��ms��+,*��AqҊRsqaBԃ�D�i�Qք��/�X{DP�
����3�u8���?4�t�s�F��N2"�]�|�u[u.V1�ur#� ��6�k�֒:^"l��6������Ҁ3W%d�l�l�p���:Gaz�(s���#ۮ:��P�O��D�igB׆�r;����YP�qR��QBG�fDɳ��]�r����}��$�o�:�<}�'*���/��.���,������	�G�k Ř����:f���ᒤE����̖�v�W���ġ����(h�[��?jo�1fߵm� ��.�5e�(6��o(O�g�خ�㔥�����g�+����k��\v�&+Rb;���(�Ja~F1y��l*���"U�ڝ���g&���z6]f�r���47�ʅ�(�hK�$��@��	.B��,.�$�&i����B��uA�
���w���L:�����t{��)P)�7������CY@�>����޸@�&\#���B�Z��-�] 5B5pi#��-�w�gD��a/ȳ�k^o~�&���?�뇪�cn����ԺV�fߴ���;����x?��(Nތ�ދ"t8�u��4GLؙ	g�h�R"sU��7��k��*a�����S��Ej� gҬB���i�8X�Q[˺ -KCK��[\$8F�E��J��J���<I�H�,��u�N�=�F������ڊ�FuT�}���NG��g^@2�q���î�|����{��E7Ec7���+�?���7��~mŋ�$D?~�8�ϣ5?r�©jXٙ�Ϥ���!S�P+D|<�s	*�sk�1���W��S�}��0���-+�F4"NMU� �]���r��gl��]ߝ�����̼v��lf�.*��Ad� [�j�$ �Q�i��`��%LO��9�?��Y��\ׅ��l�D��-�G�Z�Tϋ)���y2ய�8T�3"��5�53q,�T��1/��XYK�j���@���@�({����^ՠ��t��5�Fo���菢*���^ts��`5�|_�I��h�����M0�("��_��=en"�{�1x����,�Nĥe�r�,��VSJ
h�����%��JM�R.D�W)�m*����!S6+���}7G��e��C)����z�LAkS���| �k-��^��4�[���B(��i	�@-F��u�c�t�c6��6Ge�����p�Avm�x%i���#��0(�}���ȯ��4\��Ϗ����{�D[J���9�L�f�ArA4ZF\�Ԭ� �ȉؠ7�Bٵ��qK���/~�
m8��å#�-|F�'	U�<��0��M�YE�W���D�`.���%��Z-	�F�֚��`w�D�S-�W��N��l���*�T���+�������ٚ��CnL��n7��B(�#��4W�dr�@Y׬�[q�q�b��$�a_>��=�����z݃�ߟ�٬�Ӭ}��~u�¸RrH3f�>sDo6�~�#��#��eL��e�*�HF��H]���֓�@4<�F�Oӟ̓D�{>��6��ȼ`�=:fB$�Ί#T��I�懲1{ �	(W�7[�Ğ~�����b��(�[&3(Oa�����ᔹ6&1m"R7���{�*\l��f��J���\�-����s��gʗ���X3��X�SQ�*�>Y|�g�5��WoZ,=>LJ��ӔU�&W*�hї���c]��C
.t)3�����V������A)�n]��]`���':7`��]$�4�	�9��!�7��[��WF��|@�����Q�כ���5���9��n���px��Pws���'���1�$IR+XBb��E��]���cH��Z�v՗2X������fB�9��*��POI͚+)Yl��[��g��q��N�U����o!ܔѧ��G>��i_�������
IR���p��_2����#s"���z&����-d闵r&�p2�s���&_b+�tr �����>����?��P���&
��,(�t���FdY�8s&_ 5�?c�9����!�����yb��,7���d>��b�x1�0����	!�;��HɷA/��fuS8|���/��su�T95���B�S��~�a1�A��`��y�M������^��HQ��)3#�ZX�yk�ኬ��×����^�?(����H*-�ٸ���Ț2�J���#�0�0j�<;�U�w�O��f�:��H�4��m�[:������@���!U�>9�N����8�y�������1��G�@�%~D^��E[�1G�*����}�ූ�,�B^��kq�6�?]N����_
/�����h�f�M����qP�����4����l�n>�G��HH�dԞ��By�X�Xu����D?�9�}�@;F�֏��	��5��zLA`JoXb^�~`Cg*bo�@���[�6�iH���иo��٨�7u܎f�ߚn�������bbj�Z*��~h����'�FWZ���J<����YY�������cmMA�߷l�+�@��P��F��Q�mȦ�"@��N���!��${/;t���)Nj��d���ڑ7���I�߲�l�u�eC��Ѻp��҄�1O���#Y����sCT.��՗z)�HG����d�Ťv�;ﱬWPs�J�yoq��yޅ��I�7Y>�����&��S�)f=�d����νp�s;�#�r�=Uظ���ҷIu�P��۾�ܖ����F~F07-��n�1=�0�����'���,Ӻ�9�7S:�v�ۏ���-2k1����Ӫ��k����Ⱥ�z����ֻ(H�pUW+N���T�Q��7  �.'������ZW�q��������U�B��[�X���A��8��F���	�gO��<^&+`Ͼ��N��/����!0��-�	*�m�����<�z�"2�ꬬ���(v�0N3/��D���Ø�s��`��bم$�҈l��0�����*V��Y3����mgOW��/.��� �/��7}�:E�?K�@�F�J�@�%� m˻�v &i�8�\�-�N��l�N�Z����&Z�ɠ��eٟ��&{8���J���-�U��
�.7�����>d���b#jHKx �~�R�P����2��$i#�ښ<�=��5=X:c&�����ٔb~��ڵbb͑��.U-%t���߻����/�I�V���զH����H��!Fa��_1�$0={�S8Y`����\�m����'ILB��s� 8�F��s(v�A
��u���Ԙa��D(�E��GЙB�u'dA!U�\����b��=�2�׬�&��I�(�*0��a^ir�<��@wl@��-�U��Ć�ѕ�ڧ%ST��$����r��+�D�u�.��ţ��RA?�t�j捈��� �>()�?!+�.0cs�c=�p�6X��W;[���(VГ��qv���NC�=-��E�L���хz�Ō�R�c g)[�F�ӆ�J8��d��WL.����]״e0��Z�}�Osv<��1�z�ƿ��In^:�B~L�ʩNO�WPeA��UA7��'2�,��	a��O�S}�qg���f�B�"G�9B9�VE�{&�V��=��q�E���56��t@uz���-{2V/�q��	�_2z�/޽YR��l6���U��(Ku����D��^�k�I��W0x��mG(�q�bc;�^��[o��2��k��RDj���6��P(Py��7��u��~��X��/����1��)3�h��"��H�.���ϴ��u�(��b�k�5:~Y5��D>�B!	�j��Y��/��p��U�k�C�Bc1�Z�^Z�`�*�NZ��Q�Q|��(/%�5�M�!4�i[k�ي�Y-�`Ɏ��f�=(2TAڢ&a����n�������P"���j'x�L����z�����[�I�Tq2'�����޼J��'`�"��*�q�+�fk������׶Gb$�J_qX�s&޸�W��r�N���h�؋n�[�U&ߏ?0����N��ާ��.ZC^Յ6VG3�l�c���BJ7_&B_��?�@�:��Z�.�g�b5.���}�%��
z��Հ��M�;&սb�ɵ3��ZZ�ǖϩ�+�o�ۭ�WDO�T��}"����h����<����T�hSi'n*�N�o��9�
6��� �  �оhW�E%���#M�l���lP�(���vÊ晔�8�Ĭ0[�B���W�����D�wQpΘJf%�C���M�<���P��<�P�S�v����B�F#l^ZQ��S-\m�-�w���wz��aE>�~}��!�J!׸�\&����R��j��aW� t�X����������F�:\����tE��j_�'��{a�����Yd�8ہ��ם ������6�{X��I��
�w�aU�!:%4(�	���8��G��HO�	������f��
�$��ƨ�G������dP ��7Lx�۲��{�%qA�f�{��P��7E�4�Lr�l.�ou�x�m�wA�[lEM��ȋl� �h\�.!��1>ʥk�J:�-6���w�}%-A˻�I�o�Q%��򕥚�@>�хc���S$�{�1t}
6p&l����S�Bm��W"}�9�f���'������#���M��^�MD@�pcb٠�l�?���mV_e:+!�w���,���B���X�<>�N��$$-E�;k:I~��	��r%��ν�02Q��T��2���z���*�Sw0Ns�:�>E�sE�WB�9�x�Sb��8�S�t
���%@���w������>ݎ���DW��bA��y�^E7ݢs���,�����Z-�ҙD�\���%��4�[�̒���mN���"�֬��~��|�z��7�zŮ���֗����ur���PIt�6�y��j��?aw�������޼s����G�A�m�#	�����W�!U#KE)"J����@]�u�""��.��ܿ������q�jW{�����׏�[�&^(���me�����yX �[�ݶe���8!����k�-�'�d��.Ҹ~����5�凪��R�>֎���N������՟�f���B��H�C/���V�4���/�D	�����¤WhE��@� �U؎0R���f���W}Fm�^#R��=Y��i�"�V�c�t��u*�5̞��y��=m�+��=(k�n.�$�s��T�S]svٌiW����y��Q�Bd��:+���������Z(��ENL\^&�K�<��T�L���Z��Ir��_{zF�bJ��y�NZ�,�$o��-u���B��q��a'�BZV^Lj?�#&>X�LȻQ�7*%p�<�}�3�ѽ�f��C�_�'t#����Y!�V�
$E��T�w1l̟�glq.����]j�zj�1*U+��q�/X�͚1�����a�����Um:�O�A�W�7׼ә����?R(����k&����Skwy��%V{i�O5���S>>dd����w�����
@>�Hz���=��`�_���0�7`F���n�К���DV��y ����/�U�m������!�G! 鬭���-xӣ�'����~�-���-��9�Fs�*������L���^4TT�n��͘t;z`n��?ۂu���ydA�)`�<&��`�)�LzTF��z��2Z?Wm�����C杗*B�C�O;����|q���Pz2�l�x�X,Vs�~ʄ����N�t����<��D=��Tc�zh���OV{����7�؏02�)���I��0�0\�Y�a�m	�F��<�l���ub�Z�-f��������D�|_A��hp!e�,�2OA�t+3�At�V#������N��E�p� ���&1���
��b�BC������ 4���ԙ� ,��\�&9����p!O�<XM��aT/ݠ�<)說k����GXL�n��%U�-���&ɋar7$�*�,1�}I`{Ey�H�Vn�ڹ���+�֐�&�^D|�&����&+�k]�$�rt)�6�;��`���P:�M}�f0�9SB���^)Âl�������zɱ�5ns�+�>��)�Q��/������~�M:z1�8���~ӱ���Xw�'�a��l�꬜{�l����y��Az:&8W�dS���{%����ID�� ���(` ��4���1޹�IVv�0��X�{kc���'"����u���s����HV�2������ǚ�R�Q��x�i���
)qU(���� ������� M��=y�p�&m�j�l��=��y����o�>��l�֠����:�{������ÎQ�"����jju8�e�T��~��-����@�(�S��R+A$G���@v<մ_����ly@_�)�i��)�Hޓ~!\�E�0vr�G��8
�/G���%��'����z�>!������$#��گP��َ�s�1����?;��%e� qͳo�!�}Zs+�	��k�F!�n��ޒ���͆O��v�__��:�{w Ԓ�fA�,�.-�<����=,��d���㦀��j}ݺ1�x��^֣玆v��9�H��DfXI���[8��i�9eB׌NAD�u=ME�s�'\��~�|1�&���A$��M��S��Z�@]���DVeE�F�խ�T��+)q6��*��I��Y�j+MvHϏ�mTx���.���e|&wRN@M�A��͟�����\��pW��x`�����x�F%g��(q
�w5
�������|����@[�@X<��;�G���}J���(\Nnf��8���u���i�G����9��*�k�:��uO�,��%�`h�:.�i:�c�)�.�p���9�~��]%ݑ�����/�io0߆�U3$Q�~��.��#z��}Η�(�wj��8|���㛱G:�-�d�����R�i��F�G3?�*���1��~��w%Ջ�yNH��]�f肧طV��g5��{������'\��-����������)�*�w�laa�8�LK&�b�o��q��G밉	�f�ײ]�� �8��r9=��i��l��<�KҨ< q%m�;3�QtQBSc��&.��!�z�P����c��:YnGHG/}5$~��P�gj��Z,n�i�@��
X�fF�۽N�J��(�4�y�Q�.��<߯b�'�B�-��оʥ���a�'E]Z����j0��$;�.�w\p�t}�	�{lDw!�Cѓj5y~,:,(z�Lf:K��T�(㩙�����~�D��^ �G�n��G�������̺m��AvN�h����b�4�6{���	��h�6�����J�[O��JS�<�a+���-z���@?AL�Hh�l4Dם�.�\85 �m|ĕ��H����/��	�#�XbaG�؁סΫĊe���'�蜜CP�cd������2i���/�+IR������l���;EDrZ,b�����^_��n�F߁vW��b�;+8kv�U�9�t��2�=��Ku��H���?�lOr�5�o�yc_��G6���|�o�ڎ�Old�tU̙�2����4�C)2p�C�k��3)ʖk��S/��\�^�����������Ň�K��@�P�Ð������pKe�)����nO������F�KFK׌�"��!T���4nqE�ۃ?Q�;�*���ߛ�_:�T���:����efvh: XR�yk͹�������#W��꼑u�0&[W�B��ק�`�9�P�2��#�zeIr'T���G�|��֫�VM�;�͏�T���C��n�;�`�lc ���!s�A;BI\�I�s�5���c*����6yXL���S��$a	]�-D��@���k^w ���χ$���|]R�R��H����
u0��۵G���������Cэ]NƼ�_��l�&�����x���z#$R��,�=�߲}���R�
-��:)�3��NX��.�9Y�J)��UE�w7x!I�f��Z�Xc�-"<�Q}y8Ri�nೆi*J�o~�ҿ@�� �k3�l��!�iO��ud���),6�(%�Wk;����Zd��\$@��ѐP����Q0�=�-2��Vd�D�=hȤ�Ӄ�U?UE�}K�F��:�YrT׍.���_]>�u�շv-j[z_�"
�����ɺ�g�3BS�$V��~���$�x�)S���@��>0�S�Dxy���˔q�켪�!iX�`dr��E���SG
����ŷ�eAL}.y0i㎳Z�)�}����w ���B�lP�w[~�f;��g
�r�����0�PC��2�9���י@��@��+�[���=lߗݬI�5�"j��!�D�����B�����6ٓ�`�l�8¬s
�Wc�s׏�h��X�zȀ2!��<��'ZGOz���m��^+���毳+
���Q�/M㿢�'�(Եͨ��Bm�E���c��k�i%~>��!��X�q(䣒�W!� q.�{��<j����� 1�wr�'�^CAga��g�(�_Ր̮N��H����S5��X���O�g:'���\}'�mhA�!����y6g�S�o#1=�3.�[3�T��M9�ԏ5�M�O�}j.����@�5|�1fK#�L����zO4���a�x��F{�:�{Zb�VS��\V�0�p4̶)v��d�^%"8g��!���A�Q�Z�	� J] .@ҩI�mjI��{����z}ZeH='��և�|�7Xѹ}���lG�w�t,O��������$����4��-�	�ъ�5�s�����<��xl:���ʁ��+����nD�j�/�Dӥ�c�?�A<��"C^�ˢ]�oݨ
��0`�	u��ȿS��؞t���,/��I-a'\��+�������,v)��nE�Ӛ��C�����ʍ@7G��↿Y�0�ԩ��x��6ٛkѪQ�rL+w��:���^k�=��x�`��H�8ij��@�
��S(:R���s5��g�0���ig�>I��_�exYN��ϕj�[�l�^ħ=?6�zk�\����{�������Sh� ZR �R�\�y7�M�o����s��g��e3^�z�3�jY��5�4j!ji�!�H& ���ɲ��"�Էؑ�as��Lq�ǳw�*�x2ڍ1�&�Q�ԓI�����[/����/)�N��0IYt��WEܲY��ח��وs�Y�fF����uX)(�Ϭ�M ܛ�%YR��� �κ�n�4�	Z�N����Y���s�=7���!�>"&MgT����|�6��	%u�	(q��a��g�L���� �@����%���K�#�L�`t���kq	zY
g�B��
��&jO�;D�\e^D����\�)�O!D�k(�L��O��W��؏� ��!`�lo�*���`~;��yr������A����s��F.�AO5�[�@�w���n������L0�	�~-F�F�J��$���?�v��!WN�e��)�`��Tw�N�}��RT�'	?�퐧�C1��y����>���|"^f2�7�����Iq�׻u��7x�3]��нذE�-M�H�g����c�כk�(;���� i\�d�[gx��sx�q	��q�B�&P�ތ<�#6;�Z��{,lY�ܓT�@�nwG�yr��JR	�ǉv��Q9\�Z��Y&�4ZqØW�3�փM�"�l��VҊ�8�1�X��m�|O��V�s#Q� �sI�湵����LX�YɉOE�$p�]�z�/0*K�	���~'��!_�W�g��I?��{^
'�X��|����"���1abCb���yK�Iӝ�f?]��ȸP�%�[�}R�`��>�{��ayM�<��w��C����B-�J��ʢ���M�0���1�E%γz>2ٸ�J��kׁa��o[t�-����o��j�v��[�_���!��:F��O3v�J�8�}n�ٵpP3���i��y\��)�ᰶ��1�ָ	ȅ%vg��.����zǎL)���0�����gB�_��dv�F��rQ������D���ǈ+��2@�4��g
��*�Qg�ʑO����+�?����t�f��!>(I:���+����B4�uo �m똫�I}N�3z�!�&���s�^J���b'���|8qØ䟅�Yͫ}=�ndtx	���e�*�� ���KO�0o��@Uy�I��K)-]��%��Cf;> 5ք9�F��def����#_�I7Y��
��\bT�f�N�U�+xO�Ej��\�Yx����y?���<���8q^�֨]���X���;.8����k�7�peU�a�:�N�T^x�|4���.3�5��Kj�cf�o�,㪙��� �H�O�!�lx��ZW���lR�$o�ĕ�5���Y�I{�H�R�݂�YL�af;���0׻v� �]Γ���OT7�y���ÝdN�ܘ��v��Mu�PT7�$x�u�U�w���9�(y�ѩ����Ař<u�i�Wy�[c �Yه0�Su�fI9#<��"dW,t��ѩƓ�-��d�S���@_]��k^Jc��ܵ�4�˲��9� Ν�qU�(D���:�-�1%^�((N$��J���'�.��������Hz�C�P��=-���GU�鶶�wV�RB���6@�{������ݒ?Vd(qU�Ҏ�������U�~���Q��_��m�^���L��Nќ��|��l��161]����.ꡃjM�S&�,�@�	��U�%X�h�n�b>����QȨ��� 1fLy�L��mN\}���q5}ÏO)�nI����0
ކ�4X�.�&����ZՈS��D�ܩ��f�hg��q��!H�Vd��7膫�$�|�}-��b��b[��O� ��,������:�}7�%��_�9O�;D�*�K��X�QӒ�^{0�p��>/�~���aR g���Ŭm��`����NcI���a��Ͼs.u�t�$K�� ��w�K�� �YN�壡��=R���FZX���h��Z̠((�{�
�u���V��ʗ�Ϩ$�q�z�{u�\�]@n����apxg�$%�ˣF����9�|�K~�I�����W����#���&g��t
���kB��`F���w��R��b �>#�=f.̑��yr�_���֚{�D���K�G���W��p��`�<�^rw�9��`[8p�Z�w}����𴤱��@m�P�<s�ףz�� �I[�_a��_i��nSC��a���.ll��$��^᧡�C����B��y��$�dV��_���18�uV��!]��@�F,m�w�~c`�".s=�� �NB�wI~��X��#����it�i	#8Y3�����_��[/3�h+a�!�z��������zQKS�m��Z�>�+��-�"đ��v�=OvPU���S�cS�^��&*�K�{��C��K�>�0I�Ϙ����m�v�Ao/~�#��xzD=���]��a �d�I$��x�sŷ�7v�s���3��ub|�k�-��i�Q��j�b,��\ �z~�b�k��L��qM�c ��p!P�7*�`.]�Zudox=��Z����{vP].AUX��8�s5��1�_�wY#;�4�na�=1�Ď Xx���M;]bz�����L�yz�J�!xZ��H�W���X�Q�q-6ڌ�I��Rl������6A#����2Mc��eh���$���߷� ��&'(Fp��Â�?��h�R�Y�'��O'̎��iG �$6Đf�{�3��#�PJ����WI/��]͐,TM���r���=LmqS�W��^�&��%w	�۰hU1�x�N=Q�ծ�����f���e������z{Zg<�l�8���W�����_u	� ::*���Kߵ�=΀J�����yR��E�h�͘��b��cc�'
�Ya�Ҁ;t3��"%��� A/���R"�o>��/�)�td��ў����6{�X�����ޚ_"6;����/<�a3L9O���qvc�\�[�r&HyÔ@f�%//�h�5���1�q�(����xdne�-�n����"����d�^���%�h�穮/�T�w[�XS���>k��iV�)�ˠn����!�n�w���/��tp�Y27�;����G���/��;lf�k� �>ūE;g���źp�FÜ�P ��φ��47k!�b�}�y�P�V���%ƹ�_�Do�4P��>����wZ��ZE�C��R�v��8�,:��c�5��܋��	rP�l�u<2��6�\]u�����1��;=�W0�Y�SP1��U�"�%��--HS01���T�;��B��ɵ6xo|�߇���Tꨐ��ۍ�7�}8�ʆ�� \��+0S~H`{���f��X�>�%�!d���4��n��5 ��8�m&M�5����ej �+�lK_���/��6��Մw�B"�,�M���"�\�]�Uv�^���*ҶkH*���LY�a��l="ot�ne^r���~�R�H�G�K�)5\��[.�L�����n�o�t�p�>Q���:]$r�]245p�w�Qis��)Ɗ^�=?&(D�ei+~�������G:o�D��sglup|�I/�ao�^y)�*��[�F|jNS.����g���rUj�ҝ'�j��>o��Ю��v9���υZ��3GQPI�I�U��N��ҫG��ͮU��s�`26�Pm��M�T��\�),T|U�B{M�}�<^�ͮ�Z�E}1�+���I�*��l؏�I��3��i�W�Am������ϩ�� x��iW*��bF�%?�rW��r����-
J�z�-;�qD$r�߬x��6ڦ�׿�:G�R�7��vZ~�c�l�N~�nP@C�u\a�C�)oa-�T-@^�ћ	���c��e�{�@Z�+H��%P�0K�V���P������6���S���,��H�o}�g�{�YӍ2����/����8������*��kUO~U(��������=�VB�a�}��+m�ӑ6�H>�,�B��A�J��Lhm��>��9�P'i�Sgޱ:qh����� ��jc���y�H��'��2*��M��8�b�>��y�����ݘ��0��[�~<�sVd4�a�A{��l�����Qݍg�4o��Зt��WΓ?�:Y�����?50C>q�* QS�J��4���K�f�]-$��*��[-?���C�t;wџX���J�[:.h/�Jbnˎ�hD���]�=�q��jL���f�M�ͷ�P�E��"�u�T�Q�����[;\Nb��k���t��͌{�Ύ����A��*!QD������j�Yѵ���p�]觴�v4hk�0�5"��3�n�-r`H�����8��J�U���H����4b�5*�x8D�kq����6);>�q�peJDV^��}E%�l�+SI�?d�Z�x;!�g����S��"�)���5�dΰƊ�|"f����V�	�$B~��))4�P��2=�wA�dB�E Մ�1%��Jm|N �#�X�3��E	�DH�P�c;������0,�cMK�_�S�G��Z�"��V��B�DB��s튕SU�2�7-� �7��O�50��mn��0���9�wD;9{���5��%�f����ܟ�R Z:Eg�2Sp����)������>r�I���s�{|�W1�sM՞/�^�Ɉ��36
�wxu{҈�[������Z����n�%B?%�6̇t��W%o�h�� ��\y�@f���qC��I��>Phe������Lv�KR8��I��z`��7���WB(o�35y��;�"��GJ�^�T�sL��v}&�dJ�]��3�o��n.#T{�����4cܑp��l��o���X:u�t.I�~U_�8H����c=�SS'��ΐn�:j�5�Ԥ3���ي(Vv���7���은��1�X��.��m���V��������[{�ϐU���TG;�MAJp���\XSU,)?~�y56���O�&��$T�QѪ�.2#����K�����w2���܏�����y�,��>��u^�Z�X'ʎ~cu��J��r�ԏ@o���o�o|�@�*wuw�Y-h���{����F�yJ� ���j%DT31�-ą����sJ���m�I�"Z�$C�SR�h���<�i�&f��4�L�^�wX*$ۏ����>�w׺�/�������T+���@�
�� 0����ާ!�����$�������D�k����Sj�S�cB�"D8*�`�.�j�㐓�����엌0�$���� �V�A�_i���AYӼʩ��L��,C���>�d�P��u��<uS�H�৾�+~x�w��"�NS��Hh�2r����	x��b{g�a*��)dģ��9�8�A��J�7���̻	���
�����N��1��q�Nc����z�Sg%��#$�S*������K���{������~~>s�5-��	��pn�&7����sџ8� �w�����ax���D�
��|'��9__��@vV�H:�#�dM�*}�9�rb$��H��f⒠�/Ӕ�6·�i:���7{�������.�rL�����)�9�nN�4|��Q�j���X�5L����B���]]&�)���DB\�o�����Or���Ǔ���"��[��j+#"eaP������
|��1�R��J�<��]�Mf�9����n��".RhB�$}'�p�� �M��b;��q�7R_9���{!�d%v9������re1�}S�6����gVo��1���nU�O�"�|t��;y}][�3co���@�c�"�.���K�e۲�".9����'k-��ݙ;�%��i	}�ǰ[�V�h]�T�O�:�d���|���H����D��K|�I������|����vF[_��rX��D�9~<jtn�Ւ�H[�	:-�A�×%�Y�~��\�#j���`��"��	�^T3H�y^�ǧ� nm��F{���6�Q[P�b��^S'���������k��o��l��<�be��,#�Ѯ�Mc%�-Hmk7(���*H��@k�{\
B���4\C�/�f���{�ʲ�q�cv���{Q+�T��g�ɼm| ��6rl�#�t����BJ��6�r��ư�C�#��ph�(�.�⬵�������m��FN����6�~1;����H�YT��`}��.8e���0�&��e�#��n\)+���8v��2�U��ٍ��
Bw���:N���wF��Ao�*��������Ͱ��Ɂ����/����2�H0&����[��%�Ĵ7�T���Kv��[ָ��+�tp �����˙G���n�~�RH=p �S�Ք��X��cv��g����P�w���4#�fJlJ0B��R	��
)R�2I��./0.)�߭[m�OD>���i��蜕�R������,\!�a�6�r��XFv:5�I����gj�,g6��:�C�oC�ՇVB �,������~��ђ�@�`Mu����A������؊�CL��a�4D���5�Ts&�h�	_��S����r&k^��j�����ig�K!�t�^;ݡ�ھ*���`�D��҄���鼌�ɂ���
�s�h��Uʦ�460Fx�F�l�|o ����)��R��f�"�����q�<8�v2�Q>u�O��h���g�O_9*�����Ԓ�5��F6��fCӉ���;�:��9תZ#�%��ܡ5Œ��x��fW7z�ߥt�l~e�<y�Q7�n��Zo�bTL�CC����Ƃp�6�+����A���O���Q8B9|��h(�^gxRr��t]W��vI�[�T��v�YY�]�a7d,@���5[����Gw�� j����D"����RY�|��lf�V����$���$�� �G���gT��,(�V,�Zѯ���w~U����{b!đ����'_����x�0u���Y�G �����J��2>M�WǬ܀�'���o;����m헡������>��mi{���^�w�*�#c�hBs�p����"�Ⱦ'��*�,��%7����dH�+�aG��h*����Z��h��©��Hp��2��j��ȣ�)[��|�'��*֛�=kDasة&7�R��(<z������̰��P;��I���$�7I�޿v-�s�9^A�6q�z�I���HlƆ��|��1��1sr�I�����YJ�� $��6ʼލ�y�U�}��x��	d�U\���O�0��������3�N"D.& D%hZ<篯�eX�7{z���)��щ�ݠ������E[M(X�`�-Λ.�1�瘄�p��C҅��;�&�:ɂV���pfې>0��\ Ft2c�|�|(:�1ڼ)�v���PO��{�w����nk*_��Y�/+8@det)ɔ���lno0�a��2^�ӱei�e�K��o�[�	���,��T�� J�F��ƛ���������ʽ��8t3.u��\���"���Rȶ�x�>Z/В���$�CHD���{���f�,�۠�z���b�l�����Mχ z����^�D��bޠ�-����r�_�&�~��+r�*�@�i���f���q3 �3���� ܽ�I��Tj$��q�Q���L�T
\��!�]��hS���hq�0y'P��Ng�2%LHj�����/E�-uߓ�����^B�z���a��$�gM�s�,�)���ߗD.�X�N��ͫ+��|��:{�Wa�g���`�;8f�����),�p��)f��D�iLg�Tj�[�BT����@�̭�������A1�ԲP�vj�&?���Z����&z|�E;2d��CR��,�S�B���І�^�# u�2����7.�t��y�}hվR&��q�@���{�9ND��\���CE3�@��"9Y���Nv��000sVN�n�m�#��W�ZT�XX��o�c@��UM�"O�W�D�+��7gI��j�[miN��kbܾ�4R� ܻhشێ[pƹώy�^@9j79�6՚������?��\z�8C�$)�����8TΝMZʑUq1����~�������4��x<`������A�W�"�'��_TC]�<�]	sa7f�zTZ#p̈�O;>�%�C�wJ�w�����Vb�H����oLy��ݐ�T�,�)�����?D
s**[�Vs�9��#��	��|��V^�ȁK�?֊�ҵ$bo��U�,SH�Y�Y��"�}q�e�@�sЂ�O��2�Z SK�3(�^�*`^��8���S����c���Ė3PH�=���|�0�?"b�� ���D���gUG;I����C��vHeE1��	���h��d�#��7;C��a�{g�z��8un"�����"Oȫ5�|�0�P&�	Jx��C�Jǭ>�o̟%~̓2s���/נm�vRޠ�*��5��;5rɓ��nR"'0�?U���m#N?�=���O�^zb-/����h��(�l[����򪘽��p^{=��p����\�2W�/N�*��S��N�lӝt�rV=���#�q@���H��P��͛��N��7Nc��p6a?����~�y@�a�%,��A[���}� �61�B��`�3�3��n�s]����%�5?�sWD���˜��5�=�p�����M҃z��SH�c�ss����j���q.rFt�%�*C˝u��<�؜�h�@v����H��T��j�8'�]������h�	|Z�J�8&��_@N�z"JpFD�hW�!��#l�#³»�2A-����MŁhG�Wt��uߩ
Er�8�8Yy/�*�G@�+gv�|�C��GNە1���[�)����n��$�J���/5N�W5.��r!�"�!v���t�I<V�4,��EP@�����պ[e�{W�<�m���Um��$���	�Q���ͮ���v�|��8:��q��y��yɬ�}&�J��f�g$�[ߜ���lc�7��3��>������;�`�1�A�d��;P@?p�w���oc��/��M�:Fj�ԗ�Et�"��:Q�]�ⱳ���5�u�{�]ڢ6�CM����
q��>�YLi跈�n$+��!32�j����\*��(��!d--ׁ@��# ]u�_�|�7_:���B���/��Z��fx����ռ_
0h�QX��x�+V�=zOe�Q��Y��,�Q*�fjx�br^����f����gr� +x0ƅw=rtʫ��G�2�?�se��Z՟�$�|���evЀH]�ya��������3pҸ�إ`?��}ta�5('����_d49:��x����&{c$���h*j?��;pJ��TT�^s>�+Gv�0����N̷8H��Y����7�3"�����F�rxx���%����}��6�Hq
��JC�:��.���c�����*3�#Y�M�]�\�|�T�t�b&�R����[�12�I��xrf���SO"�7�����K`�N�f?"$� �4|�@����+ N�q�@��>�!RO0���	Yf6��eUR0w8�+ƀ"�X��V��v�v��߿�L(��y�y�/?��__x�3x3�Q(Mʏ��v�k����?0�hig���2Ц��:"T᨞���}\�S����c�M-�,�����0w�+�k> �>{���;`A���N�K�[0t�R��B��R�@��M��$���۱`غ�jς���l 8��}.�R)<�����h`œ�(��9
b{�H��Rc�jHG��%n��W��#���U��N�6��� )�S��.���ʼ�Z{V�A�p�|��L��񹭳�.gO�D~~X�xĳ�S�����$�?M,�vtV���:=bt	������[�bĆ0?T��gb���*�Q����t�\J�(z��o��Z�kG��PJ�~҆RjK�í�UY�G:��7�M���,�$`���$hĸ��'�0�!�G+U�`�qh�yM@��Z��ѢL�L�л\!N�RÕrģફ�;A����R�f�-4E�����֤�����d�C4]%��Џ],�Da��ڜQD��,�|"���4G�y��g`�")R�����CFs^ư�?I�	�笌�G��Yt�CXB{c�1b)�+�iV�^s�)4���"χ&��?;mņ�1(�j���Ê"���X$Lo2!/뭓��0�,؋���Y[<3����(�{�A{N���=��d9KӇD?m+��x��M#絥'`ѭ~W1�{Ǧh.ڛ�����l(d�vv���w�Ѻ��bF)rն>{�_"
��U<}�0��??|�!�\��w��\�;����͋�"� �O�K瓖��F�����uɞ=��T9�#�M�OOiV���TUM4�hl�|4�Lw�`Hc�u,��.�_��λ�"����*w�&��V���-��:��=o���+{�Ο'헪F&_,�����Y|�O��B-�ց`�ø���|�g�/�ÙG ���U�-�9�����?bZ�댟8����~?y�ߤtR�0�?kFǱm��Iq4�[	�����@'���Ci`�d���p��_��:~cXH���Iʇ�u��<V��crA,B�5�$����mS>�!���JI��7.i�=�	"�����-@<1�ZE�{�A[t�9�g���_����j�tǡ�qT�y�֎3��0ԁ?�O�F��h׻[��ʮa/u�y�X��i�'nGTͳ���!�š���tvH��\���OTEV��ѪwA�Uw�^����%@<d��P�e�UO�b��I����x��4
���O�!ڇ�4�	l���.%v]�o�bb�	��$��@$)��\�P��SW�Ӝ����4�rQ��: zūk�K&N*L]�W�jh��iJV�?�o���(��I��t���1R�܄S���Ž�U�}���^�s���iء﹨AЉ������4��-&N	�?W��/�oZ���x�n�9ؓu�pQtL�\�q�˳t��LW�D��Eǝ�I� >0^#;u#ĺ�7�I;&S5���������8
F�P�CҨ#�k"���G.q��[hI�q�V?� gZ� ���(�"��`��ԚvO �e����"�1E؅k�`኏QVLm�#�]��۶HZ���L�?z���Fl'��.��wq�*s�0����t��� ���~�Q
T���!���Y3�ɴ��Y�B-������{�n��[*�(=�����
oPh�_�g�i�cXD=c��7G:���UaP�_<O�81q��Vr`����V{�t�K�
�U�9�����̏��|U,����
E�"�<����] ���Q#_ZD��3�>T���d�A�	Z ���G4�?kmo/��
��)�{p��՞��|Ip�)Q��Kk�@$�|u�l�o_��@����Ub���#Y�U��g2���Vz\�ݒ��z����6�4n�U�	����}C�-�+�=���l�dGB6��QKq/lp�"$�|�Z����uڙP/e�#/=xU�s-�<��w��d�A��)(B������U�^���'�s�u�0%pI`�.�ʎ5`O<��隗�X��1(W�=�b���a䇆aɮ��|�U��.ֺ�J3e��������L֊��g�U�s;�4��0��*fg9���2ϑu�zaY5]U��0�J_�ː��\F8��"Y%gc�@L��p�	�Y�F�L��&:A�vr](E�l:t� �ҿF���~o܎��I����EjV���0�Y���X�5-�	 �Ԏ"�8�k;a�# �lC��Q@rw�F�����K��=�ͧ��pS��"�-Ӄjn��˻�*�<x^i����6�v�+f��4p
A��Sk��.����D�N���5G+ߛ1��l�����qƞ:��ŒlO/�0��'�s�(�:Lj2��'!hW M8��[LO�Ul���T�З�Q�O�-�AS��XY��^'B���Il���<f�~i�N��z�GV��>���xm���U�]RZ���%�U9��b�����{K�g�h���55�Q�b)�b ��$2������ѭ�c�W��A]�]���cK'VL�y���4�C�����'l7������O�$u	�m<x�uY�>�g2�
�B��/��5�t~���T�-ZL>��)�:UW�(N��:y.����Ǒ�-_1�gfl�
mX���3���^�����?���6N���z�m��{��ٚ�[#���G.'s���И�S�"*z`��);J�C0
�@�	��� �;w5��0�4�I��&��+�2u�F�CoQ2�6�I�H,����K����s@z�$	���YAx/a��k�d�Q儞�3ڃ�>j��
��Y3�����CRF�q�Gn��@�q��8� �V�������lWǮ�C�X�8>0Vnr�v��"4�H���[���/8�V1��՞��f�MM�4YW�/+(�J+l�#���M����ߊN�Z�IV�e05�g�R�f�f!ޖ�X��2������x��3�]"����6wd��Z�.�=�)��V2�y�v�萆����l0����t�'�����R���dYv<�0S,`�~��l�Ō�-v��\M�0���箲��.����ܵ
��1��"�]C���_�x��I-�0�R&�����򒊀����,Z��$�S�0[��@_'#���ݚ�Mq�.�h�����w� �o��C�HWR��_������]���K���"����	�@ ��U��A���)���֡K&/ ����鑾T���o1H��0^'A��L����Aԓ�F��C>7� �2v�|=#�f�M���5�Rc�\�9<��w��{�F)u���	���a9lS��bO�tv��W;�e��ǟ�@~�&�����'��
��5��h3�5��Y� �����KL��2`�Qjw�E��r����=$`��|/>A�W�����ώ*�H��Y˟c�O�+��9ȖEU�/�*jx�1�#����.�m�s�r� �3rh�T���s���/�ǎ�ʐF�8�bg�(��]9��˶�G��٦�Ƙn��[1�x�mc�<R��J�\�E�F��vq����2w���h6��7�������8�n�c`5wJ���IF�\�S ON-��:�%�!���q��`��[!N@d�$�F2Br�W��c�zx\��Vd�vc�#B���0˃(i]������9����u4&lS���?����T�(�q�[�.��>5%*۱ vp�u�FKb�����,<�Axذ�Wyu�����ip�?�|YsL ;?l �1B��ĕ
?%������Cd�\IWۖh���}��ȁ�o�ڧ�p�A����5��M�y䆵d}-?t]��'�τ��.��bYk��1Lwu)��:Q��1@�X�ٰ�����O���`.7 ���]���k!�7�Q �nc�&"�p�xr��pK�r��Y���M���;���>�~����`;{�!_�XʊH|Tu_�v��2Y���BdG��w�I�ٓj�[D#����_���E���P���g{�Edv�#�7s^C�/�2��R��A�����j����n[���6D��V&4ҡ�+d�#��{�G�2wG�Q����n*l��5w0�.���8��(J��pX�@X�h%�I�ԧ/�����l]5y�iO-tM�)�X3��ǉlGME��;�U��U�3ch�@.8�q�|�J��1EeUF���:�ϸlM��bR4�,�Zmk��)����'��]ٹv�2�� l+��|�����mej(�hh�Y�^ �3�vM�'�kك��[���&�&e����V_����A�4	�q�;G@���-D�z�3t!l;/i0â���.�dI�c���(���E��P�hӻ8T�۹%�X�vK&L:�� �{X�çu�"V伖�?��Ԛ�?F��\h���nݮ��Y�	>��07�M>|�Z����:�. �PFr��p���F����FF!i�u��P�\�d� �F��^�����9خi��Q�n�;�j.���E^����R����JK$@��gT��$*����gfl/�.��*�����pJ�ǃz���ɴ-̉�,��s�#�9����{��k��ߍeH6�ײb��M��#�P�nG{��~̓p�1و��+����1���GJa���J�����3q$M�/A��u�#� ��^;�����1P��E¯��;���!	+�O��L�k$u�8b�bI1u.��<�w�Zz�vw��W�����j��L����_^/k��b}����D�9@�ч=��Rzi{�^��f-A� �d\�0�脒:j��N�&n"�ڬ6�����c��u�k��&a���F)�%>"��_(���,ڝ��`
�4حS��=�?g(8#�n	a�3NӶ=���,>?|LXkdw§��a�� ag�
V����+V����T�����f��k��i��)�ԩ���=��I��yKH!��a
0P���4R��R34ṅݠ�YA�V�q\Vn�<F�~�kQ��&���z��&����g�n�D�ak���+��`	(��h�����O�n�K<��J���Ap��^N�6��Ξ���&	J����pz�f<�p��
�r�[�j��in�@W
Bw���L�(se7ŁXN�w0{�b�V�A}ŀ/-ㅿhp���:԰w�YđCxZ�{�.���zi��_>U ��;��ډ�e e�!X^DCE!۱�i���G���dX��mw����/2���z�V��脸��!�ύ�y�8�yT��."�
*���Q�9���Y)rn�� �y����}}c�Nlm����H$.��!m�	+��wb��AQ�ι���� ZObגԡ��1��&�E/_���������f�ī-�Sa[�!Ϧ�#ٓ�#���m��c�f�)�T	�_�|'\W�~�Z7�'N�A;DM��=����>hj�$A;��6�H�ztz�u�(�H�HW�HW���z� ���:��D����8�a��O���ߐ��`��W:���.�*�#�;Q;�`�	����h�X����GP�\�j��2M���f��+�˯��	+2���t���.5+p�0�q�6��{�۶�2���|���<��,�L�)�5>�*�tDO	�ad��W��𺹂>w���b  ����+%W*[ǰ�+�՝����}ޅ�C�P�y��v�l�:i�(����l�i�UF��Rp������F�ź��q�y�Ϊ*�R��gr]=m���%���V���K���+j�HҤh?��[p�\ờ�3�(7+9+���?���[�B�#�����J/�B�Ү�����M��N��8ɞY���!�>�xemM��D���P�qFC�P�H@.P��zO�a0�8�Ž�ϊ>l�QI�c؊f��}���KJG�bR������a�������A�����-}��.���ղ�jA�7\����v���.:����Z�����`���S������2W����\,ǀu�w���Qd�񫘌�WF�Iߍ=j�~ف�K�Kɕ�ci��ȸ�W���F�m��t�,Ȉ��L�1��bM��j*��G�l�<N���#.�f�Nr<j��ŵg�+��_䥛a�|����q�YTĕi�2B�J@B�@L��T�O���D
̹����6]k_�L�Y4�!L��1���|�!ŝaT��e��	�v�ew�U��SH��55�*�bU,��Ӟ�o�4U���	�+����h���
	;J����e���b��u��N^�qƪMM�7^����%�B���tL�M���PN*b<XN�̍A׮V�h0	�`t�A�cB�_Y|= �0�ł;ޫ+W4�i�^�e�c��ѥ��zc�w�5���k�h��9�W3!��\������4��Rd�%/`G�q)	s~�N����۾��� �=��lܩ���U,Y���-�����߰��E�%YqZ_q;��d���|�2:�$~�2[����Z�>�P� ��pu(Y9�΀]a�����KqƱf���毿i�A�R�J)� ��o�x���`�p!�rI��%�Q~mc�^��9������ӝ�;�Ѐ�2<+�uU_��4�A�MBx	��p�S�H���i�{~G�E>�V���~�~�>cS\��;��c�W�&��_*i����45JGI����h�}u�CLX<i�? ��~<�C`*L4�:T:{��nĀm�E,��V���~�j��/*4ܢ.��Y��������P6pl�_�ya����qB�}������)m4�[�f��k��H �Љ�O����q�/A�+�	��L	�b��Z>&E��T��N�ϵ�i�'7�4T"5�|����2�Gڿj��ɝ��-��w�!��' }B��޹�����O2�<ڶ{������F�U;��(|��0-�s�cR�(	�������T��D�͋8�}=/v���h��L��1}��e�B�&7��2�豞*;�)�����_Е��aY0l͉8��� Sʛ��\�-�U���Y���EI���F �4�G��;Z�K���*��u�c#�Hߞ������q;Œ�~END�t�����3��̭���#`�<�w"�x~K��s&m��WU���"25YJ]��Ů���?���@���G�1A1I���>~p�0Mf8O�����=�ߢ�|�~�g��#��`�<�)H:E8�дQZ�٧Q>D1.�l�V�H�n�201�+����e��%ML���H~����:�@�o�`��ȏ��+}EH�U#����m���duN��E��$B�#�$��b$����w{na�;��Kx���ߣu��Q���/=L���ߖ��J'�+��$䡩t�#�<�_:Ks\Hj�j@��dU�e��o0��/o���m��({"�#��BM�n��nj@�ȏ�XL6�p��Y�(��nX_�a����5�o6W���E��f��`�H7��.g�\6j��}�+Z�(A����B��t�3���
��:�)�&*�s�D�>�	DN�lD�&^Mb���xkI���?���������g��b��t���|k�����Cjr��|j'd�ʺ����:�'�gSw1{6?ЁUx����ן�۷-��=֬Щ��v<�W�Wo�^���rJ���%��R�4V�}\%ESA=J@׳�DG�J�\���6f�*��~W�_6��5��G�w[��/׏�e�1'�"8���
x��S�hᷗ�Ɯ#z���ԣ ΅84�*I���pFl9z�1�'�o��م�P(�|�o�>����d�S�}�6�-i{�f~�N5��I�~Ll�M�-'�,[��dW�������ոϺEviœ�^�����F鍐o���w!`�:�K�ǥp�\�է��L�.`��^�6[�)d8헚��΂9�Bƨ)>��;����t���x�cµk���l6�8��GZ
Ѹ{˿�� ��%��u&=.�W�dZ�ʵ�W(k"��2-�P7i��	�x�׬�g��G2C�1��7��/��.�ܼBz3��N�!9D ��Ԓ�~I���B����M�'��X�J�Q��t��xi��C�M��	uHS]r�{#0�q��m�ఁ��߳`�V�p���Ac��i�g�i�&Y�}&�u���U�y/���|b��T�2�0�}� �r����u�T-��0�j�WD�Ep�J��P����&�9��ka�<�&�۶&X�{*��X���������ho���]z-m�>�~!�5�`Ɓ;�h��s4�h���˚�F�V����7�ix'���t)�i���ڊi'�o:(8��z�+b�4����	)��rͱ��զ����x�.�N0��[-�3_�c��/�~_���E����|�3��jv3j��Ѻ�Vɕ%���	8q#j?��&�L����u1n�^F= ��ig��E��QV-���3�ga�wd���x�X���ˠ���ׁ���=���s��3/#W�Vo�|lo�)�I����~6��F���?�;+���Kt�}���6���vwi|:��$���f�j	���Ζ���N P�"��^�>�f���+��/�J5e��Ę�t� ���i׉/c��rt	��[�Ь�9/�(��G8��$����z�[�(l�"�XE���Y �
mke�P.����,Ued�F��}�c���&�6���W���HͰ=L����L��7�j��}��O���Ly�-�����~;�����Cj���bص�������48^���������M��	�E=pt��rΈ�-<���I���"�����z���8�'�8�#2/�B��*�AW8e���^���>cZ�g�
?ju9Xm�G�XX�˻S���=�\���@�c� �fp�ќA�m��tX�����e�����(J\��J�%��X���ۮ����4l�c�1�BdI%"�Xt�|�	&�X�/ܒqo>V����oZ-
K�������O6���#�P�t�O����>�9�)Vs~�"��.�Wmb��^=��&($pe��8���$��Y�ԥĿX������ ��n�"f�� ������!{B�'���G���9�.B\�� �,(� ��w�Y����2P�V�{%:M��f���f�M�G��I�s�m'�IMnW�Ĥ�R����- (�C��+�����DkB�N���*M�#�9����B�����M��O�#���^h3�{}A*��2vu#������ѯ�������!��i�T��DI���C�xzf0g��J�_���qv���o89�qq����F�WZC�md�H'���#�g��+W(�s����{՚�DH^���X7P�tF-5!z&���b9��4��0c��L
"I�f2�������ib蜬dy���0�o����5Y�с���'����R�s[�s���%��� ��[��,�������ޮ.����"��,s���ߡ�@�n{'O�M���H��mv�!r|	njǕ~�Ò85TE�)j��IR��<0h�UcD&|v"hU�l�1[�d�$fjV�1��a8l�U��d�c]S���H�.���(��dr�c�j�(�=�e��ߏ�y}�����D��(��m�Kp�p���ز�5�7=\���~�i�M�&tA�k�'R�e���v�-k��wd�fYWr�Y ��Y.>�tӼ�]��R�܁T'ʊsz5�xeGU�
s�����bT��¤iE�� k��͵�r��I�]0M����zw�V/�Avv/��*u������S�x�l����T��Q�[���jLF��$;k�R�r/�1L�u�����v��R�L]����%�-rt�k��ɰ�:U�d�ѱ�,�=�!U}�)v荲��HҰZ ��I
/r"�(��^	8; ���;0=�B�I�={�a_�:b�r���pg<\��yz�t����D@/���K�3cs6`�H+خ�����KqB,ɗ�,���&���}�u�e�hx�h����k�m�8p�:k�K�Ogzn9��) �[#HS��^�~K�����{��Hjm�<�ނ�M��]p�`ۚ�(E�l+�j0.U�b���˽��j�Y�N���f��?���p��W���-�2�$�X�N��r��b��;�%X�ki7g~)_ �1���$�A��B�1�E�Q�~42Q����Q�M���T�9�rZ��L)��ښ��m�����������җ�jt��)zV3k��mfɍT��5'�[��SeB����/�Hڢ�r},�g��e�=niʽ1���x�h����P8/q���40�1���ps:o�=XѢ8g�Apk9��66��-G�*���z+�Ăh��~�_�C��ז:L�=2?V;΂jl���IϞ*������3��b6��PR	.�S�tU--D)?�Hꂖ�<�S{#�����p��s	�م���f�L)�1����O��&����"���R|}�ٱ��g(qKQ������g�4�-�b�>XA-�x����+K`�Y����3�c���*��	�-<� �ڨ!�gE��j��O�G'r}Q������DPK0Y�S�/U@S&�������Yհ&���F^
�2R�?�%�I�4O��>S	�r�D��0 �w0�n��t59��3�>�
! �;_��fd!5����v� �(:�����Z�V�T��kј#�A�&7�����y��2��<�&�R�����[C����d!3�ߝ����v��g`/t����QnW�eF�@3s���!h{ٟ��<���Er�M�" ��{�a�����ѯ2���!�uR7��*��/�OSKO���.V�ۆG���j@$�7��z�*<�[ge����YV �g=���D�3�҄��q�2���^]�V�~h7eL[��W���Op�G��tǱ(�[���Ԋ�M��A�'@�����
�TrIP;�������P��F�1Z��}��zk�I�ve�Ԁ*�f��t۽Bо�k?�un
��憶J�0S����Wog�22���� A�a^��{��� �e"SNۙq��
���;�9��r9��[���5�Z �p �������\��,|�~iE��ʞ��I�/&��&���Sț���w�m=�������<ɏ
�U�N��]��ҀH�ͱKn��ab 羞�E�.FFÁ��� M4�oaN)3�m)��qx��������%��b��"��F��i�H�˸<�����@�Oȏ/2�`�Z�4�����:��Ft[��h͔0�C3�
�=�$�&����yU��mՠ�5����Ϻ}�$���ߒI���np��!y�.��45���|�M�sԐC��b�P),����\/�]Ua���?3�a���}�d<{�p��0!x�����
��dE�JȐ���=s1ّ�P���dmH3�`_�>�S�jG�[��R_��u��r���n�W��;@aǚ�'�̛Vp�T'�j|q�9wV�L@�f�~��v�6��	�:��k78C�tW�8�.t��{��I�S�����Qv-�dk}	r5lP�lK9ͥ����DR}��@Q!#`�ŶX�$����<����6�+,V-�'dBv�s���=Yau
�_���N�#Z�s�����zVx���E|��ѭ�T̊�C�'�H��H�A(c�|���d�'��fi���: ���R�e0/�~�a�"c(K4��K@z���S,ҭ���.!�D a��?q䭂w3��-�9Q��!���1|���n���U��/B���%���|	]��Ф��� ���:Y�������T�
��v�ϋ�S��3��Q���x~��"v�\�����
(	�Nd�o���ذl@�ɹ.��G1vΤ"rI�+���0�?8�5ZL��>�{1"��)K���t��D�0�i���������r��O�u��jy���omY����� ��9�:����,�`���̄ǔ�m��"���������7�W�Y}=Uƹ�����=���߰����Q�d�᜖���`R�`1�{BLuV"�+���<��c�U���撿4T�l<�\t��1l��OH�)�P\f1&����톺�w9����[<�2��:��<��~�0��l�W���jxJ��^����s
��"$����Q!�����y	����jB����8��KN���b7^����@��(�A�r�h"��eX��5���lf���UK�t��=Gv|G�pr�𱥣�MU+V��֋J�ٯ͓J��[kZ籋����5*���:�%�Co8b
b���	�J��$��(�F�����(F;�	�u<4�Drꮜ�����#2�ƫ[k$v�,��ޛM�s����t��>��*ɘ[�������`ϵ
�i#���K�C�y����q�NgV ��D<����@����G�k�L���m_���O*��	�N6ь>l\���_k�d���p���:!mj�o��&����趛���(6d)�P��Q��.�\Xu���7�Y>�CEa�����f_eG,��|�~ta��>[i�'�nl���q� �J�z�l����~�蒩;F]��7�#�v&su��ez���`���A;.��0I��vu������f�6�@(���r�.\?(V��Z$�+l�k �^xw5��.-}�7q=rD�ꞧ��SϮ��.Q��`�pg�t�eq Mk��'��Z��ZY��I@.�C���v��_PPA�7FS��ȎIj�BR}����h��]�U扐�LDd�6?������9_�W;�+�*,9�;�/J�Ũ����|UWI���$�%�䌅�$x&u�ʎZ(����PV��L��o����>��$�}���}�+*R;G�0� �6]���g�a_޾�b�$V�9(eND)�lƛ���0y�d<9����b�+���6��2�i������o�f��3�>��`�:������P>63����$�,~���i���ы��z� tl�]��1�Dۼs���u����7e�e�;�6��CL�:]��Դ$;�1�;���F�Gm���wE_sy��	�5�F�Csj�lC�m�%6�To���2��(ɩ���|F i�{�o���:)9�?R� 53�x86�X�1�/�*��-�ǹ�5vvN9���.�;�p����%�&k�w!�-_�F�Z�� �3���r�|n�VrT�N�P�w�sE�l~ �ݨ*��ӕ��	D`���N���|�=� ��1t}�Lkw-�� ����e�t�[l���qxqj@w_�����P(��A�ܝ�Z{x�ȝ���o)�r�����q��A�)�0P�c�}`�k��Ƙ��j�/�y�oX�ʄ��"U5��͋BF�{>���9N����d输Z#*�$��9���,b��~���3Q\��ЋP��ř�z��lV]f�S�K1�:��VNTᆥ2Xug_1����W�����Xh�[ǐu��(ƀ�1��e��e0���г]����ӻk�"����r��ǁ��w�ǎ��%&B&��A�p$h{�?W/Aq���Q��;,�$;��5X��U���$�������A�0��#�Ƨؾ�����yr}�KV�W*Q�0c �r�0u�N��3��]}X�iXAhf훤����\T,y�	��.�$J�����y���5=�Ĝ�uzh��FIL[���ؼ�>K�I�#Rc�r_����?��<F�>~4|�غ�1��i�KמpnEb؝a����"��'��$��j��b�i&�7�Auv�=W)�.Z���g�˲/��\�$Z�6%he����0T8���wR�/�[�� �i�[��j��0�8�,K���`MO�ơ��|;t����f	�S�"�,��=�hB��������#�ŷ�ol���4sn�!�����;"��W���@$��7���<*~��q;(%�	��Ta?�t8,����� ��K��G��b��ek�ҡ!���V`���`�0To�Ft}�A�I
VՈ14�;9O
{A6h[AN��.U0�'[�P������C��V� L5Z�Wr�O�/����l�|�?R*[����>^z�����Y����F8���X�,�U��Ɛ��n#^��$=EL�L��(�`�Ũ��� �pV�WԺ����dj(�R�ޮV���H-�wr�M1"��t�]U�7b8ސ�.1���Mg�J���pK3��8��\�ӛk
|U|)V)_���W�q{��_�|#p)�re�f��H�m�Q	}�Œ��S�������������֝���hBHE����a?@5�N�����ni��] o�/�Y���ĥ�V�u��_�'	$���EZ�/�{��f]�gL�̆2���k��=kR�##o��F��v̐�'h�Fs�&�7=W^_�k(�8آKs \Fw��$��4zg;�I-Q6����!��wvwj���B�Ho��8$�ҵ �H�2#�:��<V!" �<�'۩	�-�d�Z��K�����ui ��f����6{&,�lJS)�5ԍ��?���{��z���-A�.��c����Z��j���4���7�]�#�	sg=��I��r��L��hh7F��/����nT�#+ӯ��%�nZ�V���z�8~�e6S�䗛��u��}ɫ�c������@�"�7� sMecޏ�E�"������U�q��Ջ��Ǹ5*��>��aa�������Q����7�z�b�<��C�+{��e%����t��^%׬b?'��r4��R�L52Dg�.�UE�@5g9xm/����v�#Fs�{M��G��'V��g��G����q�L�ʯx_ȮS��v���xK�D4f�+ wH��A�܅��b5���%��T1�0�W�ޑ���R�KK7��_q�і�]���馌�O���CH�]Y�;�d����<3�]E�a���+Sd7$��/?=?4��4��\ƿS"bE��Dde����E��Oܐ�OE0����K4r�cs'����U�;0iRc$q^�@`�E���8��f��*F悖���iu�����{Ŭ���3�p�hh͸���k4�S�->�yFM+�����m�� �$���@�Q![�r@ί�?�+$�R���f}��MrF�i��ZV�Y���NC��H����Uڸ���v��k�ڣ��3�H����1)��$���>{��x�SH<-�~�ج���b-�H*r�c����Mh5�a�����Q^3�HP@"��D�bB2�;�,�3b�h�����SNQ�ü�Zy�fE"0u�>*���
��X�3!_�j�ƀ��z(�_��8�+�bp�YP��n&������;PFBf10�nDA�R9N��#��t��Yy��F71EA,�\�U�g�/XEI���Y�ϴc���붹����,�x��� _b�����C�d�P$T��+kq�:�hU%�9��|,�h�#zy��6��s���H�O�
�Y��$�V�[E'��[��������)�D줏S�~��<�w�l�ED�s,�8����2p9��	��*��^c_Ȇ��\f��"S�/���+xb^QF[�(�` �9*��5�<���@�M��
�B�`�qҵ�e<������M����-� ��~���F���Pݷ�;�d���Q�V:�ō�ǗF�.O����St4���4͚���B�j>Je��y��f��Y�|ˈA��1R��GE�����Ce�x�H���7�{1,�F,e�EQ��~��[�X�1C�����=È[m�%sV�GT�ف��(B��#�Nz�i�A�-M���|�9����
�� ��DS��9��>R^3��~f>���kO`�v�/R�In��A 葬�����;�h����*��s����M�=��1��
�������
�c���17��0]�m�[@d���6�P�oz��nj��:���	Vͬ�2�t}}�'Yſ~�
��%96��:�n�0�&���U�U����W-��.�_�}*mֆ��&�q6��@V��Lo  �\�QU�����A?ȁ]��2JءJ������F��q/7b���yHXg�ޙ�5DK�T�2=j���0LYA�+�7݀����������U���lR|��
{_����*�~Q#Y�t`<�*j��	l�հ�$Z�,w�	S`�
�+)��$Ex��~^�(U* c)׫
u�N����nk&2q��NVξ�/�y� �,��U�7��|��^YI���p96)3߂����d�D>Ѩ�V��	ק�M
lc@5ּ�����?	���3���.��/H��%���H |���N��_��{��:��k��A넚/�w!��������H�����B�7�z�xz�N��8�n|�0�L:�|�)&6P�C�1�M�z�B���z~S.�e�6���MΒ#,K1Q��0/���# *,-Jo��5��%d*�mA��nԶ�[Q�pt�FA�����
�%�m�j��Q���ٮ��
����S�ˁ.ޮ۶/�`XR�~>�'��r�7�:o*S�&h%��*�+~*W%��y8K��	s�:�?��@j��p��*~����#��]��>K������fH�鶍W��D�I��v�^�ƚ�;A�`D�{?�x2jм��ھ���9���É�ҥ�Ӝ�0N�,U��Z�
i���"�'/��g���gXxԻ6���b	Eh����`�uz��kV�kj�#�H�������N��H}���J�Cegb���&%��������69`�R����"'$��;��:��B3�)����C�(ի1����` ���$��JMlZ5�*��AI�� 
:�)Ȝޙ�E�����#L��M+h#�S�ؽI�/�rp,B9�{8������j&Y�k	�8�B ����S�)�B	#�7�K.?��x�߉��xk+�D�M��i�F�chgR�1g��9w�X}�1����
�#2��L�2_�0�\dNE�桓�	N��V�5�]y��;���I{fr�Mǵ������6n�V��Dɼ�Pc����{�'��E���õ�]���=\ږZ���0&}p	w--M~@-��gQh�f�cU0������G�m�ҡ�esЁ �=�֦�OZ�kl�#��qߤQ�?m>���~܋���F(A�fC��m4`�XZ�&K����I>�����}aC�����3�+W��*M�v��ZN]��fӇ���@hX�����7�������'��Dp>fF?�}G���s�u��u�$�A��#��� \U-;�Z=��󈑂��	�sf��]��go{TM����>���}r���lZOqw���sP�4q���Z���H?���וj����;��BԞ/5F E�ql�hs��S��k���E%����kWZN��@	��X�&v`X��c�k��OZ���2�M�܇u0�ʞ6���:����b�]�)Bo���Qe�#%���j���|%� �q��~�WQ��$�._��%)`D`tj���)k��	���'�~Óz��v�-���PVm�9�V�M{����ճ]��w-sȞ��y��|�Љ��_��ɱ�]~��x�+�S��?�!y;�5' '�Aa��g�$���+;_�x���e�������=�n����$�����M�Hg)�e����'�5��3�k(��v��%oTp��%��DuW��|��:��%&6�#�B|G%N�P��|�w��<�{тO�S�����~��[V#�K� ��"����e�Z?4�[-���\`d�a��Iu�L{�W������	�tf5�!�REf�S��A�T�\���Q��D����.4Am���v�$6T+��g��<��ڔ N�`j�Y9�>�4ԥ3��V��U�Z6W����&F"��T+lD}c����Nn "'�[��	�����ϒ���+0k$�ʀ{#�Fh�J��w��}_�.j~mA�z��Ba�D�,�y<S����o�2TMI|l5\)��gߵ��{L	=-�kj��q����ʹVƄ0A�
 �ŬN�7�"6@ޑ���a�/�X8S(m�)�3�Q!ɬ��:q8ΰ�d����L�\� �����b�ޗ-/f��%3����}�4��K�;����\:� u�{�[m�i�j��'�=N2�0E�?�5�r7��OJ��Ӱ�ܳ�l���Z�n�@��Е&�p�D��.4�����3k�r��.>_H?���� ��SрˆΔ]���MT5���ngM��e�m!砗����0��������A��GJ��z��Bڭ��+W7��\���>#�<JO���4�5�>�).�FOi��^9�gR����1m&+XW��{��F��Y�jڭ�E,L��@�j����4Mph�O���jv�+i������e�VqC-n�γ��zQ�D�!y97A���gp��\+�:���o�q��m��v zF��ᗤY�٭f��b�Ln����JE�-,��!�S	��h!!}��� ��^�ˊ��浰~k������8`z�č0�e(+��IJ�Y������ ��Jfa��r5�)B��SPh���cPB�G<���w86>���85	�c��z���J�y�%��5MnU)���?�Uv�[���Da������0�5�kØY�r�|�����2}2�#��9X)��V��b��R_�rb�y{��U��|�Wۂͻ���3}�����G��W��R&��Fbf�G����XS�a��u;(����l6����H�,ؚ�:�˿t9i�URt� Y��CD���0?��%4�d"��q!ɝJS�1眩���2Q�`���vF��k���=?w���ѭ�������⪱OjΕà�o/��}�	���� ���\�z:�7��h8"���<w9"��֧���- �~�K��Z|R�Yu������1���;jKw�/e�`�Ului5�րit���p�OZ�X���10!+�9TZ幛;ԁ�E���r��P/�Jߏ���׫?3�c�ݴ�a(�g����B�y���9�b�7�lk����F�|z�KcV�����E.��!{�,���:��>v=�L����xҽ�Hۧ�l�0���P �%dHf `��u̽�_��2fD�t��V@��+�\�o�$�(~p�4���M�>^�O�#��Q;��ºf�8k�K���;�冥���'�FV@R�'�����\l+�*/D�ZZ����bٛ���o�{RI��_L���a2��w��I�f�
�����O�РH�^�^��-汃�e��&-�y��ALƋ�|��%*ЅK�{�	ȬPFg< @�;�u	�΢�5�W�V�؇�����X-	P����%O4�CW�Mz����{|kC˩\Q�n*��+1��3��M���`q��e16N!�!M�{4�Pl�j����SH�pY�R�ʉ?u�� R�e'%�xdL�&�����T�.<�-��!H9X��iF���]�5�b߆�y��T��C}�b��)|M�'�n��x��t��d�f����|v���<��$�2�<�Pn�z�W^��CN$MP�ޫ2�3:>�������^Hl��KJ�T�Nbܼ2\�I��y��约ϞWM>��O��l�5�u�b���̚~,�p��`�;��B��/]�;����`�﹏�{�Z��'�"ZN@X�ۼy%/��:Rg�2�Jf0d���Q-@l�;�	�[< u��Z�+X���B˾��Ǹwj�dl\QZދ>Jܒ�.9�.��E	C���]��Q���,�2�����Mp�=��dEh�fL���cH�Xֱk�{�
<���g�0��g�I@S)��_A~�@qfWnsf<Δ���R��Yʄ(m� �~�yq?$�*�6��ZZl�/�[\�@SD:��Z�?�:ơ׊�f�H%MQ���h��zfez�i�!�)�*'C���)����0�{�.��[�Ɨmm��_�p�h��_'4�[�.���6��t7-��+�*΂�fk[�96�jt�8�́\k��4qRdA��e%6����E�u����"J�2��J�pZ������\�s7����J�c�c��-v���mr@z�'�5�<���D${\�{BR�)�~|�����7X$Q�_�?l�����RB�e�ʵ��1��gT�U�;�䆙�M{7k��ZY�A����N����Qj�Q��teܢá��\��	g��\��k3�
i�ż<��L��o�ٲ)^�}�/V���*CΌ0??d �j�0=�z����
+;0��$\Re�<�i����҂�x���6+�I�!z�>>?���us�"���(r��g*GO��q��'u��c�,'6�a~?�r�k��K|j"�|�\D��2���C	5t.�H}ɼ�����.��z�\ǑO��^�n+��"8��=�6@�0YY�gbR�5�ҝ
D�)�� ?u7b����d2G��oL����h��?Lfɑ�7�X$��\�? 28t���N�BP�q8�X*�<��!~���:E���`��~R0�,Q;��ߍU�vwc�?Ԍ�6���LL����(�K%QDjs,�v{~�o"՗���c����v��g�����~���J��ɽ�+��p��>U�f<��� ��I�R��F���]�=2O�C�d�'H0V�P�ھ�D�����I��5Y���N����,1n�J�XuY�6!�k�C�5Z�J��`r�����̤�Y>����W��њ"K�(Y ����9K��t\��1v�7�Q�N���Q��*�Ӟo����<�^-̪�/��kɄe	�a���43����'�y�����b󣹱��ڹgr ͩD����q���i�@B۔�W�t���[�&c�j���(�f�"�~54Q��[@��`1��\����1������#~4f��N���+G��AE�	�ȫ���[�~�^� ͣ�zq�jѥ�����B���]�m@7<�3�z=�	�d4��8�ơBkb���c�.1���ݜ�F)�=�����]R����i�+s=�F_��8����S����7:2J�m��K+V��LV�Kw&+߰jG	�И�7����Vr+��@d��],�}0V[,I���u�L�Ƹ��P���az�aN�O� �j����N�	�þ�'t��N�f�̈��~�� ]��٤q:B�C��c��NGH	��b����]I���d�2���p�֌�>����#%٬&6UZ�`I�L�_�����U�F"���2z�&��N������O\WgM^�l�'��^b}o���J�j��l69
�D闹��*0ét�y-�?�h�Cy��M��9bҪ�θd#|�������5����X��q��L�iC�k�da��������/�%�`��2��O���;�78�o�V�L���t�V��[?��^�H���(�aӘ��M~�s�#tu%ݠyڻ�KZB�m���?p{�Mm�����u �����J���l�S^Ǥ���0<Mǘ:M��Pd�P�]����5�ek��V��*T�����ϣԽ�V�n��&���[����MF2I�����G��	q�����n�����t�X�j�w��e�����;��%���\��$�X�\���y��/��Ds��bLU ;�d�d�%�=ML{������Q|�;MɆ�>��r7��]E��F��f��_cY���z9V�*����7y����'��F�n�2��]�2�ri�ٷ^N��YP���+�ɸ�NM˺[�"�|[(��RUuذ�z�G���Hޡ&m�\��F��FXn�P��"�0��}մbl��}Hھl��S��¢�*�\1�:��R�\�i�u6�Q:f����dew#�ٰ
���4�h�͍�r�s'bg]��d�[�Pnv��3����������@�ko�f/����A�?�1�@}����U��T��J󒫮��j~y%/���6��.��Er�ˠĤb�K�u��e���i�)��g�
;�&f������%�k����t��)�!l�9�M7�<{b>�
�nez1����5�uq����>Y_���곑r�Ѻ��TgT��Y!���;��By�ᛱE��//SZ�}����4M����ɉǸ+.���N�^��J��ˏR����A��RoЖQ\�j�x�Ϝ�_�s�R6��U��AKG�"H^��#�(uӖ�׶�Ӳ5E� 'we�?��In`Xu}LىM�����σ�����w�H��B�v�o���@�� ��2��]�����pF�˺%s�z>�������yr(7�w�8�L؞��m cIl���]!��Hosi}y����lPM�\����^�YR�%�O����)�v�M��==�`ʘE����rɒ�ݑx}U���:�[o8�|�)���v��ʔ�TK_k"��2¥஍K�eH��`ͣ��]mJ��!hJbf��O�ꩭ6�j�	�(c��9YV^��V�@:8��'ݩ늕0���l��Dsi������5:Fn�o[��E��3l���p>�)�f�5�ƃ-,^R��h�W�)(��B�ilpE�TSBl��H�`Ԓ�$4�>���e�/�پ����P�o#�\�*`�G��Qr
T0��_��Z�K���n:��+>`@c\C�-ee��9�͵0�a�j� _l��&y_s_/B� �v]����z&»�<�W� r�������4������+���Z���/�
��"]�#�P�ru��~+	����u�+��j=�>����m�5�t�7D� ���D�d����.�G��u6c�MN��m*��cN��թ��[�����5��9����Ǫm�������������Up���Nv�,N�j�R�"���`.�cC�	���d��!��O��F��m��ЅmN�����<�J0|L�^�]�ӆ���D���[S���]��H�9��j`�Q�� �s8�o��OW�e.l� ��j�U����޹j,7�5�TbO����N��b���I�(��\�{:[M���+-��Ւ�A#�L��?F3����u�%
h�.<�K)��~�^��_
p�3�ܟ��u�҅��1�2C�	ln�dcA-ۻ_�Ɗ��� k�K�ĝҎ�U*r��v�=s����P�(�Ueu�������  ��}�"�W�[{h��N�S>����]�p�8E��hC@��N˩&��~f���y�d&��d�<WE_�}D��]9��H��\�!]�b�����޼��^�=���8�/���������t���O
%����{Ъ��Q�
'	kP����o5>Mh��6�茣��U?繕� ?q��q� ;�#C>�k�qw1��Ol�{��;7'x�P�+�΋Ex�lQ`<#B$G��l���AJ�-���,�Cp���aV<O���\��!I@�^�r�+$8��'�Wf_rq�嗛V/>�����һ��}�5�		�t�4ⱦ{a^�O��{]H՗ȱ�{�ev��Տ�D�0�-��������m@�3�~�3�a���ɝ�˄Of�r�[�C~jj��.u�9�ȯ2�u���!ӄ��/�Č03��Z�w
�(���9n� �hfh&0i��|�C��ɘ�Zk	u|E.��u�������+ow:�"�綑����U�;��$<���r��%����������K�HB����%�pK���KT溹^bR���W��'�Ҧ޵�m��(Ot�N��d����\}-;φ����T���+s��%����_��Gj��U�_���b����i��v�z�c2Ϭ�����F�>N.�vZrt�ƛ�Q [W���D����g���D�-�q\�����'0O�Ń>���`�GF�#QPĽ��kqб��̐���d:��u��ߟp(��,���uZ���_��?�V9����9�Iֶ Y�w��c\m�x?�	��#�f%DW.f,�svP	-򴋶E���?�ls�������Uו���>2r�]*�^��q�<E�s��H�x�+Se���G3fʬ����5�Otu���E9������R����Vm�	�
�4,�� ���ۼ@�|��[y�S�X�����:�k��Yh��X�S�-�$��ix@I�K��v�8���TE=0Eo&��9;A-\�m k����*�&�	��+�*ӗA4�ڝ�F��~��ˇH����̘���K�I��K�PT5�����ʯ �}4w�R�{��k+v�/��.��oD�6Vر�nԴ8��?|���O\��Q��ٓIn,� ���}Y+��eߡAppa�F�F�����0��S��� Ǟ�x����JMr/�QhJyѫ�mx��#�4]b'��@�e��{�q"��}�iJ��KB��@��5a)��+���y�j�oZ˄+��:y<�̖[q˴�T��)C�RK}~^���ɥ�oL|�?1�JX�W_V\���:]�_c!������(�Qښ�3�������-�HR4�a�~c(��	��Ŷ��u7m�f�{����UGt� �Y��h=�3������3 �68Y]:�
W "����'o�K�������a�b{�`��$�8�价B��b�y,h@m-T�O���3k�"�uE�9 ��ڍ�RE\���4�sc��0���M�39�wb�Tt���j��-V6�
6K��Z7���p�C�n�OU�m<�������ߙ臓<��z��aT�F-݁B�d�� ��������i�����j�샻ic�q�>��ͪ�����7�5�)&����z���}���{�K�����i��?(�Vtr��������6^�Xd@MK����yG��"ϓB�qX���9�N�y͔�j����ۜ����O_-CƔڒ�����i�P,�"L4'�6��H���hg��)��b�<2�^��>��ōg�,IL4�}��G�ѻ���'c��F��
��S�9v���{o%��;��K�,䶁�4	��p��-�=����HYS�3���[8F��5�8WQ�����&�΀$0 cdϨ7�:#8x��$ـ��v��h�d"�ًxxa)i�t��+]�x�hC���a"�_��4��^�q4b�g��ʵ�\B�#ǐ#{��?�����ϴ�q��{���=�7��^���0�y���-&�����f)ӥc����\<��P�uEyr��Bp��
����ة�d�]#{��n�����ј��	t ���G�!���v%;u�!�!65総r��d��Aql���������b���9��=�3����}�LN��t�X�J��w�ÿJ�����8����UO�e�Mi��Pk�lCT#t3]�;�Xx�d:���y�'�cF:,J��O�2Y���g���H�`)��t�
�ug��%��Y��25�
`�d@%E��B��Q�vD���TX�ս��Qw�A{dػ᱋ܖp��Ű� C��剾L���6��.�x{ehp�ʠ'��\	A0"��[��,�Q�zuD��١��-%�f�|��$�ɍ��|����BĻ.�~G?����b��@�y{Z�1&�Z���1{K`g���(��
=p�4G�H�&��$[��/�T��|��ݿ����������< 
0�����H �Âˁv���O���O�ˑh�O���wJB
/�#� �����w�����u�i�h{"�t*�p<��5�7dav}Pcg%��۞J<Fr���|��D���M�¦���
�bR?��� ���2ٳ@*Л@�pGȃp�g��������'�Ue�U����5w14�,Ub�^p}&��5�+qpT9��a�]�\4)}��
a��Wl0���9x #�Z��n �^*�C�����%��o�/��RSKb���Ԡ�����By��nKʭ\�Y����b%�Mn,�,Ҝ�`�W�T*Mg)B��[M�Yf��L�)�d!	}�g�\�2[�4'��d�є��?8��m�	jM�!LB$-v�1��D��Z�JL�T ���b$熋�@+|�l+��HH�G�2�n�f�=TJ�ȝ�Azb�����VR��e��~�x��v<��ǆ D$��I��!Ӹ����ߚ�z7����Fw�ch����$�M�T��P�+G��b�1�¥�vmɲ�l���w����SH�3�[ぃ�g�m|찍C�N�B~���	�x�Q��}�h�2�aط谝|�{��X&��Qh�Zք�s�����n'�ɾع$8 �w����4)W�3]E�� �B��	;��ea�c�N�����/��>������5�;^%�Q	y��&|��G�,禒%�����;�ʙ!�R#��]���
���M#�{h� ��ল�*�r�4�#o W��'T�e"�w��b��b,�$Q�e�n����sNy��l���Q5
�n{Č�&T�5��r���y��p0"�Q����b�˩;�Y�(h�4�[�����wp�	�Ql�C?�(�\G�֖�U�p6�� ���`�����'�z|��!�����-�s�U�U2�JK��Avn�n��8M�7B�onh�.��mZ��c�ra�E��o@ �wA�D�p�͗j��/1�^��m�PcX��G�2�<FĹ���O�r��4>짃��4�h�0���һ��PL���A
�w7|f^���0
��$��s5��e�;C/�#�@��ܠ�U��O�d���Ir��Iǳ��Z�H���g�H�"��3&�v\}c/	1���l���L�L;_	�DA���⽋J�=��i�kp�3<1�� ��^<	�P<�"/Q��E��Ѳ�C�{�u>���r���G�����,�iV�/ɬ�n��[���c�(}���,	�6�6r��Nu0�TmiϡhV���L9���@ц]��%������E�gi�I;֢������=i��{g�[9��XӜ*.K�UUi�>g@@�Q ���������f�0���u5�����ɣ܏�C�U�������)T��s�{Zb�C��fX�m��9��:�k�!�6��)W�"�Dx4��rA�K�?]B�U$���g���� ��_���*�(_�hBGV�E��ڝ�0�Q�iFN��f�Чy��L��n����
�`{���±9K�F�T�"�}p ��G�g��;��=�@�������6X`���E�"��! �\��m�C�;Bc�$�k��=]��Y۰0���D$�)7G�#1Ђ��\'�	2H)Čyd�2Ih}�q�ޢ$B�/D�A{I����db7V�<|��pRb�<���ǳ�/:���m�Ҭ�u�;��q	VC=B�LfWC�TE࿰��>]���z=�:�4�D��jtjk���Tl[1�u�i���.�ļ�� ��Һ|7j!D��7���}b36�.�Л�ק��ܥA:�-�8�;�	S�����&�g�	�Yp2�DD`�B�b���	TG���4y7���mu@7����R�4�H�����c�q(e+�Q�h�X@=s���|��> ��w{�^���
5����梋�m�p�)���3S/f.=u���OJJnߥ�Ɍ:r_�jL
���1�S���Q.{V��L�ش~�K��q�Cs��c���l�[�b���׎��-hȔ���W��t�wCR;^�/���,Y�Q��9�Xh���	����N՝`�7��M�KV�W���y���4�4z��Uۤ������ڇ���7�R�%�L<�o!-+ �)-�ʑj��K���-��@٠�����lcG�-@�{I�[��z�uE����c�l�{kEG̝�����[�E�/����S�`a�����[ʞq�%E�,֣��&I)Mj��wI� M��W�8Ȇds𳷆�2�V"����Ǜ1�gWL�BmX������X8�)��o���T���	Xar�t�	��C�Y�ݏ��	�U�X�s�{o~����`/Ⱦ�2��B�q6~�PGU_��&- #/4f[ID��߸�@�Y�.���xW���,]a5Np~�|0��OEũ����߀�����I�@P����-y�ZX��w�����������(�4}X��RG%��eA�N0=D�b�#+�`6�ZA*W{+3��!9�a�N��͇M�<kbd�I�h��iރ'ݍɞ��"��w�8�1E�@��e����-�66eO_���ç8�L3���ml��)Sn·xV/����nHv;�|��F���@�N��썐��?ܼ<�H��>⟘�F�p'�r��\l���[�n���,�"��g��<$B)пC=�B���9���������7=3+�i� 	O��H��1������bXٻ�y��/�d��x}���,�I'$k,񪳦��	ļwטx����z����aD�ׅ�#���{ Ö}�.)D�܊�>��Q���S,.w�F^�QV����c� ��fY�M������R���x()�,�SdW���zs�_=���������4��{��4 �&Xꪍ��j�������'T�w),S��$��0�缋1��MVG��[����5���]H�VPAx�]�&����˶�Ďk�5?�&�����̉NVv�\�c��3
꾫F�.1�σ��Wߕ;��X7dI�*e�;��OrW=�w�~���2H��$Ȣآ��򯯹�3A�B^��˞}݅���R#%�uڌ�=9;;��7%_���g�ΆW����4�����N���8���BH�G�l6���r� Se�bYbo_�?��~E���zl�r��tH}VLMM�JB�����XIY��m-<�?=e��{�K�U�ݤ�j,�Dnk��XD��:��1A�OF��S�M+����)p�p(���3�c$Ll�|�3�+�!�z�M��t�K)�!:��E-$����}J�p����k�J/��e��iK��{[s��jҡ>Uz�=�����^"6��2�����Em���1A6��$���N'���b��1�{%�}�?#n.>�e߮���3�.���jkg�~N�
x�r���#I����xx��1Ԭ�󁦱N�FO2d��j:���"�#o���3�� \�A2�g{������}Z5h.�R�0�hT��v;�p�C��95�1K� �~�~�'0��{
�ڈ��ƀY.��_�,�h/�@%@2���g�\�d�����#�k��<G�}Mf�%�$�y����U�Mg�6������СG�Dy��� �﷔֨,"GP2�ڮ]IdSm;X��2G������J�Fx�:J�� /Fs	�#T2��f⁡���-�����&j)`�#�G12��i�H�e1���&���(�B��v��;��b$~X���߄���ٛddH� ��l�-mO�jѵ)���H��P�7U0r�Q][e�nҏj��]3�'��(�¥�-��1�*�X*f��A��Q��l�k�6qL0)}b�aIOiTg<�If<%tD�)����c'�k�Yy��*�sY��f������V��Ƅ�+}�K�+�d��ye����ń��D�J�Bթ�=�ʹtU{�mDV�K���sf��`Ǎ$[��av#�,�g�U�18��գDi���������~ۆ4��L	��s�h$�+x��?����0I*�s>t��SA���v*�ջ�?8��o+H	U��|�)���8U�hґ��y�C���d_��ސ� �k��|SE{�
�ԣ��u��![� ��d��k1�L̮�X!�ɤ0O�5Ӆt�l�INp*�*����i%'���tS�uơE��x�:�(,]HS�n������Ke�*�'�n�$�c�d�u$��:��u�I;�d�^p��fE)��3�6��j2��O�?[��g��=W�I��~�2��$���GHQL��Q���د����0�U+���O� �~���q	X*<��#�"����5��U�f���%�Z�u���H^�.��y+s���{(�e�0@���t,�����cK��can�#u�P3�+
1Dw�WC��ݐE��d�c��l
o�,�q�:¢�P��T+���I��|C��}*ȥ2�.I�y�J"d}/!����n��X�e�.U��z��ͦ  ��
q�SPǶ��s�;�@}����ûD+��sim�����aX���gK=c�Ǚ�<�ֲ��X��@�t,Bт%��C�רj������Ȅ��p�a:�}I��=�v�,7�T�J�]*��>*.�K� �N���e�s�G|�����Lp�� ���.����l�O�ݟ�C��ƈ�W��G���9��y)������EK���G��2���D����e	i���d�v9(�¤�wsogr
�t!G���"W�Ts���/�)�u��tؚ	Uy-N��egv�/P�c�6�Ɏ�0�a\@b��~I��!޸؟�r�e��|����ש��H΢1��I�5Y�ϲT�@��Ǩz�� ���f�:c{�٠�	�?Au7�0��{1Gc���>[����,��M,�*�;���_ވ����i�|��mK�F�S����%|3�RO�V-zd�:�W�<Bo�9��Z�V�Nd}�*)/�BrL2�o�c�Aͺ�E���@5���G�VW>)��P���HvS#����+��9�y�U1q��P����
^'H��c-ڋ	-C�s��S���W�{�~1����`�j"hV��[����H�/>��ɸ�l��v?��$9N]$/`���@������Z�H��O8H������`\��ҫ���:$�T��(bl�Iq���5�Å*��y{�D�|�\�=���|�[�{~\��*1�2���XNV6j�%O���y52�4�\;Y�t��p���&"6�����~o���Ryy��@@[�ފ������N|�5]�>K��#�P4oyɐA�V�Rp���l5����4|������/���a<��RT�Q���ۜt�{�9�T�<�LV0+m��Yh��M9� �"���t��ɧ KE�b����K~M�n����_�z8���v��v��Ch�&�b� �
|��h����p�!m4��]�I�7����(S�{�{9R'ko�i�n�A~p�p	���5"<dӺ���-��'�Z�B�`om3�Jb�vڊ�Qg�����x���i��iq	vSZR@��YT֏��\I{i�5�o_��mE��ǔB^8������ֱJ�p=�Lh��AZW|�K��Q$0`���`�������zz���6vP`� 	��z.b��;�ϝUJ�5[w���]M��PBnr{�D�\;s��Uw!_Ly��W�r������|\;o�kQ��N�-��a���o��>+HPIf�����!G���`�:���c�=٢��C��h��q�x�	ۮ
+]P~�{h-K똙*ڷ�Wۉ��5�S�0��2���?�򱐂�&�b�-��j��u���5�������2N�H�l%|���P�^o@�4��,��c�O��j���fs���3���M��!�A�;�pVm�����N�a�C7�p�7����\��u�X�R^�*�_:�N���sҹ+�~��_���5�<a�7�R�.wc��~�L��ۚSx:����)�d��EPY�ZR�_]�^P�l�Mg�w�L��W�V�n�Q�$�9A�Q���$.'�@6��A?#��SB�]�
���+�a���Ԉ����ZK������7���<#N{m)Rq��qBXs0	\��9�]�
�x{|M��- 	���lA^�r2w�_f�`�:{hF�~��>j�`��nv[4�)B��-,�YM����$F���va�)��B,r�k��$��)_g@N�e��}��w���`���+>7��R����a�����g5�b�$��Y�CW���;c���]ثL���'΃Cp���N�3�oAwz���y�M@�g���e�S���,�Z��(��"��!ȵ���f�+������x�"J#?Gg�a�"ư�(�}�'ٺ�
G7	�2��A|r��d2[=���_�B��P&ȡQĜ��ٞa���ʭQѽÜǁ��\VAW"�D�8�,z�MoD�$B�7Y<�
@�4O����G���Ib?}B\��|�d>w��U��:�R�w:{T�} 7:���R�n�����������xڣ�L�=�^f� ���������Y�&���ͽ���+%�0�+�0-g� 5Z]u�d�A&�E:��~(z�qY�Q�m�K7Bl�<�~BG_���(Ә���5�QN���"��iͽ<S�0A`�( ;X�+f�������h�=(��Qݮ����*��5��ٶT<�����ܖ���|�r�w��z3��,Hb�j�w�K�!L��w��71�����ɱ(���a��|���B��M��X�Mg��u�ٹ?�ߘʪ)�c�i[��/F}\�:ĭ���K)fy:2���]��h\:a�2�<���r�=(]��%@3��+?�����PM���G�x�U��XJ��#�h�A/����!�T�/�K&찇¥���)m��-Z  �qDT��f�k��"&H���g�M���Xj��D���� ���`�l���`�yQH}�1���v�y���hرfI|3�-�����3r�`���5���F��SՇ�J5�M1
%���T2J��pcqe<��5��н��N����b�έ���l�-�vs���r�6O^��W&�Dq/��s�Bo�Sa�vf6w2��[����??�R�� �A���%b���w/m ��('�D}�:���i�c��a��X~���vj>��+'�9M)P ���'��.�8n�Rot�i��V�	/�i��1aBdR'���Eɱ�>���#k��fg��dQ������V;oLM��םK���9DQ3��1���WF�<+N�8�/o�ˋQ3�B^�����*1����Q\�?Pp��������A	��չ���H�T��}�x�>���U��l��M#�im��]��^�;������������S/l���!Br�F�9mD��"�&���I+��w+�8WJ�gF4Nq����=>�2a����~��� P6g�Eˤ��=RA�1�@vWk���ܩض�l;���k=k{۩[��Rs]٭r�Oo�L�_\�i�|����|!�fm/��6k�GD�G� A�l	y��|�Z�M=���pSR���E\Ǉ��L�)���G�e��A!���2ո��B�4�a��P�\�4P���Ƽ��	S�<%�&��;z��F�j�C�印�����f3�d-��`�h���?K�fy˻��rJCwd�Ք�y9�s	z���Z�#s�ܸm��-Q*EݲG�}�wj����Nh�m�K)�%  ��k���i�X%��E�����5�?CL^r���0���t [1d���
�_kr�������(�I�^�����㩈�҉ߛ�гS���Y�����R൘��ӆ�б<���_sqVas6DE���?�"���)�(�f�Ɔ�`~�@p��i���p��4�$w����Y\n�ԫ���"W�=1�|1�㈾�\+�	�h]jK��"6�w���S�ݬe1NG���2�]�u��8���x�{���7�=�{��?�Ԇ��(��F��U�\�#���yҒ���ؖ��f��������8S$�{�E��M'd���p���&��ZO�G���w[�S��H����zƜ��>��w	DAo���~vfȥy[����o\t8��	O���9���{pW�r��o�.V�7�6�p�0����3��Ԕ}]%�O[�@"�x,�bB��zr�+qc>BF������N�ݳ�bUl�z��q�dj��n�j��?#஛υ���x��/;GY$V�����<���J$��B'7R��%�I��,��������<Z|�M��qr�������q�J+�p	�e#Ш��N�� ����~Ħ*��-�,��ݓO�萃� ��yl�- 
����;8�n����lH��`EG����;���ݟa"n%�@�4II ���&`��N����]�u�k�(�����`�W�L�ρ��n��~�V&Q�޷�J��xIr�
����q���G2�p�#�Ej3���ˏ�ӹ'$���",��j�U�ư¦�Xħir�)�i�́j[mX�����J���|���	&L�Gz�\�6%�p���Q�U^�@��]59S���~�O����/���=' 3�vO����av�@tR$&_���'�8��}�P�Q�i��l�ot~��D=��5v �j�5�3®���)A`sQ��=�	9�ߌ�G���h��}��B��/6�&2��*&�<�1�����ì,X���	ٓ%��TgOo�����>4�´�z�f�C�P����S � m�=ƛ��?+��q�b'�X�pp:楬�n�(�|���2���vl���ɲ���c9_��t:�y>�v��I�iK&c���Z�=֏��/�Y���� ��'�q�z�yQ��m))��fg	a��f�j���g?����nV����F�[K��Y�}U�hi�P�:0{��lͫI}Ғh�`G�h�@v-���Z'�� ���W�NC�=��8�c�ALo��"�(h�ϓ��]�{�GL��K�����JT�Z��Im ee�"�ಘ����A�Jc��%?O�|T���dYa���:u4�`8D/�LPS����w;���Z��W{M���z��0ş,~���� �o#v���).=���TJc���K�O�����Yn ZS6[cw��b<�:��<�u�=�ig��8�j���� ���f�w�O��cN�==��G> �J5ou�pF-��l��`RL$��V-r�Aw��V~�z۪�W+�ƍH�ѝ�18뒈��S�a���
^�}�G�ް��Mo�V�7���^C���1	��DK�W)=�U�յ\j��[��*��Mr����m�+4�D�X�}ª5m2C����$�q���f��?��s�evط���l�W�N�ɐ�_�����Sb�di��1��}�������礊�d�����ð� �s2��%���o� �zXaf���� �������Sa!V�?�}���k�&̢�*�O��f#��)W^?+�3<��w����j�5g=��o���BMmV�9��`�A���:i��B���|�I�}`%˥�0]\ZD]n �L�V����/=�۶����,�1��-"�u�-.��r�Ӎ5Ⱥ��p��?j.��=n��8�9�^J�f�#쒥XX2���v�T'j�+^���ݳB ��hZh�_�R���ة��3�o�_U �����8����8<��VkB�q$��Og�-�OG��N�ȣ+[��B���l_e�{�<���B��`�b]�;>����osk?�9��.1 ��1��戳����Z�sa�B&l�(�+W��D �sba7&GP��*j�B�DG���O,��K�AQD�շ��A&��w3檜�Cuʇ}�{իϓomu�-p��<�j�{�:�Q�p���"<r(����m���_C�O�m_.�]"u��8֊�p4ɑOy��h�	���1�#��(�'���>TnX��u�s/�{�uv��mHa�C:)�=4o�g[�MƟR,���U3�֦t�?ݛM&"���q�`��Z:�4���u$op�`D\��h!�D�M��o�>!]W�h�h8���+�I���g�5�ǩ�[�����rPH�O��dX��� cynx,�\����ĝ�v�Q�^UE���^L��I��_��a��AA�)��O�.�+ho��)<5]�=I�¿p�`�F�ut����{<¯�0��Fz���(-n��Ѕ�8垓3�������O�/�gf��s�7�Q�duxBC>_�hDW}^��R7�2�&����4
�6���ABNlj���>/.��[����%�^��C�������b�?�H�?�Ӿ�I��s��-W�"rŶ��H����[��i�F�wa�$�y)��E�-LD���r؞��ln�tg?�AȪ�67xP��md;H�wU)��J
b�o�s
��l�=G3E����L�v�u���k������JU�����4�l�����xDSX
�6Ʃ� �#���y{���@�Н4�[7�NО?���i�L�A��.4����, KZ:=�ޕ�|� m�(�_��#�q��Ow�]O�ܾ|]/����� �0yͩ�$-ڙB�k�N���N�����9&a-G���_�ЊtqLKD��Ok���?��\�+�bՃ�D��J����T�!
�y�j���du�)��eco��s�|rbɛk��?��c���	mE����Xs�CY����Af���+u>�m�5V!A���,S]e\��mb_�*D�c� H2b�q��xV}��: ����^��S9� A�\�A�j���+p�������D+N��whѤ`�J�#��R�N��	�]?������ڰigf���U_����(��#!(�5Fec�fKʫ�D^��`=<K�A?㯛�;��r����;��7����w<JW�P��%E�L�r�av�#�R�}c���B���X=�b)m��6�S�7	�Elۛ���򹄓^$�<�Pذ,q�Vw ���_��tC�<QQ��p�Fa�]�[�tه9��9��R�%�ũ)R�\,�)��Ld&@��_E:�yW dLjs�^)!��tA^@���O�	�(���"EXx�Y�4�x��j�>B7�Z��e��������}yY�5����
.�\��T���ل�}���튀u�Q�l��15���̭S��M����_MvhuIQ��4[��{½�߷�*6��,	����:6�<+-�gQ�H�EL� ��$7�*�a[��/��5�e�O1d�Z絋0~X��Ccy���ى�"��'A�Y\�f*����n�b����ј3����FJv��N����C��w]�8�f�)�<)j�`�&f>i����� _�U)��k+AQ�H|�be��HO+Y��j��d�A�я-�A�������`�;�W>Ĭm�},J�q��L��g����#��]L�6SK����O�v%�0�߸�]]9 ��y����1�"�)L2��4SIw�e��q��BW$�*�u����?�B8{��0"�z�Q�h�>�Ɖ�&/�L!W���56�'I��}	�F\l¶��<X�e��|I�T���HƆU�oކ_6�:G�ƺ1
)� wx %����e]a#����S�䈠�
Z��gcUM °C��6���Ѭ��y�~��h՗��v�[�q/���Ƽ�^j]�7L[�H���h �&�r�&�ӛё
��Blv�=Rk�_�i��B��*֏�a������"�E�a_�E{f�z/J`_xj��yy�6}�5�G�:/�. ־6��;l�v�!Vg�9N���3X�c'`9��\����Z���|�������������;���C���Y�i����E�(ۤ���uyѕE���t4fY^C�>`n
~���������A룄�\�TC����X^�4����D���WK
0̑x�z��:&�>N�?�IQ_v��m�����&�N5���X���vIO/\(u�kB�g[�b�o/��s���>�+M�<��-�)Qj��d@�����`g�{*�M��F;.���&�yVh	�3P"hq]mxQSĀ��YT_�h�����7fDD��u�i�ۆ�ry|�d��rg,hP��ݕr皩H����ùl�FbD�A��B�yG�V��V�X�N�Ȕ���I���;A:>E��LJ�ֳ�X���%	,��tKg+k1�Y�&������X�z�z�J��Ucy�N깭~}�b����0$IU�+���5ҙ����J���yJ��}	#�̹/�$ypvY��j懳Ϝ@+������AS����k��/7G�y3�����kg�Ɍ��^��3��'�h:}��X�`�1��)���+�XTuD5���g0���T���a=Kk( ݾ����.U5H[5��Mv�B[.�c���#"^�]p�F�*�('	c�ޮ�Z��]��ܢ�B���@�y�\���۴�a�dXc��o�rX�տ셠a.2U��P�߳$	�1��I��0t�C���\��=/�H�J����Nؾ����oKee�b�E�(9�T1MjITC�9X/�US�@��[��y_��?�2�%/�q���7�_�� �4��~�ݑ
B�w��A���[�2�Φ����L�FT~J���B�K�5$2�1ד���/5�T8Ӡ|�����!�C�?���߬p��4����\�nq�ȃ�����F3=K�����%�Y7��=H����ߍ`z���T��8�*!�F����'{r��T�Pk���r��n�p�=C����o�M5�$�T$�9k�āӣ�}k��Y��S�Cv��o�F�
�9�7~���h�I���L�'�>�����Պꔃ<e �
��>��t����I�vz��[jII�-m��I
^�R+5`c�+e���[J��<�`!����/7O��J*��,1p~����
����"�RD���N���}��	;g��	�������u��L�n��?t�c^}�T¥^]�=��<����sgz��m�u1M|�� ����m�ķ�*9��`��F�1{�T�W��39Ʒ}#T_5�Ŀ;��?L�4_��Au/��<��[4ck��C��W�V����Z���^�%�i;d����:�Wm�9��i+���{�W�l���tf��2�H�[�p��s�$��/!p��q��)l��N�eh�ӡ����g
@5��\	�N���?�n&���B��B�AfO���J��÷غwT�j>.\�������6eT��Z�=�I�1� 	�/�z)�+>����,�SSbMv98�����E2вE���0���8����J�$8�ߌ|OW��]�1f��Y^���0�f@�6. 8��.��(g\��zĨ@ �����/H0�LOk�n��dy$C�.%�'Y[��$�;�^o�,��ЎH�)�3�@��_߱�F�D���h��UznQ?���=�0mdK������>
#w��#H�p{Z����?����� ɬP��*ן��E�!~풯e
�o�Y��>Ic}�M�(y�j8�ֽR�#��A��-���)#�-�㧏p�{Q���E�w�cc��(���r�'3�d�Q$DC�j��{��@����T��+� �����V�V(2lY�[�e�긷	��]��zW�-�"�6���g���(^�ɷ�����K�-���Ck���9ښd3\ #��L����ڡk�,�n(b��3JGv5(�X�O���胁#R��DnR��hgL��|RQ�D�s9������է�9=��-���RB*���,��$��=�jFLKº�nF�Đ�q�ne��~`mU��E��/����{?X\"��3S7��FߏH����9ǩiV�5`G�u�xv�z+A��yE�Md%=
�D/{޲�748�e�9�4��PG�ܾY�hr����@	Ek�'��q�P�߄d��2�v�`ź�%�:7*l���w�{�q��buw�A�f̆fNNy��I��"�U	>�h�·	��Jlnˢ*H4�s|lf)jZȽO��x�K_��f���G�hLa�e��]����M[?I����G��fd�iò��ۈf槦B�m	�[�p�= �'별��?{��շ{�Y�ci���>37�ΒM���\��$��Yqݼ_�x6;tuµFU�#�!�%������x�w'��W��O���~o�z�S-m��W'��� �%2t�Ќq�+5W�&�������v���L��{Pp�>��\+�j�Wil>َsa ����ґ�.���O�����wIC���Zp��ځ;����$���b��r߇��v�'�T[����o� �!|]��aEe�Ǹ렔W"�j�ą4v��5���˒.8��݃�-
��7q=hy@��M�x�iP+G[gO���Ƃ���Nf{���V�aO�I�J�v�Pr0��8V8w�u��^��@�i
�S�V��X�E�]j�[�����u��jc��4*<'df�qG�wCNcء�$AXG�#��������~||\��ٛ�.�f�e�m|Ew.K�B,�|{��6]+��U�?�ro4�o5�F5��U�����F�%{�ÈP���wLAǘҎ4z�ķ�ۮE%]��x�R0%?)l\��с�ш���y��_hg�"�*G��>���b=[#��Q��!oC
d���l�9v�1�y<_`b�#6��ȑ/ 8X�l2��w�Ƌ�I*��v�S"���C�1�X�<`��SwǨ��r>y���2w�uTc�}�̮�?��_F�4M����F_���Nݫ�I��2yVO ��@����t�z�r.!T�<�|��޾�r�9�W31�m"�1�Ki1��;W�l2�[�rPh�RԊ������PN�ڪK���.�F/V�<LIʞ򺄐�<�������VOB�n���8bA��/-���=�Pp��+R��.v�Us�등ڳ8!:��CN;�o:(��tI�����B��Qc�w�0iP�gW���QJ&�sak��X�ȑ��sD�~�
S�AB1�g��^���b>x���q������f��d�n?���lۛ�v8Q�*?rf�j5f�z��Z>� >���/Ci�g����'��
5���S��5���?��x��d���w�B$O��W�m>�CԔۚ'*W�d�03U�|+�83���i�G��\���
�B��{��쥔���#Ӆ����-�caxK�c���i /�Vv�.�M��Zz����>6,�<Bx߃�-�ߏ ~Jlm,����	9T�f�G0����'(@�u��/@Y�L���/p�[5��ݷe��e��+4��/��)� >V��V���0"�K���'{+w�VR�����5�XQe���x�1�����:D��]��=0�� x����/D]���,��89|MXS$H�CL�e'�������]2�'/�G�����=jm.��X[h\"�yuĮ���J�h��Uq�A�q_��>�����xM�R��0��`'TU���������-���Fo��4�R���DG$�c�h ����� 0�����{-c�U�sN�iQn���"|><�"R�:�^��U�3��ir�2��
(&�+|};���ܨ*U�Vpy ��!d��jk�zEp�)#Vzϲܦ@|�����Y>`�?\:�f�% ������yQ��d}�8��n$I�WdTw�S���ONش�"_%�b� �x�m'�$�X����y�(//Q[��}��[qod���Mqqx]�x��Gq5'D���<�'���T������:*o��#T=VL����u0�h�oz4��3�;�YYu���A������]����z�GuOgy&��:Er��5>�Ο���>�
����)�$���R̈�$ۗ�"���53��:E�<��ߓ�	ԯ�v^�E��|@���Oq���>��ˬ�����#t��ui[
m��Pa0=<��<��5��`y�,��9���茆'�v@�.�*}d�k`}	��J���!�b��F��� %F��y:��߭<�2��z�B��j�|5�B}ɮ!�A��N�o�Ȳ���le��D�NĄ�Ñi(U	�%��ٺ�o]�����>Q�)�es���r��a�*�$p�k�i��H�I;F�����R���G�b<��N���P��ݪ��+~V�-;��%��ּ��H])�6~UZ0s����U�7�_F�� cf�����G�mW�eA>(8�@E��8"HqÔ�ܳ���d���{DWY�R����B�������н�#�g�L�A7^��H߻Щ�@ت����yX8�4�K�9�3�ĵ$&2�_N	+6íR�rP�jK��;c'��j� 5��RvVZ$���?N�!l�?����G�=�!_��*�d;��D�6��R5��<9�?�dK���s=��R�ԒT��h��e�'0]�?��+���zq���)�G�%b�K���Lj�F�K�g�?o[�yX	Wπ�nL���,��H�H4v�'��y����0�㻺�$��|j
������.�͋������Il--��k&PSQ+��Qbl96E���J<��v,���
ó T�h��jd��D�\�^do�#٤7�~/s�%�"�1����"P�V̈y&�ʿY]Aܫw:C�$�S�������غ��8���y�>�-�'�̎}����#�IZ�K�th�n��3sf�G�$�r�xbl[���v��"��I��,�ٻ�Y=Ey<�H��̼% ��Ӫ��������|�@���K����Y�>���ێ���'�� ΏF�F��~X�C�!K�ߣL�!,�_���J&��F�'w��!�!L����@�~���qg�$#P���)6L�sN�+��g�cߎ�9CtZ%��b�ǒ��a3�>�,�u�W0���@��%4����&��˅z��~8v��jt�[�a�.,�f��Y�3�\0�],r��4�~�B8�t�1+�W��;Ӂ1�� �sn����EW5����@67�K���'���MZ
��K�d;�ٵP���IlxҼR���V����H�Y��xt��3�
b�@xuL�`��gv�ɛ_�cj��R�Q�C�D�T%q�R�]�E���BuB�!.��D�2=jߚ�5���B� 	\���<���#������"�U8���T���E�Q�)��i��3�~Kf����5���f��_f\�*5fzͥ�t�j�e�#��zf|,)�v�qK�}�d'�L�c|�؊��4\�+��k
1��e��2�c��P�dF��h��B������ۭ��?B�Lrٴ}<�L4�Y������,0���t�T�&���y5��Y�4X�#�H��|Hh�����9��]������M�����ܛ����u��޾����{���M�gn��������Ws��'K�y���	���I4���J�>h�<\c�A�=I ��
�^ʍ}:������'"�$əZ�,������Jc�R9�_���^9���f�`�d�+K'Za�7���b�{��23��;P2�_	���rH�d`ʘA��e�xUm�v!��`;vw�����I�����b���$x\ҧ��O�J杫��ش���Ñ�Ƶ8v3��ah�|�.XU'��T�8/�%��d�����tF	V����#`B����x?�
c����)<��|Rz:�ı^� \F?N��lK�ď�:S&������D7�ı�����tx������uLx��[Y�}U�ky�7�����SP+~�7,��1�Xm���2��M�5��V������7�IM�|�V���>��b6̙v7%���@uFp��1�����E"mL���qޚ��^R%8��bɤj%v*_GG�d��&"߹-e��t�O8�lV[p0����zҴ���vt��������^��^��HF��[^���B׆���/W�V������m3�n�=4��rG<�)��鎴|8)�EjQ���1��_�{���{"�<�lG�����d�ۛN�M���ekeh4�ƙ�v;q=k�TFg2�8��CG�%�<V�����6�Gj��xkj؁B�v�x9{����K���w�* ��@ͅK� P
\�`}���tߴU�����3B��T�}�j� +�0�|0��o��� &�jp����������~4�S�s�o��'�(sMxt�h�*�
�M�GA	�+�i��3t�^�w��O߯�~bWo��}��f�l��\�'4���ǆ�+8+�I�1	�sv�#Ģ� ��ͮ�I�f(Z��ݚďo`Q�c=���z�0M������!�����'1�`���	�GR�pe��.1`gg	��Q�Q����ʨ��"S�9J=Ѐgk���!�Kkf�X�A�Q�@6(�N�NP�n�ln��+�&����U\�֍��g�1�4v�9��/�-��4@]gC#�����{s�_�C�"�F�ҏ6��O���䔻�>�sj	W#d�d�60���0�Z�q�W����~�:������A���f��U(&��;��C3U�LCռ6�Xv�����R�6��ف6,��Ŏ�s��bBO�s� �E9�����!�]í �z�- �xw�yy����f���h�T`�b0�����*���c���y�
�8���;�n(��������z}w�1�N7Ϳ%�,E�p�!�u��E�����s �|=!�.�6ȼ<]�qQvEr��,	M��S�`�>UدbH�h.��:ȶ��ӦȌ4F.�&6�"�`�ʕ	�������gZ9khk,ܡ"�K �Dڪ�<5}Вs�ٟ�07*�u�Q.o��/n�r{È剶	oSHM�W%!�k ���TG�?\�'i�B]𧃽f�Eq�ZdULW�J�V<�wF�v�U�U����W��׊�Q�J�]�la%͛D�!��Xs y=Q��-.���JT����ٝ3������s�]�����5̄��z!2�z��5��j*{6 ���?a�d{1�c.�f�@Ե�'Za�o�lGݚCK�`gJ�� ��k�Ubl{�=�S�{]�YZl^ȴ>�Ȑ�����HH�'���
TR*��~9�������9��"C��w*6-g�i��8j��[��H���ˋq����M��)!�3��6S�L�&�k�OuN$8��K���=�� ]�^]s(��Z7�W0D��((�|�MsK�u��I��˚�\�_"�F
E2��O�$�4=�f;}����j �S�3���,��mU�Q�|�)���w������S�!md�����H��<}
����2��B�{S��>���K�n�đ(����IH�>�uF��¦��(w��A�;�]�X�Q}[r�uO�bg�����)��QWs1k�1���~	��>�$��
���k�09�����U��fu���y߮�Ya�|�`��C��&�����4�c��Bv4.�L�	逫�Lh�	!��u�C����<P�8�<OڍEn�"��^�RW��xs\�ǰ$�d_��*<��݆`"�"}6%=��u72��4��z�ˀ�@�ԪEp�[M����2%�*q�������c��g��TXL[ى��j%��x	��f/�2"H�n��F_�c�j9�׃�n����}W��<7�5���co��NoI|��t4�Ù�q�܋Y@N�>�M��aV�G4�N��4 ����*^���^-�΃.�mq{?c���eQ�Dh������a_���ߚ{*��Q��:0�쑤��0�NH����I��k�X|�/���w�$���K��Z�b���N����1��9�L*s�_:�Ɓݜ���xi�Ğ��qF�*|kF���w5c5���(S?;�5���7��As��v�U\۩]�RP�U���&����ԋ���Q2/�D���7�,90G�<Æ݌�V�
~�B���>�I��6O��D^k3/9F�1�'�d���L
U�>[�'���_�q.~ģ=D��o$(�GܐW-��m��t;��ធ��mF!VqT[-�-��� |*��p����`�Q=�i|�F�!⁋�{=�G�a������U���H��X��t�S!��Ĕ�8��߯ة���|T�:���k���7�)�qn��Q��*�O�����j����ehT,��Z܈%RIǌ?`��g��_�Gޯ��PO������ll���Ӭ|d�����?��Ǡ���z26�c�E�)h���܏^�0U��x��+�U˔I��.���Β�n�\O.O�8���� e�^&}�D8��;g4���`����Lo|4�,�"����,\�FA?ުd|"�2O�aI�ē�9��w��f���AV��0_�Qm��� d�k慒"�̸���զC'�;���	���̧h�;~{J���O}2�A߆}~ߚ&��$�P��(����C#1I�b%��jtzyHQ4�
�Ԁp��d�@#�
� ����@�v�šV������)��l�a�u��t��*U�3Ų�z�Q�x�o��l�/��}�ю�/q?�i8��ޖ������d/a��ђ�b�*�<xw��9�[�u�Tb�%�XK�.p��O,�]\����ۘ\�·c�R�~A��l�UZz���_�2�w4>k��*�cso}�"�a���3A�h�LTA���P�Q�����#���� �v�)��.�[��c��/�CF���ʋ�X�-��XT��E��c��V��~��\2{��˴��.
�\"���1�%��	�<+�8D0؇����;#��)���~�M���qPq�[�r�ۋ�/l�XgW�7+�e�U���06y�󑦅,���at�!vڤ�z�MM��0A���O���D�g��P� �����������1��88��m���ě�:o]�8�R��RH�u�贕� p-B�72�-ULy��B ���w�PF���(y�09�����	Զ�3�v�N��Gr}>h�Ǖ[��f�.�_����HJ~g3�w)�	,�;�|�fx��ť�V��W�x4Y�t�L`Vl�%D�w�����+Z�5���kUJ�e��j.�;Y��w��$b��aG��t}���ix(V��?r�=ov�VYaT������jm�$2��K���W�B��3)��k�9l�Z4~�yw�R���}�	P�д�%J�e���7M�BUJ���8�yBw���E�l�'�7�$�� ހ�%>}�]�иvnv~�����1�TV���5���H;�N�?=���l��wn��1[���91+p��l�\
U���ˢ��Ҥ.:Ş�ݸ6�4FEwj�1�m1�B4>�1�DTrފ�R�U�jD�f��(h����c��I��������S�V�*+m���I4O�L���)a���'W.�\�U��cӆ�rq��e:��� /C���IWk�-:Q&�"�"��ջ���;�*�Q��{�8�r⍨d��k�ň�$LY�LQ�lB�0�h�I�A���9+w�(q�a�d�9]|5y���Q��!z�`#������u�\L�4�A$��h����\�i�x�qu�q�Ρ'#d�H��p�p���#9���>[�]\'�ު2��p�_�s��;C��C�߃��j���!�tf�g40�V �3JT\ Z�`g��`�|H���
pS��]@-�H����h4���u���Bﴑ�"�{���B�+�3�:zT�������w_N�Haa,�_Մ4wF�aƚ�F�����M�;��y�#D%Fz�����[M1Q �)ڐ��^P:���	:d���x�㥆B1p�9S#���b���kb�l}��I�M㱵r�!ri�+�t���;���eb}/�Wu� ��p*p�� ⥏r��ӓ������s�j��1�M���S�p�=R���wk�S���<���ëk���W��&��!�2D{U
���[�^1�2�$G!K4À��Tx!�l�c6��\���{��pGA.��2^�Y���}�v��G�`�R�ۅ�[��ߝx��?���a&֕`�ģ@��x�U�����:���'t?zs7&���E�{�)�4z�s�����B�����p���ҫn����>ۃ�D����e�!C$�ݶ�>��K~����Ʌc�d`�,��)f��H��G��}�w:���w,�s��"Z�~ՐǛHr�0G���BY�ܪ�����	Q�M�L&��P��g���Nb�UT,���#�¬���ؙa��2<��1�N���3:|�������<��q�s��zC����ۣ&?,��p���Q�M܌�?��X\�N�f�Y��<��hQd�<�$ �j�Mo������Z�vB�J�5^�ѐ7�R����B���ы��V�u�̈,�8�@ìmP�۸t��V���j�r�>���!�-�X���k��gs����H��^q�[�~��u���!��C�Q��B(��%%���
V}��M��&�JD�I�y�ގ��໠�C��KNDK���판�P�̫۽�?�ԛ�aH�I�5Sa�h^�j}�)�3�-�lG��kJ���n7w�Kͱ^��;1����v+�ߡ2������֡�¸�gY	���v�\���g�0@�+5!����T��T�+�^Qkv q��ǿg��@�r�:PE�@���̜�n;��x6\&����9L�meN��%m�8�dN��vs��!��q@il��ŪL�S~����r�r��G�k��	i�0y�,���3��e=G2��aO̫���W�&o[�D�>RE(ӿ�OD6�yN�&Y�����<��8�]��H�B؂�	�����N���~��p�(���1�`�TSv"}�'Ƴhb�����J�]ﲐ>�xaӭ/�re���-pQ��3��xcѝ�]�녞'��+? �3b�Tw�Y8(5�+���9�� .��F�k�H�&`���ڲz��(��V�1�4�g����w&�}�ߣ��Y~@(��|�F�+�ϲY]�B�j�*�����U��6��
<g�.r�Y}�c��eOY�H�mBX���Y�`_�c�J�-s�0����e�UGV�g�i)�fms� ��,pk��a�H;wgS�'Ȏl��e���z�w�L4��G��+�G���h�*�/�m�>K�^Dw�1|;�#���u.��"9tG&�!���|YT��#��.��N���X##���أ;E�)ˇ�P�j��s��ZZ�~�)rsg,�o��c�K*dw��X-��d����,���A���3FM{}�i�ؔt���̊��h5�,Z't�!�lh9�OQ�!fL��rMk����yJ+m7�7���/,���Ps����
C�;��a�;|9�^,Ɨ7w'����c�,�m�$�k�AZ!D>,~c6�]>�}������xan��$m>���E��<�ը�֫�b
�y2Z������v���:
Τ�$��� ����8f�,q��E(P�c= -�_��2�D8�]�	9��n�l�U�w��i8�Hx#���ϙ����ۂ6��T� �>C2�G��I%��x�樮n��v��.���g"hm~��*RM~w��/���Z�A�Q�	��Um�����cB�'��-
�g���|�*�{.���@�$����ռ
ʧI>n�X�񒥳2)�`�����(�A��.y�3�-<<�bVC��O��3�Xy���:@���RIh-��ٲ$)Ձ�!���B��_���|���Ա��/|��ӭg�bz���p��kM��)��5|רZ��f��<�J��u�V��n�?
�7�_�l�N��gˉ�2��F]�	���V�k2ˇb���Eټ>NF� �R�_X'pw$]����.��9� ?�Hi����XWp��2M�b}C�',�&��ƭ��.Am�O�3Wv�Ry_���}m��,r�h;_�hݏW����wM�tt�~�~�U2�)����5�%�K?� �?��ˤ��fu�o�y�sީ��ƣ��j�L0���67Y);����G·y�!r �2�?3���h۔sL�'��(�٦4Ҡ�cg�ש��dwû��7W�e*��U��nۭNgJU���j#��H��P�k�Qa��Ȫ����>-��\�:�>(�C�X�h-B!0wξ4i���;���J�]Lg�w�hS��7}�0�?`����ӽ��_��F-d�qR�<�vWK��|��TA�K�h�G�e���vٜ�Q��m�7N�����7HU$���Z������iZ��A�.�_m$y�2'6�~�,qT)�B���IF#G��8~��3�y�oU�6��b}v�Ս>���9N�����Ȫ����\�Q�I%L �!_�kks`�B~{9Չ�p��!��S���y��v]ǎ�#sJ� �×3��G�<��[���bj/�$�̘�y�������{=[���S�#~���ï�����A���$ρ�]���i"C�1��g���6c�����;>I_$9P�$$]�w�m�;�툲_�f�I{�݊"Q�煮���5�BF�9�+���̢�w;=@��h�3��;�Ľ�κ-Iv@�m]�Q�:�ؾ�!�:����CW�$<ϛ{�\��d|g�o�ζ9}����v�Z\[�(�w{�9�#:4#s��W�7vO��eX���"���a?�ۃX��F_k�L�Xm>;�װv-��;Z
"�Au��QX�o+�L����,C�g�m��G�Qx$p��m����2�~�.ɍ=�dD�U1d� bSW[DڸS�Z%��X��H~@��ә�W,p�*��jB.,��E�e�|N��Xr�����ջ��u��H�97	��WN`��$:�=��m�u(�#���k]#g�����<lۘ��`�D
���y��%��5�fg	f6����܆J����_�v�X�=2�}ӫ����^gӧ��,��2�B�S� ˮ�w���+��8y��'�kd�#��Vp	әmC$
������TE�V��	%<��S�N���>:��5����,'��4��&��D�l^q���{��n�z���+�}�[~�>mkA�
̗�_�.6�E���.Q2�D��^��F�	���B��YL� /����U�ϪPR��2}+9��8bsK�-���J�+K�u�r�(���-*�ƚ�K��Z�;e<��B�@�c�ۿ�@	ȇX���V������L����)��Ճ�ț��B�4���ul,xr:�H`���qҊ9�ڑ�p���&�ꇰ6����+�8�=?�9�-��t'es1�a�9�2�㿼dZ�pk��֗�?4L����-��e��7�֘�+,�����r7%/|>&R����Y%��5\Ҕx@�:Q=,�� �������bD�i�t D�7��wb%!Va���,�o��������m���ԺvO���8���V��	��3d���$��]��!��F��������0��)��-J��W��/��6�P��W�e�D���Kx��J�4�ŷ���މ������4R���T�"�g�TW>Gs��^�6UDd1���{��d9U�\l>�m�b�Jee�R����\G�|���d�D!Hj|��O8�N��Y;��� �a���!`�`Fi��֮�ޑ`Ҹk�7s-�(�ey����k��M�c�];�κ_�RB��&�΀�:����D���{{v��b��[�=\�9ҭ��ۀ��w\ȣ2�(>�V��,��9����$��'u��a�k�	����C�1Q�
a�|xܿ����W���+��;�uE4!o��^x&q=�)�ģܕ���X���B��1�j�
H��9��v:�$���V��Hʩ�t�G44娉�c���zpC�z���-,Jg� 	�P�o�R�TY���*�&`I�R�p�L����0�YF� �'�~�����_���W&s$"��=!q���8�ED� ��z��G�G[�ڜ3�&1��l�l�l����rŖyI�q}�zﮋ)遙
MU	6OJn���I?N�c��5��@�$�?��z���=al���R��lU�jB�T��p��_�0�|��FlƱ����ޑb��@����'1���������}���:0��%9�r�0��=��:�.O���E�ˉ풼V����ݟAe^m=�zr-�\�	:��b5�uѐ/4N�����a��[?1���=I� 0ǳL���QݽŃ�����MW���D����,�0L� ���\�-�����L�,�/{��%��#�B�KZ"�����_FW�%�I��)���48IP1�����tG��s���ʻ��i���X�n+�"�"�e#�b�:��Yd\Ⱦ�~��{��7jD�H�E�*��o�� ������{!�6\�bv��f�d���'�s��}5Lk����vh��w߽�A�o���O�I��<�|��a�}ӎ�@���V�\f�q~�Q��z�T���Id3qf�r�yS!��c)%�Cm�8ˍ�bqt g���[��a�������f�k�h��m�HH�[M\�r�k��@w������֡�BP�Mci�x'X���`��̸`&�ƌ�"�C4Ff]�Yօ��'b? ��V4oNż�:o %���V�1�	ϔ��+�����P`�.7;d웍�
��j�N����{���ΒZ�I�<�M8Yw��,|V��yUJ.���,�#�1�^�Yơ��sS��S�O����o:�4���F��Da�o�����-��r3�.�'�F	T�N�A��S���B�'���@�*(�z�,�N���;Ѣo"
��.=���s��`��8���OL�X�P2
�w�	3��S �H֏����f�E���B>��^E0�]:�d#n�Q���w^��"v��p�ɒ{�03_�kx1Fv�C�e��2V�
mم*�%f��K�حn��5�.��>̳��x������Y����y�����A���
���������b��[�ó�w-��T�q�aS���%ߕT
���!�	%�� ������-3j�������[	��v8Ā�@�������r�g��ᮎ+?�����fcKw[+8��mZz��\V6��ߐ�k+NBE@)ER�d�����iS��N��rW��+����'��v&�C0�|�����LC'5�ϑ��)��)�
:�<rJz�	���jކ�S�|EL��n��C�mb!md�;(��:�o�����[.��vǇ���۟�CfT:��樄�(�����xX
���Xۣl���7Ԑs� �,m�b�z���7���R���8����t�]T��a>�MX�3k��W�\xM�r�Us���k�MH�"]Y�_ݕ(b��������䪤I�Q�/��{��&��}[2H�0`i�I���Z��W$�?d���CQ#�	oGl���3��S�Jۦ=�Q�G�#GB�C����%���]�M���#��vUw��8:�����v��~}�Ʉ��֞����Q'iO]�v����u �d˥8�A4B�!M�tx�_yz�o�Dt.yY��3�Q�w���j�̂*��:��M3�UѮ#�U� ������"^�~�ma�혯���-]�;���.��k�5-��l���$>���"U����k�*���&�吴q���g��Mg�/�uܭw�*�o�Wdα�~�߶���uSK`����X��$�^V���V�=�f��^-�z���uZI6��W߈ME��o	�M���� x�0;J*'�h+���vuad��#S� 1��u�Մ�ך�I����ѓ��^���Y4b���H�*^����tP�Lܣ:Ӗ�JJ�5��GQ����Ua"�����y/�� ��V{W4��˔[�M�??�_~_��:^��/�q��v�k48�
A,��s�����Y���q����-U�(	����o���dcG̭�8
�#��`BaA��8�VO�x+2�~Qk3��,�f*LF���Ѣ�-!�e��B�p�^��A�^#�uq�o�GQIE9���]r��Cd �p����R �����i/에�z@`��m"<�轘 �P4G��\��L�B V�!X��*��UK�\�/��=�~�Y[K�2����
�<^�6BJ/��m����E�b<Ӆ�n�/�J�I�i���X2\S_�T�.#u����n�/����q?���c =���2	�����Q�Yř���[t�:�nB��;Y����*Ol��>#�Ɨ���������T��ȶ'��}`�1� ��ICv` �-�Q���c�������4S/���?еBI�P^��!����.4��<��PB���KEL�/�y]7�PA-�nKV L�~��Ƚ?:����h�^���Wu�	O�`[��AF�ݗ[��H�B7�I�N���DƜ��ZlK���y��2���<�gb��2`G6�y"vS�`6Q���'�cJ2!�c������^�p�N�0ak��f����
b���B~���]��F�ڥoArq��<¬��^"���yX�t>���_bj��5R�������ʺ�c�$_�8
C�O8k���8��!ds�a�?s&W���%��N�M6�оo��K33�U���9u@Zq����w#���(4Q���֌���q�$Y����5n�q���~}�Z�C�2����V5�/����h�8�J{��a��l2vP��>�Ww3zY[ �Xъ���f!���P�xgٛy% �(i�"����|4!�[j�(~}�m�~N�ܮ�ُ���o��!��@i.���	�)`���b��-���4��N��M�m�m=����h�l�F%�m�F[^���R�����FQ��O�w�T)�چܤ�0��h����܂:ϱV�K9��]���Ч�z6�=���ǥE��{2#�vk)��-s�lś5�wO�E�q���K]��Q�b-4!��h)��2�7��lu�@4��Ӡ*����iY=+�R}/Ο�|X��L��Oey�_C��yY�Yq���h��V�\�'�'���=�h���#�/�6qf[�*@�!�s�
�aV� %�[.̩���K���D��Pg@c'��"��=�-��O��w�:Bu�*
�����͘����j)��	?]|�kSD��tz�А�%���栰�J	�52^���������Y�ݎ���	㺺St<�eㆦ�d�m�#s�D�KxX��z6�2�j������1�[3�믘,����V�B����U�1o�0,Y�0��~.�>��D|k^��݁��۾㪎�o6��C���С��`���;���DM6��K��5y�j�Q�#(�ދn%%P�q�ǰ�T]5�C:~�¸�[C��'kAQf�Z�T63�y踡�沑����\��Fk7���Y���cGaF"�7r�-�6[X	k.�nF@�jO�R����f=6�P⎡�"< 9~lC�M�h?0�Q�G���|�F���(�2� �\�;>r�8t�pV�\��Y���x�7���u.�,��ֹ��AY����pV|Y��m*������u��,���+���I�������y�#��PpR�%ȡ{ 3u(�آ+�#d��K�q�q�}9�V���w���ފ�ƈ�L�ya65�|����ҁ+�ˌ������A��������6�5�Uk��/s���*!Y�}ɍ}�ʐ����@$�m���D)Y�}/1z�G�(�z�6�_0��
�W����������fk6 IK�3��0���D�{*}�S�쪞��#`�+5�n���&���?�]\�������t#�G%=lK6M���}ҋ��,��*����يg��]�-ȭ�#c����,q�3�Pu?mr����)P�CQ�0��6E	��!@7 sV�IC�;�q^�+Sa�����s����b�"Rp�;)�bÒiz�-�d;�!r� l,� �vA��������u�.-=]=��o�Ί
�#�g/}���H�����lh���cyݒ&���C)�c#p�j~i�0���ӹH�	%f|!j��M��Om�^�i=ق6w+gp/m6�P�X��W��0����f�G����4��˝y�tl������2�)b���޲�O�i�Ѓ/�ĺ�e�^<���)\�`{it�M����(h6uX� pb�i�x��D&�~9��]��`�'DJ��iN<��Zh��r������T�PP$�
�멐���P���]��w�
��I�¶)�ˠ���H:t�w��UIj��� �G��E�'3�D�߆����)	̮~0�#r���r�Z�� �=��ԣafߤ�Q&�k���/��Y�P�*�>���dQ°0d�ԭ!wC��QS�#�ҧS��<��fAu�7��<� gf{���>�Q���|n<*/�~"��r{��)B�� S�Q�7K�	e�x:��i� �}R3b�u�q-�}A�:�����^�O#�h/��|��[@�Co�4y�b'`l{�� ��m^�f�+��|#����-Y�ʨ���G:r��ӄ�_vM���`_�:�N��I�IZ��d����;���b��`e��~�^:��LH]�*��ݽ�#�n)�(�������wM{�!���c��Xu���L��;�(�%�t�ZUy'�&꧚��%�P�T֡�BB"+�2r2gKoN�vF�dQ(��9��!���v?($���+&#�M�+}�ՙn�
�o��]$�ӳ�>�G��U^ui���iz��b7im,�������V���`���9�h=~���:��đ$e�v��g������a���L'ed�
A<cZ�"8�KZm̮;������#��w�o�'���6q��`���dBy�6���9��~y=+�ߚn���R��Z���ΡM��<����3i1��::)�	������#�1���@ޣ�����i�ӆm-^��	�Q�|@��S��������--��(�d���S�W%�8ֳ,��G���܄g8��1j,��ki޵X�1�{[_2i�0`��(ca,tB bO��2�#���*�x;U,�x�⨈h|q��:b��|�Z;�2��T�H1�ûRF��Rះ�t�=��,�9��#5ɭ+G��kݼ��乷����A�-�l�L���n�	�H��1hW��HY��o�����~)�� ����[s=[��-���$d��������ߧ3��Fޏ���u�~�S-�7R��6����
��&�]�zT��[$�Cw��S��Q\H\\|���������ʉr�v����+�y�io!��٨�j�4�`����oc{���e1�����g���O�)��6�����oW�$i��꾣 ��ӫ[m|n��&�z&ן����\{�^:�y������-l�է��3ۦK�G�Q)�Y	<��o�!�r�e��;h��$@�w����&j�w��UyH������ �ʾJp[q���6�� P
�����vR�:"�?�8��|�B��.�+}�C�1��;k8a:ůq�
�`�x]������uz�s^�����!e��l�1�j�+2Y����Y�D.Q�jŹ0��KO�':�W~��q��5�俪�ɪ{n���.�1^���!:��Q�e�+�f�?U�9���>k?YXV  �7ai>�E��v�����M���rU)���瓼��%L�E���RP�����;��� 	h'X�z�CO������w�&�h�z��i�54���Z�ܳ�t��.^>�G�/�s�I$�I�Q��܊3�2���[���e1���O]D;b�ݿ7v�@͈{���2�nq躨$ Gm
Dtv�.Z4Hrbq��)�j�O��;.�.��v���.�Lۦ/Gs!��I)����};  �La]�sA�Ԩ eq����f	������MI_;IB�c0�F@u�_)�~� �*�0{�e�Z��l6M�1<F2�v��Μ�&���ܑŠ�ԽO�Ӟ;�Q�W8g���>5�����4���_AO
]����%`��?T��/��Ko�� �$H},���Q�0�'�F�o?s	�o�֙T��4�xj�GN�m|�G���dJ�@�����V&����M@c��ř�T����_2,1��e,y����#{�O��'3�\�9��)��]�% �װ$9��,nU���I��K��"�i�83.��xcJ	�9>�4����F<���2�i;7�v���!;� NP��\{����]���|4<�C��R�ćUG��,]s\��B�����|�PdA�g����y:��N �]�'����qQ�ߌ9�,/��K�B��.���U�\�z�f�ǑدƷ�oPq���mQ}�x�~�V���(q�&�Xe��o�6�&��,�QI�4�N �"���r,<V�s0~����{%0�q���Iz��oV �h���m�II�/�P[>���0Rp5���<[��#��EF\��1#8`��8�ج�[�2��!�tـ�dO�R��C
y�\!_�CA��E�褱�ba��t�Q��.k6q%ɫ%�uJ�b���Z��5`���'��g���7q]���J%��i����˖�4k��I?R��gS�W��'�P.y??��|ɧ�����_T�2|��ǤL��'�04�y����3A֓we��r�xu����F<��g�|y�9���6(�R�E��uNT�g]��X�W�w.C)OF��&���#�P�B]��%#��+��&�9���Uqk\��%�P7l��H7oU�O�O�|���e`=�;M��r�:�ϕy�$ n���}gy� zK�'rE�S���R,���ķ�9��'�	�]/E�&��d�l*X�˱դ&��A蹭�f����&L��ԯ��U���o�m���kq[�=��$�����Ed�q�ɦ9}���ģh�7ZJ,X$n6kQ-G�'!*���3�������8��*��MS� X���O�!*��|L(��2A<)���D���35�fr	��%�0*`�>�L�X�9^1��/����*�����<A6/u
x�3���*� =2�^Dn_��p~�!>A�68���L�w6w�c�}�L�Vz�F��6h� �́5�J��h1V^�� M�+�4� �=�W��\uM�� �7�R4z�;ez�$�x/�m7v��fX7��$��,�i+���{�l�?G�����E!;�ΩF̚��n]Ƙ,���Ǭf���@]���Zp�X.g����pIz�fp�$)���u�/�8"���E��p׵��-�R�cx[B6L�S��,�P���C,9�8�h[�A��3����F{��+̎0��1I�{@W�����OjE�K/u*OK�����ڥ|��8{oSAl��q��������l�����xgc�8m�'�����=<$�,�pK�j�J�ȕ�:+����l��y:S���?XJOk���p>���o����AQ�.������;��O_G-��K`�Q�.�DW�F�F�"!��V�w���!ş@y��fd��lLB]�e-<y��T�D���
P(����w���Z�T�e�"���^��8�m�0^w`�������?&Z6&_@�����)��������o-U��s�C�o]���x��w��LZ5��RE���SI˾�,"wPƩ�����3أ�)㘖�{g�#O�.�¯�׎O��hfP���~���.����)+׶D6��WCMfj/�����U�:t��>����ߑ��R,x�̽��a�lj�\�w�H�:;�;�%v�2�|��^���͸nދ9�~��_�Cu��yĥ��+y|��<�g�z�����2���
GF(b�Yn�x>���h o���9��G����ٿ4e�ͽ=��s/�0;Y:ܕ[Sn:s�հqiL:)aw o����ٗI5�F�t����Y� �;0�~]��pW{f<�5c�t��
wY��Zlg�/܏�
L���B)F����>�����#V�m�wn���<΅�uc�>^�)B�J�[���0���Y�c8�f*'So��{(s6�����h^EH�l�ƨ]��-�oАsW�Ŝ���#x��G7�~U?a�#���]j�0��{Z�F^��e�c�@��ҮM���V�����vƦƅ��c%�����wJ����iz�kB��1;Za[���y{�GY��������lB�`�,4�~��\B�gH�3���� :�����<��a�$�>�A� �΍��(����hS&& ׎�?����
�_�!SqhGi�$І�1r%8��n��r���^���UZ	n�ܨ�t��V"ʻ?�������;(pgw=hn�l+��ӢD�Wx��º�K�7
��#���7��9~B����Tڂ�e��ٺ;�'ڃ`S+��v{�;��3����<r�vN��{��7��U)E"�;�x��Դ�3�9$��L��1Ms�7̗?.�9,sa	K{6ѱS�L��q�ns2�M�u^����E���"�4ک�hnlﻩ Bw0kn\y�PZ�������v�tW�܁E�ڵ�=�X��~����l�V��~�"��;��y�3��FGxÅ�{�z�&�ʋ���\v8�����IO2�9S�]�ϴpn)��_.4b��ؼ}a��U`��1h��p��0��p}�U�]QGѳ�I>;���]fF����5�pM��z1;��;�Ճ�D�y�/�a�,��5cZ��d���n}����5�"=7�<y���l�L�Ԓ4��j-�_���{k�H�5���r;���7�j�iK:B%�0��!]�5@!�Yn)���t�Jg��l�^<M}�	ĵ�O�� �z���H��>�i)WW�БX�y�����Y��mV y��n�˃���5�i��F��᧡�f�k�7�m�n�0�M���C�3X� �D�[x��R*}T{��t-����Q������K�M[��1�~�6�i�9�@�{ip���Y�o�����9A&���8D�qF:e�G6@���j�S���0P��<��5G����a����t��X��x1���������`�81��Llm���N����V(�+�I��	���;��F��Sc�`0l���E�j�0is��Y���
�1eg.�f�����VιP��)��J�q�'r�o���Z�~Ec��f@l�2 ���3��c,��g������c�1��^�'"����7�TUW�7p|�v�Y�b�]e\F�>��A�Sw��Hk��e�:�Fl*v�^�{/���j5Fۉ6r�2�/�W]H4��	C!e�A�l��SP[�-N�F��Q̵����#¯�_t�X{�XhE�v�����V7���Fd߀�e�hlC�X���W��d���8,E�{|��`�\5�����(`\��3�7���e���զ��C�a����7m�$�V�	z%�MblT�t��㚔�hD{f���+�
r�.p+��m���[��C���FM)�8���ӵ��؛o;�~0�C�����I�'rf�o��>6<��>�ZT�p�yo��n� �Ϲ���#.U� �v~pmƁ��3�X&lX�Wz�=�]��X"\Ɩ6O��B����d�q�D�!f��Wc��Q�4J��0�f�?��=<�7��ָ#H�#�y��C�K�<̟,�w25��Y��J��_h]�#� ��^L�e�u�����r�fe�c��/��ʩ&���%r'�1�iz�Ep/m��E+̏X�0&��`o�5i6�G�w�+�����Peu
j�m@W�����2īl,��\L�T8�i��3-�0�����Ϫ΁x��t���<t��eų,�r�	��S�!'~�Z�h�!�ۦ�[	���摀6�K�g(����ZY�o�c�X��ں,��K���E@z�o�x9e��;;�v��PS�aH�KC���J��|�4�K�.���סu������_�GL@l�kU$�
-׆w�}�`y*z#3+�$?�Qg�!J�2K{��2ÌU�SL��C/�6��A�:��K��d�r �]3+3*"I�"��)��ޘ�(|kQ��vw"u���2RLD�ĕ����&'e0��2;�_�"���Z�)mC��`�:�'f���$������9�ꨮ3J��K?���۴�MD�$mư���nFd��A���_U��Y��~���V����m$�5�gzʮ/�,�ĠB0mm���g�r�_R���u�NW!Grz7�#\�EF%��D��V�/4��^�RA<���h-qߊ��P��c0�ƌ�� ����3G?K81��H�1��U�rN9BL�ϻ��}��zr�Lq���Y��J�(����[�p_���1� .R�����L ��(���23?�����0]AΡ�WĥET{�j|H\[RV���HVj����	���CU���	�qM�Q��k�;���j.H��x���=�oī� ���*���䵈r):;r�K?v5�?�G��U05���vE\�ڡ'��a�-(�&J�-H ���F�]tB�]D�i;?�S�^
0QU*���jc.ʱ���kt����p�,a���N�X><���
�}z�;��=�4�)'®��t�P �kwY��Q�\�߽o�O,<������$�?�(MbM��� RڳL��'@�Y#�����!"�Q$뷰�����s���,��ST:B��(���F�����
�=>�����G�l���7N�k�|	d��P	ʄ�K�Rz?�S�R(٩�8�%�ىU�o��,�(%Z�ٝ��(38f6�Da�zֶ�4V��-��D�lؓO�R�᝸��z���;�3�Ѣ�<�&abF;m!�䭕����rw��$إ�M�a�5Gxt����������R	����w�Kp]j�d���G�+oo�J�B�s_�Jr$���s�֣`P\�P��_�mv˫
�3��C�4tA���@�a]�߫2U����D"s��+ڽ{&G�D��kkW�H��'�J���W�ѥ�V���i ���A5�]���D"K�l�Xz
^�׸,�0&ps6Q+�>d�͌��1f�ܘU�5B���s� �����7��fv);SI	���-��JCg<�6�֙KR�w��Y��h���&\�L�sǧ�������B�
]y�A�3
h{����=��E��f���}�G�eN�^7���ٿ�K�uC�`���Tio�'�5���1ɞ6uh?���:d��E�L��P�gR=��l{���Q�O�����#R�Z��ĝ�F�%qkC���3�SUJ��e8^��]3ӟ8>X<p�Ur�C��0��C@�j	��s��������|��J�G�y�a���jdoσO����V���w�ġ4ylU���uĠ�N�9o�t�G��{�DJ8�y�	Ѿ����t������{|�h�ƌ =�]&�a��=OB5�G�K�E�}�۾�����}�qAq�Z|K�[�^
k ��H��6�/�k���.<^�����0"����x z��<�FbjA��۽�mX��m���� �hVRы�����
�浪t#b���9�ķl%'�������wA[���[Ik}��r�F��X	G��  T�^oMc�q�yZ���;��U�3�a��B�d���T;������{u���<��?9���쇕�"5�k8T�F�ARl�#IDh�8g�C.���ֈL[R��Q�A˧����	,k��%�u�u�V�IF�u�,�r��By��6���1O�$���c�s͞��Vɾ�}������9�^bP�2���6�Ϋ+��79bj���l�X	���l�SJƃt�j�l�����2�u�'Þ���֓K�2M�7��6Jbd�X��Ό�#��2d�� �k�U���@p�ZbOa��w���CJ�{�C�vA"���)�[ӀmLQ��G��(�E�CЏ`�G�1�:���P^�����-.��@�'��s��cI�J��^�-���ⵤ������CT�!��>
0g�2�]�P����3���eS�b+�o��Q�5�}%�}�˔h!�>�s�u˂��G\���bZW���;>73�U�� ����3�ƺ����HXN���n��a>�W"��+�P:SK���L�}:4��Y���s����=J��x�*T��I�y�!��o,¸�R\í�YOJ�m�!��7Y���x�Պ�Sw,&�NE��z"�[�ܤ9@_:� RE�΂Q!9/����ȊQ� ��7�pv�T��WV���D�`������at���"(ǜ��\����_���rSӓw֞������^mH����5X����ًD��C!
s��'Ȉ�
�F]<VP-����`:�H �`������%�e�P�	���k�L˶4J�ʥ]���t�nlm�0�ޤ���_��&�{�}��j��P%lk>X�6}�W���Q��ywԤ^ImZ`��93'3q�{��9Vt䩕���⨍V��Ą���#�s:2�xҠ��>B����D+>4��H����P�!Ws����,�X]_c��~�5�$%Р��A��[��fbvFM59�Ȍl�I�D ���Ͻ�g}��`����S1j\�f�C3Ɲ��q�U�0)X��w�fh��U_��{���G�ʷ{��!��J#��d�p�=e܉��3���F�:���0��u�l_��s&�$��ݬ:���^4Ȉ�Z����y��v I�� si� a'�����`,Ӷ��Y;���(�7aqr��.�2�m�:�QR�~��A"�WԞ^��emyͤ�E�ִ$��j�Dc��xq ���^Q�.��a�������mh��B�` �� :��-��.�/и <v�\�ЉfT�S	�U������z@6O�Ӊnt{蝛���U�����C���RH�p�f*�+�	r>��x#��1��	H}\�&1G���j�C+m[��˛F]7=	�AX���,.y�����@%�(�e��8>�I��
y;����1f�`<"E�`Zl�\�띿�)$�4?aI=_m�1�V�a��d���j�{�(>/�٫��Ql��Z-X��i����Q�9�0D,�L�w���Y��V��M�z9���}B�dSɜ�^���ܸ���:�����Yi���<�(a��(�=-I?���	C`��8�T.�s�Wd�pN݊��}&2���'�0+P8����g�}�F�k�"V�7��9$�wɼ*�63�:��c��WK&��ۉ姡J�|bi���RU�i�Azvi�ؑ�	�0q)�[��hc���m>�zL��z������yC�����*�EMK��o�����zpxY�%_�N
� ���'%��_�Ƿ^��>��U���Dܥ���(�`-����{ 0�VG2+xF�WF�����Yʋi�Y�	&�������*�:ES�J�"�t�HU��`f�Xx�r1~
\����ε�K�sT�JwWt�!RI�� 5`�����(��(�j �y���/�/��&R����	�bZ
�w��[xȮ�Y}�Y���_g�A����V���;�:������?�ٲ�2�&�\����:߷��_�A-��m�0����M��JV��1'��4��m�̤�oi�ʙP|��IK�)�SU�m��W�I�O�t������׷t��0|Q)�uO���<2�C��^�r�j1����H�mHEɄ���o��E�!�zxS�+��6Ku�6*�;54�d����( �{�R��ܕ�v�1�:,�i������fo,,�����|����+��Pvj��[b���QX&��%����p�1(�m{m�������v�p��fҍH���K2twGP����w(A�Y�Us��}�$�UiKG6�e)���-R�)�T���Dq+����B�TZV��1�i��I!`5�T��&X�~s�C����1��3~��/�<gC�MYeΨհ%>��J�NnZg[d^.�?;�_R;؀�+J��:S4r��ȅ�����I���t��]A	}h�X(3W��:(��iI8 +-�Y\�B�"OOc$)�b	�*;$4íb���t!J��[]	�2�Ψ/�@�&���+�I�q��+�u;��p�!�E�Ii�0z-�g�[��_M�ӈ��oSW�.Wմ,c�G7Y��mT��)=N�k@�F����ۗׯ��
��������^r���6��ܪC��P�s/���t��uI�RcH��v��M��PV�h��%m	˻!�^P��(ύ�+D���̽���.T�0��v_h�˯1[_�}��ǀ z_`��R2�-�a�~��r�m{q�Wr+��1��)�n6�z��|O�5O�0�Q7���\�k5�g�AhH�旨0(��5��ﵺ	4��Jx�2��MzLgvDt�'�Xn�\o��!�DM����z��͔���3��r���5�fYb�Ol�hމ����\pPd�Z4J]ј����a�w������M��(N~��/��O7�>7/|����,?�Wn��'f$���z�'8�G�G�V#���� 2|t/:�jq�_���v��jr�{��_�N�g�P����|*�j�O�_4��`r/ A�D�t�`��1�q��fy�Č�v='�+¢[S�3(ܨr��94}�5�>`�'���/4�	�b�G�M�AڅX�j���H�?Ssv ɖ [wu��l݊QдCjjR���Ȣ�-�{��pDD��@�?e�����O ��'Ǜy�c�t!��5_ ��D]��z��P�`15IG�_��a����	��I+Z��<`�Y�����w�������� p���B}}�4����˫�ޅ�� ���hY]�R ��o�0Ĳ��Qo|�I�v�E��hO��bɶS����K�
σr��djY����q�9�^���s{grݱ�.Tf�3�R	a���Kl�~����-;ɗ!�0&<���0�#n�>�\��{RO����װ��M����w}�ͬ"�`�U=ջ�@�v]/N�yB|O�7D;�>��)<ܣ.�6;�/#���~KC2�磧�P�b� ���-�����ޣ'e�FQE*8P����7���eq2���[�������t��l� �߹ox�'P�5L��z���T�[[���)P��(�)���O��3�#�Qo�4���	|?ؙ����C�1�ͽ������G���c�A�I�+�89���6��{��h�>�L�L��̚�nAl{�����2�}qJ��p��+\?�=$���&���w�R�6 c�兙�؏���C��t�_�x?��Db�3/JB�� ��!��`]���XCU�EL0Y7��s`�f��9�<�z]��_ ��k�7�J^�W��H����5�/�Q���γ���u^��'����=���@��엺�4�[�����`�
 �d�jj�x���i��Y;����M_޼t$.�2��Iۀ�Q��j3��)1m�y�������_��R��k�
�5�����,ޖ�`"Gw�!
IK���5=�WXi�vDJ�0�ڿ�7�%h���Qq�O�0얀%�����t)�NsEk>4yY'lJ�Y����D��&%�LpV��3��o4��!���&n�~�&�,����MqT�8~ŗX�6��Y!������̓r�/�)_��ȋ�}'�y�L��ƥ�C�#3-�Υ+mz��NBM<�_�l����nR����Fh[���꒿��U1�9��aʇ.O�o�g	���d�
��t!Li�3�������G��*f�[_��U8ڸK������r�9yo��(�w1����8�B�e󢮶#�`\b�_�� �o�='W4���r��3�_�)ZL��y����K���m���1�Ϊ
4�6��YH`Eb�/�Μ�,I��N
�=	�!���J���|�)2d��&h-�C��t�����pC�I)�4�TV!��Bo��L
>I�|���]V�w_+p@�9l��$gck�z)a(�N���Yj&ӎ%�&}5=i���2�Y)���y��5D@,�k�$E4{�����ڹ;��@��|H7I��h�"�i�-�v�"_i��N����RSpt�;�����u�=2�B)F˞9֭��ѩ�GWǻS�
E�<�Wٽ�h\�A�3��y+%��~���5�7�_����f��/��8���,���@�k��T�B��������Ѕ�5P��N�0t_����|��(O��Ojy2aL��и��F�핷xt_=قQb=��W'�5$f[h1 S���\����΃���Ex�a����q*{�.cͭ���)n������ɏ�
O�~ӹ�	)��#I�����gL���[���+w�gML���a�y��Y�F �to�lI%���̟H"�Th�=~����<�ۀ��h.�L���U���XTTO{5)�K��^����A_[���\�ck#[��J^J�/�s����ѯ���<��}�i���h����"7c���k��f}\s"��|�n��=ޗ�ڐ7������_Ө���58�G ���(�W8��Qa�RI����3f��o���;����=�4�LWzb�%Q1����qC���F�:���Z�'p��b��f=%d���*}��:�BB�p���1?i���u5��q�`ݘ��/��l��dp��)y���c0Q��=C��1��1��tS?
P�*o��� ]P'�]�q�,͎w�M,g��ީ�Be�������3�,��~e�ږD�5����w�������;����.��^�+(������:��?�%Ȑ���E�:��[�=�uA\&1K�9w����~W]��"�g��Y)@����>�F)᜼� �6�x��a!�G�)��X����y~ul{�,�f�]{��s&�^+��VG�a���x=,�:���
ٿU��d��`T�W�z��5��&��C�ab����<Ȏn�4`����ք����%�v�^I�G�$��UrM�껏4�urO���qtx��\����Si����_�N�y-q�E9�XT
�3{��8�������^JA��k�{}~�c@�-F յm%�gw��Xp8�X�Qn�h���`�
�4�/�s��e1���ΈNp�x�u=�Y�܃�\*9�k��Ӳ��{LKR!�x[M�x�I�팙!��w�@���пר�z��H�)_���������m>��SځN>Gez���r�7E���JJ4�Z-nD���?�~}�CWP�H_�OBtT�q�� '�}`����ם�t����
��jY`�Y�,o�@!�G��vyA�,u���E�}�6�#������h'^O���6�|��|�-faq��vf��G����K��9���
��j��qe@].M>�4����ρ:�	���IK�K<M�<L��)�ϩ��;\�g<����ZU��={�
�l45̀���a�ARP��9�x�yy��Y�X8i�0j����Թ���Y�i�� ����N�Au��{ԸP̥
��S�0����t��y�{�&9z[��HpJ�d�)��{����@H�S!����v���M#Г|q��5�x����C��`�o&�!�K���MĹ*\��fǻ|��F/:rXXs���H����Rhژi�w���H}t-������
&��	���w�A�i�W��}����w�l/$9��%r�b��`j<</�T6��Q�O[��z��砒���D>��Y�(����^1�M�mEKV�����:�]|TŃ��2�.�?x�A��ƪL�gUkb��[��m}�(>�e�Qc�=�hx0�}W%&@����E�:�
��S�Q/���˝j@��X��$�f��}�&�ܾg�P�2�2o3�&�6�5������.����f����e`���~�u��������C�NCm�dN;3�?�J�h��.d��M�57鳶'�"
8D�~���LB@����nW�_ �})̈��f +�WO��m�4�6I(A�CmԤ]�(�c\����'�W�	��v�:D��YHx3�\,V���=����~1h�߹|�=n�Ր>�ފ~�������8pz�/�'H�c�_��l��o�g/�W6J�,C���:t(J���%�t��lA7��f��@?�W�y�dīH���#E�xEJ$'�~������KT�@�J�?�riVď�C^R��i�Q�=���L�lݴ�Q�Tyo�ggɶ������D�h�m]��ݻ<S
&�������T�R1*�óH:ݎ���姎����k�_���Y� `[FV�j?�[�L_f�?�>���K>G��Y�SNQ����3�!�6��d6!�T}+�W�u6s.�ߋ+6�0�z�GuwfD�&,�P�2R{!�ۊbV<������s��o#�N��yv+K�.���x.��X��u}A���oz�뒜MEB���,�>�y�($��*��GN�x@][]	c����U+���'Y̥�6���~�q~���$���b����i�V������tw&�O۳�S,E?w�{�E�����>0��	k�aST�nj�1J��>9�k��܀�������8;(#�(�z����1p�lC'2�;��0����5)Q�ƹ� �W,��I*�4e�h��5T��<F�H�-+Y[m:*��Ƒ��{��[i�{��Q�l����3g~��[�M^�����8+5��������-笀6��
�W�>4k:/,W����c gC�z���iF���@�Hb�aI�ɘ�gܥ\�i�Քސ�u��6�=��t�����ɝ�tQ.TƵZ#_��/�J�Ҧ������'���M	?�?1��Žp��t	��~�zS��T0����9�$��>��XV�/��P���̕���8\c+���T/^<X��c���=U��@K~�@�`xa�R�۞w�l䳨� ���W�9w�q+R�N��-�Rk�f�r5�]�D<���WN�'2{$�z\R(���#�X�?��v��G�(��Xi�]�����H]G�Y��X�'���GHg�:��ϻ�J�7e�ݏeSМJ`�xfhe�Fr���vJ���m�$��)�5�2H��`�WL��=���n���w��7�?\{D}�0��E��-Ϙ����`�s3�Az�ݶ��T�d&�O2ǝ�5�	#!U��ݪ*:��,⨥�����G��F�=�[�oN<�f-�4D~��z0��Rsr|I� GN" ,�9#�g/Fh�:F��J�O=�	M0��y�F��<���3d�_��z���L�l��Tq�	`�O0�ą󹲁B2[8J�EOW����O�o{�~��M�;R�i�D�{�w �֭Kڿ��$��t�v�.���D�Ь�Oi�ꃩ���x}/i��|^j��_��Oѝ�w�q�	y��������ȵ���t_ ��{j��xh������ސSg�a'W�Q`��]#3*403zP:�����R����+�:�e�W��L�Lul>��J�)�W)�"�]����3�/�1D)���O=�����D�o��}� �o*���Q@��.���$/]E�$�6S�x��^�ů�4�KЯ=ˤ:;k&�W�u~������,�p�Ƚ�'��Ό-��u/��o31��Y ���Z��� �?�yrw>:��SZ!�w�w��¥0N��t0�Ӥ��I�/ߙ��DEXz�A(d'�D�-c<K�0�H�ߨ���~i�/�!`��Iͬ5�T���g����<�X�+w)oc��>��Ѯ_xV��<��GL��8�E8�2�8ƹa��3�p���YN]�|�ߍ>ǴI�\3�&U ��Q	:��i]���4��ρ�!b�z�W����Ɍ�~� ���U4g�ʙ ��o��������g�I�H��%�'�>��� EL�����g�i}�x�H�qf����D!�u1������C2�olG����􊵭�6
��^ 3��Fh��EYn�l�9x��8Ԍ**���FV�jzҝ6���i����)�����CYi��"��V�t(Y��m�-3B�T|D3���c)����i�m���.�����.�yϗ�0��r��t�r��,ɦ�j��+�X_}���r����GQ��#;`����4���@��s	��bE�d[�K�邛�<K�ц���%gF��s ��i8���68�i&ɚ�p��닟����n-Qm�ks�꫿I��Y�s�0��ZQ񙛃�骜1�IP�6`m�����3��m�hz�w�;��J�-�P:���m�?��syR��:�����ئ����B!����G�u�sT^��m�5=��N\�<���������t�"1RFb�Q����XY$cgo�Y�]�I<9p����.�c�����T% �R�뺤�CS��x
���Q.�c�#�!pb ��i��4w�Q����zy����i���	}]����ߞ	I�i�e��.f�iڶ��k7Ѩs:�Sj�X�^q�!Ɛǜ�iR���'�o'��G��@��T�F.���8׭���/b�P�&�&W9b��uMɄ��"^�8U,����|����v�F�&���Y#j�bjXimw-Z���@����J�70�V��[z�\8�v�x�ra��"�P`��xt�?��H���؜m�����s�\I	�k��v�QlB���n��e�8������ڂ��荼�-���H�A$���'@�����ckA�hj���%����Dc��+��P9j�E��S��CUfj\PE��?9!�]�͘4�,�?FE bѨ1��#�P����^w��3��mn��Hm�
Ӷf2�b�U�O�[�#��$��,�K���&uDɚ�__"�6�4���VC}�B��=�Z''�`
�y�O��[ك[H�&��W��Q|@2���ٖ���Z��Q92
Yoc��4!S�11���@�������������,Tl�UQ�R�z�E�㲿x>ɂ٤�qA�]��hW�R	�����aEWla�Is�H���N�+s��WA鵖��$*8�����C@�+�I�(jC ��@o�i���`�f�io��vީ�.1K��	��A��u��tSi��,�=?r���"k��PW��v�6&�
���MPv�+�.tw��$L��E ���ovۅ
��Ѩ�{Q!�J ��x�9D�{�p2}��&7�ܹ>�v?�,�`4�䷚*�YU���=��`�����n����@��)	�5gdQ?h@`�/�X�T�
���9�SF������o��D�������b;���c@�w)���''v�eC��D �f����0oɴ�y���$2w�{�"�_�Q�e���s�<�D�>��Y�o��v��1��4���Jn��Z�?ї��!��<>�� ��䚸FUf�1��:,dp@YL��9w!��݂l�Պ��w�Gnq�?<�Y�V'�ߵ_Ŋ;�䮹�*�g���Z"�Ud<�F�s� ڊ�J4Ȧ�z\i���"��Zc}����������e4���?;������T��L�d +�/(����.VJ�y���ejn/E�HRnH~����@�yk�O�2��1;[�d�P���B@j�/ԡ\��jN� ���*�Ga�ʊW)�ݰ��D�����8��gC2[`��O�Yb��R�P�X����*�Yx�E�98\�d�쒿�F�o@�n	�����A��v>�=�Ζ&���`�9�y�w�4�����*�X���ol���j\��[

���b����C�GݣqO��jR9ʬ����{a;ͮ5� ��8�5c,)�~�<
6���wHG���P|�l]N W�P��o;��Y�������H�G+�z�:��=���M����������hFo<�_�f�'����Iᮨ����\�Un�	�`{3m�}�Sty����C��3&r���S[$�벪Z��Ŋ������)��i1��Q�͒� �J[���#5��
|
���*r<��r�]G� *���:��V�GuƱ�7�B��@c	�� b�{���##�� w� ���?�b�1���<\0 �2�̽Q��"�ka4kh����������V6� ;�ШZ���\z*�H�Jͨ	��R
y a�0�>`ԇ���s����^Xr�TO�������8w
�*q#����sL�̡*�x^��:�.3<���uV�xi�O��)5��uL4� y������S߻u4򆌌F*;�"SR=�%�G�%�c���`���Z�z����@�ào2
�S�]=W3*<�e� ��_�W�-ۘq��gv5��.xJӃA�: I��i��'��i�)L��e��%o�̰UK�;6����G�(ׄ��e!FNN3?}F���:k��ZdJ[
��͘�xm�Dܛ� ��ч��2��+���<'"��=ɥ~�+���<�Z	��ʒ����t���n������0
��ɠl3��eR��{_��������e���B,Q��27���Rb������d�q��JBN2�����V��A^���nAM�l�]��*����\8g�sx�OՊ�{�d�)σ�*�ݣ�6�Z�rG��8A��[Vr�&/#V���I8k˓�i4�H6.����E��jq^����S���V�I)e9�A�e��bÓ�Uz>f�	��������Rv����|u�}���W�5��Yc������h��^-=d���|b�N��$�=XE)�1Դ!�J��ޭgMz ��c,��x	o�1�]��<���dn��yuV X���aC���I�G���!b.�5�_$#M�>f�)i�����
2+5��Բo�Un��PG?�G���Ӏ>Y�bXI�	ˠ�1���������D�~��r��-�,��Ϳz!),>�=�:��B�<������0�H�	^�Bh��#4��.�
�n{��&�\9�����G�cض�Z�m0z��k����
����Jq�Y1����>�`�3�Ƶ�*�1�Aà#�0� 3*���ٞt|3��v
F���T����%ͮ����k3�ˍ81`Q�Ykh�m�����k�*�Mx�����+n�#U�z��7چAQ��b�L� #��i��2e>=֦o}���٥Y5mՕ	�pT] ��cm����L��Ӿ&���f���X��u��.n�Mtӊ.�R�d���(�
>њjx��lL�"UGcrZhq����� ��p���#��$��JR?���΂�ѸdZ}ǳħq"�J�|1_6e`�*�~�ſ@]4	Ͼd.�km��]��*ϡ��'`ٖPZ�UOF<�q�QT�
���&�A��!<7��;ͶѰ�}=R6�qd0�	dgP�$Ƹ��f�����g �z��a����h�:0'Ҋ���e7��ث��leR�� Zɒ��Ë����<(S+#�z��a5�c)�"�hGSTDC�����>�, t���4��O�R��4�,ē�R�����5�z�p�-�2�2'�MF��ݏ�O�F�p��В��E�����#5���S�Q����$����R�U�P�q�,#�q>�;�	�f]vk)�9���T㈣�)d>�r� ��z�0ͤ�~F�KkY/�8b��������ծ��N�tB�� ��+o�����t���a0��|-����L5�ޔp�DmPZG#���U��C�[ĳ�wȧ{DM��F%��VT���gl��訖[����1��YKI���Y�a���x�_�V�m�֪`�#�#�y�>,Ob,��04��L���d��+4Lf���zô6X�#3��W�c�P��2J&Z���0 S�JW�9�B�d���ݳ���B�}8���������p��L��7po�^g)Mn��.���tq��U�Ӄ��(����#X��N��Im��4�XqNw��ډ�$[NO"�B���a��g�`���]ݟ���X��b]o���w�������!�gjp����6����!�\�H/fH8	���UӊQ�����cϐ��,��+^;?n��
�0����
���4��8Qu��"�.�=����.���S���4���ޜ^uZd��6���̄��}h��U�u1��fѢ��f�T����u�a��~=k�ܻ'����-�k��}?Đ�cG ei�B��t�c���e^�Uw�+H���e�+��6p�X�0�2ְ��(���<����l�3�tC؏̴�2�2��V�m�(�쮾�j���� �a��a������<R��X��cK�ע� �>u��B=z1s�Yo�C�a�'c8�����N�d��5�4�F�.=�x����ނ1��-KۍOa�TI��GD{��,��i>�n�PA���`%��D�S�˝Be�#HO�ʱj���@�u?��T��V�4��yҰ����2�����c�:��/��dfy��;eڿ�,#�s�,�7�%gZ�:Tՙ�(sᚠj��t{���
��anN��n�n1+ɲ�~����tc��4aE|Ff<y�89��1�&C;�˛�U�a����n9[����aa�hت��w�3����Q!����7[����j�;�%18��g���9���������ɖyI?.��K��Uά���s�vLz�Wp����(����#�8��b������PI��J�gJ�=�V���i˹Z2uE��@6P�����!g6Y��ߎ'D;W�4����DY�Cy��	u1 ���Ձ�@k��﹭U=��v���c����E`y�^�0?<m���T���2lɣ�E�hu�o{H�fp�]�g�;���d�b� ��F4ԠqU��o���1�N�VP�����a�M����FN�9�wrm����B�
��P`+*6TSE.v7?o/I��򿪾��֖�7K��a�G��'��q�$ZB����L�w��޼_��]�&A G�m�f6N��먭y�h���{A��kHw�i9�,Ǫ	5)����
�)��?A�B��;+)����rxo���T����Z1�S@�P&��q�ׇˠpZG5̒�B�OЏ!�D���=?<ڶ�^<���'�.������	�N���-҄����=���!�0��gG<n��*�p��փ���7�:��	n1L��ϒ9.�Y촔9?�2��ݮ�4�~cTz� �վ�_���}Gf�������	r�aS�&�v�O��5��6�&�:�S��L�G(+W(`s.Z�����_�B�>ƯX�����n;PK<|�kC�Ԕ]8�����Dt�இ�~�����2�ob��8�d��1�Ұ��4��N�����n�x!�Ym�����d�H�P���r7 7x�06��-��Xwsmo����d+�����w"�b�U&����-��3)ƙ��މ�2"����r�ᒒ��'dm��̹��������s����a��Pi����84@��ٱH B�{��VnDe�#B����������󞶥����YU[u�f�ޥ�n��&�'6`$��NN�Ȁ�i#�Y?� ����y�H:-����:�os������s~cefڣ����W)�/,G�S]?W|�Y���Ex,��\���}؉~��/Ӓ��(�b�7�������A��`�[[v�iVg������
�koss6[NKMI�(�;:k7�X���vY��ӕF��0o����1���QW5r�g�����N0z�b\�����?�V��$����},�J�Z����m�p��$H_k�A0���r��Gd�_�X�����R��n�f��Mk)��153�X$�����Rf���v�1�5�B��������.7�d��˒�t��;D�uٍ	��H���;�e�w���B�'Ъ�]C���Kt�V���;<ى^��D0��%8�RF��ڿ����^Bq|���~o�7 ��C}XA8-Q��`���;��6���Q�h�QX`c��:��&T�g-^Vp�Į2��?��-]O��w�6����:_�f�H�v�5�����(,���b�H�x�H{`
���U�d�h���H,ɴ��
�/41��[l��e�(�BV��-�'kW���O[��h���]�i�n��;�Ƭ��̔�R2�a��P�r�~t�!K�;=f�[���aًJ��Օ��]ؽiM��M��`�F���*^�"��2^�e�K�X�Y�#���3n�����ӫ��Y�z�;=;r�F��i���W#��b~l(c�"�/val-A�)`���e5����zI?SA�M�Hܧ��	��|%mL�>��2����MJ�s��s/� ����!-�I�~0�s*Z7W'�yN}�ol�Oс�q>/���4��%�:\{�5������p�7�__�=��,	L;n��Eɸ8������XR�i�mf��K���3�l�uu�{M�u*�B����A=�#���B��"ڧ>V���s����D���J,��1�3�1O�����0���+���9P�<�ko�b����ELӇ�Ŵ���=�r^ɿ3���;���n]d9��׭�IH���<�d�S��17{�f`���>:�K$�v}�F��%pȸ��;�\��5�B���6���a�<�.Z?��!ںF<�/9�@��Ǹ,���E��c	Q#�/΀DG;���y ����Q���2%ʐ�ڙ�:"�l����}�������&����&n�Qh���7�kVu��ʃ��~HX2��+����!]�Jr��c���=C	0�~Ƞ5����t�*vO��1�D	
�;&�PGnZ`ڙ�_�<�j���J�9���݅�@�Y��U_�<�0=p[O��Vk%���l,p��X�e�ܡ�	��~�lR��M��-�{ߤ)-pE�q���8����&)i�*�Gmg�m>)Y�G���n`g5i�D�#�L̮�kŞv)��ވ||�͚;��?Q���r}&M&>������,K������3;Ëdf�tS+����@�D�5ow
�΃�����2~��h2bP�w�?�4��@��~�𣒔�0!\1�'�\��1ø�����g�~%��{�Q����wsTyZ̙om)��*A�0J�7��" 3���	K��`�0-{�a�y�g5�+{�M�����t��L�]��)7��!�ط�\�]S��I}D�E���{q�xJgN�H�;�{�4H�Fod�l�8����:לXA�2�f��x" �xٜ�[��j�"\M>�/A��SX�ꑊ���Zr�� (�٧�ȹ�H�ЅM:ˀ �]!�Y��DU 7�d�%�y��g��6��㇘0���(^�O��P�l�������J᥏���	�� 9�Τ狫;5s��ň�BήH-*���b���n`�nUGOd� ���fa�ZK�訐��*�1�xwO���]�~Q�����U���I����d���!�x]gʜ��ڌ�ѷbr>3W�@3��jv7��b5��ѐg�����b��E&�?�f�3���f#����2:����I��$�(��adR��	���)'�q�DL��X�_�2�Ӥ�)��=a��aV�]$^:�rQ����RES���#B���N�\�sE����p�p��Mc����LZ�7L[;�r�8�������%�{�p2OZ������n��icS^+LCh�+\��%�{o�2�������؏ʝ�!#��N�����m���Ӡ��C++��,��I�H�MQ�����צ��M�M��O���	��E2M�r�1*ٝ!��+��J5��|�5��yW��C��&r\}8��7dCt`�I�|�#��t&�M<%Ur���A��u=�P��Դۃ�n)��Ϣ�y��ɣ����b�5����I��8Ku�h�wB�;�(�6���r�[I��8I��C5�d�2߈���K�>�����)�t�L̃r�T�#1�j��l��7�@��?lp�<����}�!J�M�v��+�U$~��@�#�����#>��-���qMݥ\ �8W�E��3\�C��X@s�^�� SM3~s�1̓��Y�fH�'�GU�s�#*�uIԒ�~�𽢊v�X�c�wL��b��Cn*�F 9�����+�P��
5�����l���mU�}�2�=c�Մ�eR9p���.�P��=�&�6O��	��48�,Ԡ"ZQ�76����&R�u�����|w��r�L����co�	Z�ܦ�c0�O��zq|�S����$��y�~�ȑݷ\�l
]M�8�a%tPJ8��I�� �M��-�&be����],q�U���θ�E���s�\"�'���=�
�ߍ	S�n�Y��!I {�l�tRk���{R���B׀�\XS��Pb�0m-�9L_g�E7+��9�!u�'ύџڡ��x��>8ӈ��7: ,zqֈѣם�����f��E����,~Cl��K~?+�c&7���(�`����0N�F-ZDi��z��^V��qB�ѫJ��F��m���u(@�����<���M�sCyۗ
T�|\�H�����A��1im�?M���왅;�2��M�m�m(4�^<Q��u=����[��Ό�]^  �r�>=� �4/*·��Cw�͐�j�Jȿdoq�+x��� 1h����l��)�A1��W���X%4|��l;8=���mF|��Vr��:�?�f"���  Q%�����E��߻u)X��ql����pK%=�_2��=��e0�d�J���I41��1��
�^D��O���r��#Ρk�����x���Bp�WH�Z��-5��B��c�׃�O�3	���/�^��]����}Bu����#&�%U�C�!OJUw=}.*}^;L����=��V�6])>e�d3nϞ�S�:�$�P�H_�y�.l�J��������<��N\؈������R?iVz�%+�4%����q�qi7d�\�U��S��N�TA�A,Ϝ;���=6�\�	��{�@�d���Y3n�G�oz�[+6�z��^����1yv}̹6�(��� ��$�g�ė��Vv�1�
vi��XE=�qn�E0m�ͱ���k\��Gϭ�����{�v��7)>�Wt�o5����W�����)$N]���"-���|��12� 8�3�q�
!��RZ�jI��H%��zp7]��^���*�3�j_z�
;�������S(�{����p4�C�"<�@�0���3ˀ~�l3&�m����%N7�D���'zbqP�S��Z � 5je�Ꞓ����m.B��Ͳ�h4�A[�H���L��M�
߱��]�L��x�>�ElU��K�0<g^vo�[@�S�zK*%�����G�ƿ�l{�Z 0�!@��ݛ�D6��d���j�%M4԰�3C��)/�����]�N>J�E)�ln�w�تZ-'�c�w��ZD-��L.8�O����e����Z;]��i�v�O��e���85��Ŏ��z�D���� x�X�$��!a����H�W���톐u4� �J��q����6Di����&P&I�����"뙁?���?ţ�^ai����M�O�%8��_�UG_�T2��pL����%�:`*��ld$�?���m��RjM�>�_(�m�Ip�������}%�+K|͜�UW�����UDJ�\<���i��$��@�����c��1UQ����>�3 �E���K���r��-�<b����W����1\[ݑT�k�I(\�?K��[�s+,��L��c�7C�g�Pـ�1x;�`���Q��q䷵tz�u(�%j��b����ζ���U��`���Z�M����o���"r���&8[�:�y�Eo�;q��Ĝ>Ք!��{��A�¸۶������͸���R�\�!����#����ď�d��ϒޗ�,o��7"���sBAvc��_[_�6B����zim����ѢV�~ո{���2<T�+O�׷M���Ҵ�@f�$�*R��調wAC�[�F���N���(�,�1�$)�?�dZ��dE?i���r�����c7����.��B�n�or�Xw#GU�ͺZp�=1N(�7�J�������̀b��P��W>2��f�--t	r j�0�K�!�ra
��� wlir���5�_�b:`�����p�����=^q8���=׶	�~� WJ�ȘG�㵻Z �u �R>ζ�Ĳ��騤��\悄j�����*���މy8	9�c�*���1
�D�k4%������]���VJ�v�F����n�$v��Ɗ�5�&�W�����FO	���[���������A�n�(c�$^64'Ƃ'A��_���"��@����7����|��BUQ �8��@a?*�xY���$-�l0�A��X�\4V�G��6}x]=ͥ	���� DmY��E]j�^��J"��q��_:�C�ga�̗���E�8#�t���BV=k@\����R��el�<ư�^ᬒX�>�B�в�Fkhy���;%6K�p_#A��&Sp�D 
�*,Tq��$v�x.��/�sԺ�d���l
Z,�B�qgYv����{�Sbq����1�����f:�p�:E1�AlH� ��0�/��d�,�6��bJ�(�c�Ղ�;[� � �=^�R�6I*GMe���6�=Ͷ�?&�����j}�D��M�8xTQ"@��y�C.���3ϰg�������&xw��/[cM���{+ly�I����$��]��UX;gsũ�ͼa@cN-#��	p�x|zJ��s��w$7�m�>����~TLg�T�ُO\Ƭ3���h��2��R(*��([��E�A6e*� 97` $�cC�ֿ����3[8R� ]�N��,��)[ޕt������+�x�b��C%4U��hB���
�׺��Ȩ	�\��PK�v5�R����S'�j�ab�����N�� �M&Yt-��>�f7�y�.OC��Ԭ_d�I`������@�4���S��4^3*9���yT�/�<A+������*%L#�� -L+���)�Dp���諎H�F#K���IRVAƥ���v~��H�S)�����z�p(<A���@mj@�q�"�ˌ�[�f�>�bPl�R����,�ʼ��s�=���|'x��WN�3y�H]��ؗ<V����C�=�k!���K%|��z�C.�А�V�Z �+'5�['z��NG��>=[��ԕJ�ÿ�R�6sּ�`I��r�)Txu�L�O~i�2�}g)�!NO�-6�f�7����b��Q����Z�����'�I�5I�'J,�I�m̡��N���tA_�a߾��_���M��PAol�#WT�+8�W���s���6�;���@O�`7�'zm?J�n��|nT�Wxl1�����N�#NӃ��JR�c��N�i�]%�fZ٥?T��I��o�j�*p���T��xz���u��+�DG��9��笖%K���������L��:��b��e6�A�(��њ5���xJq�ӕ
�lbId������Mil��$u��*�Z�EF�+��GE�K~hR/?��5)��(�dHN���A�{�q P�P�~�Mg�I�9�F�w�B���!����َ��s���-e���$����1�p� h�����߉9����K��q	ۗ%ȕ�,#
͂#⑷�����u9m�\}�l� ����e��'�=N=h�-*�Q�YXO��8����V��^$�A��Ѥ�9��Rq;��'�Q��`5~�d��`��I&Y���t�0Nl�4��
Ų��xi�%�m3��f������i'����8�|g��s���J(�V��;D�Nđ�|մ��O��M#�.b
��b�%��0�1%��b*@qA&Ő�v'ک�����T6&y�n�)ZA�Ȗ��_%��pP�$�L���䔩��f�z��+�0˲�O�ӞSӏeom{L�r�*���ڭ���B�j��1�9J*&x��!��Z�c��A����y|����镮����B>���rdnW�~��`L6F3�U�7�BI����V�5��R�as�I(ߣ%DO|N���D�i��4[9t��
�[�gjќm���
଒���@�K%�B�^�G5��~�r-�^~����y ǜN�X�����xǶ5pE'�L6�Sw���zL��dJ���}#=�|�g�["�(���Ӻo�
M��-�L�b�(�<��T�.Z��襵�ZJ�;m������vV����%+sr�	G�3Bj���LW������ͻ>����Q�g��:���%DK�,�-�54�<2���]��|�[ �����:+m=ʈ���m�A�~fo�ִ�h�펑�FZ�K�c��h��]V��oL{zwA��-s]�',=��g��:?.�)-6���oUsG��;�<�N����B+}�m�8�8%3�T��d�خc��8��e(���S��ˌ�t�m%����!�w�*�e��a51A0{-`����괐�5��щ�~�hC�s���<v�Ҭ�!�Z� �{�S�put��#�.�w�a٬?��g��)�Q��V?��e>��"�I�`�RU����m����٨��g��?
IC�Q�;1#���_8�����(MOi���	��fk���j2��mw�T1(�4�OМ;���u��@�ַ��G�(g	��4H� B1�RE���X�V�О�x;���:|Ę&V����.����O?��n;��fH�6+;T��ԛ��&��J����1�>�,)����K�����-��9��[Tta�7T��u�6A�⁸��h)�Hk�����B��[�m�?�?���*cph,Yq<j�
��5�؎���ھ�v��I��QW�a`>g�cQ�U�-��K�O|�������}�h����!�u�+�O��������:i��?��>�W�OժG�M������')�O�J�?�=c�rm�j����[�Ż$G����6�(�+�0;��bE*�B���"%rkívz���G�������6ꉘz�d�N��L��,Y2�EE��KL�|7&��(P#?��}U���p�[Fy�\d���>a���t v�%��u�*:{�"����T��*K��'�S��$��)�S��7������=����d��]��n�D�Ir�����ˉ߃u�R��.�V���&��S���=v�ZHn����@�i�7���u�S�0g������.ަ���Pi|�1�҃����@�g�݅��T�?.$�B7��HbB����@��p�Y� ��P|�����kh(��GE|DxH��ӊ�̨N\UN_�ŋSS�� ]Ͻ��X)���$E��6�(����**b�>A|�L�O�{�߯�Q���AD� �zh��n�:l����9�zm��;V(,�z5H�y�����h��Xp9W��J�]w�?bhS��ӳJ?�D�[|���iL���T�Z�[5�u��%h%�;�ժot�"��K��R��Q�]j�J��T �}����R'U2��#
�H ��9��:\��k)/�ڌ�/�v@앑N�fyLt��w�����Gh���BB��;V�zs�?)��?2���{�ڭ�3�~'$��>k�~F4�</����=�.gIJ�;����W;0��-܎��è0�`2;�/��h���&���7B������2�ب��)�lf��/z~)W���$�[I�>�b.�	'q���
�ԩ.p��
�
 `�m����������J�^�t^^%��^qJ.À}����dc]��~����S������3���2j�6�nY�i��HZ�'�2�+��.�Ky������+�_��
���q����
��%��Ϳ!ɷm�����S'?�{�\3�-Gў]h4ݲx��3�]��4?R�����s�����b����^#jy�c-��rt�u��TO�D8��>^Q���о��79?�;]1i��MN�~�"�o)ƶP;�����֭L��˙�.UiyO$�{��\w���6�7�4~�R�����h��ǀ"���i�e�C���:d���c.�A!�d'l,U���1�Z�r��߀yth��D�/Q�{G��D����rg�w^�����7f
ru)Jd�j�	�6�X3�SN�rp����J�>岗*�5x�<9�2ޜօ�오�Dqp^ ߣ$����]�ݜ���,�oQG{�sB�2h<a��6���]7W�Y�8�t��~�< �$�ލ���7q�~�I�|�N��9Z��;��~��н'�DԺ�#�hDz#�]g5l�9] �u�˛�0'J5A�X�2 T-�9�0���!!�������լ��S�w��$j���1+W�����t��(�F��Ȼu�L#p2Gv'�� ���I�������Oj���n�tJۂ�������0���4�:)ڞ��{��� 3��qA�J�A���SE0M�����������O�i';k�:x dZg>{s��?�`�oqF$�5�A�T-��"����<R� ��Htp���>M�$I�9_=4�^�����hL�n��feZ�U�ʤ� _�	e�U�@�a����_�
����O��`���Ey�G5Ig���.�����0�|�k(��x�%	��^�.�<�D�:�.x ��VB{ѣ�-�_��.����t�_w��D�Y�atg��r�C�
|��zΟHo	���u3�JJ��4r�!Szɴ�s�xԐs-q$���ȭ����Ù��ǵ^N9�?���91�y_�mU
$ _0� gU�����]t݈�s�)MnU����ۍ�0����U��W� j!�q<˭[���Ir@I�ӟ��"g`�^����/�W���1����7�(\EJ�HOxk��~r��D�wi	mC��ɤ��* OSt�"���\����v�@�ْ�����7��q���>�'xW�;*U�����E%���?9*��.5R-�$�6����EӲH�N�*�ߒ&�z,�W��m�zu_J��>��O����ko��߁��hĄ�S�Hn���������س^d/M����1Ih�M3S����^�5�ȲƔ���f�%��&��"��F�Se����RU	�L�"WO��NƢ3�����3>U_G,r�=iU�m�p�[m�eI����q;��5d�tC9�n3TvUQ�0�?��0N���O��m��x��2#�t��'ݰ�w��g�H�XIBx8W��C�"�@ܻ���d~�y��ݐ-�Ea���H����okKEO;��S�p��E��d&�3j���8�����s�!X
�&�:L)�v@�S��x�y��w��2�X���m�I!XT�J�h*�zk�@��
�B�x;Y7���]1v��gNOMXO��9�e�S:�w�q�SмҦ��kt��ZA?ɾO���~�V�~~iiIL|�0,����& ��H$s0����]�R�����E�LD�V���\	K��3J@���v�(�*O�#/i�y�&�g l��V�ێ�B�K
�}Sh�ua{��C�9��U�.v���Lyv~Z�戶��Rp����A~��ӌ���#pi�i�˩�ڿKKC+cmj�}�Ϲ�<Kўz4n���6��+s���B����z|+rⅦ�떇��흢G��R0�f�!���cU�'=����x�`��(���%����,Ģ=��7$VNp\�W�{"���d5E��(�/pcS�sN��I�縡��P>��*��<A\� �{��`!�������3����sN���y	��$�nI�2��G.��ɘG�N�qY#;�<z,J9�Ǭ��!)��D;��V�1�����j��Td�R���W��"Ɓ�3�+P�`���<p���7T�>IN9ѡ�crUe��H�sm��y/׭�c����B��O��$�����n�RP�0�}}u}Y�Ϋ��:�޻<hszR���/Y`+��i�%�}�R����q��)��i��𸤉@�m����J�h�C��T���F]���_�הy�п�i̎���ƶ��^�
װ	=l&	en��Bl8��.���A��/q��QOU鬗�3��,[sM�!�B��7F��G7���ry,��iﲕ��X���7����g����A�B�ր�RP��I yv�գ_�s��vLƱ�Z�eD��
q�^���އL,���m��z���ݖ/h�|Q'tN�B9n�����H"�x��*W�J>����Y`�ì����&\�/��*LO4�����O��l�� |E��~>n��'�Ԉ�=��|�x�au�J�0@%}S�O�s0WOG_�9	@Ѧ�*3T�֎���)��>��x���,�����ik�.J[�����@!����RU����}s�>or�3^�����7�%Ԩ
��.�G��U�cUEmӜ�Lqb~�s���T�z�X�_�p_%_� : �c�-f�>��0��z9���l�KxJm�[vQ��s}�5�Ϙ*`�[H�TG�,q��D99^�N�����E�����~$$�B��a1����ܢvs��B�4Hy���D�Bd�h���k>I�^k#���x��x�φC���&㊣��6 N��`��i|m��ߦ��e(�~�4�Mݣ����Bx���f�듸
��i�留�(����E�O<�@�k���v3�-Ȁ�ѝ��o�dD*s�L9q������x@%�>��4щl�ʀ9H>*4~�sk�!�9�_c%0�M��K��Q��y�׵�(䜳��x�����58�c�Y3�M��K��Hg�*;��M�0��W���}(IX��=#[���T<�vP�{ń�X����c���ŀb� P�9��.|`s�Ӭ�!	e���!���#�"��V{�%�u�W(2za��=�u�D8"��Zg�QX��ϑۣ�;gn�|OՍmI�Vo�,p`*���M!2Ԟ�0���6�]���4O���3F?�B~P�
�(��fy��0#HW��]�Jƈ�8Uw'+���DP����vۄ8X�l��'�"vqkkn	T�7�;3�W��傌RX~��ϗ�˫t�H���J� ޝZllQE�ȫ+?%�1�!�1�tM�*���䟗���Gƥ�p�Ì�1Q�
u�{��b�5Ɵi���t���q��>:�6��4�u*$P�%�"��N1��-_]��l%�AMT�*�cQp"QE�l�+X����;��6���C��]*g��s�^�<Z��k>E�>�eB���g�Pd6+G{MC����;�M��.�L�ٍ`�'z�����uO�KbzHE��.���*&n�2r&tzh��Q���Y����bQ��F�U��8�	3rN�lbq���2#e����y`���&�h�xƆJ`�>�J��53�sV� �{V?lYlÎ40g��^�*�&%}�d�,�&���#�^֥g�4���-�QYC����Q��Ko���Ȋ�C� �Bb��o$�\$?��0��z���!w*�hS[�H,w4��Y�f��;J�K-�g�	!��4�0���ztZЛ_YC-Gr|ϻ�<�"Vb! ߶|E�#.c\T�q'/��Z7��wS�w �%3�ORut�fA� ��S\hQ�~�L^Wt�a���9�^~�c_���GN`�A�*Zg�JF�t�(��ory�.�_�*��m��s0
�C��74����r���9����˅�˽��&�����r?�	*�(�Uxr�
4�,y/� �� �r���e��C����y3�#	�{nIզ<�!���;[L`3  W�Y���yX�jiSP�AW�9����O�8��L����ݼX(����*_�wa\�Pǁ��3W1A���$�\v���#͢�,��ei�a��N�AL�^^_>$�� F��&�I��l���G�-�n2�1WS�B���]&����3����?�kX�D�sb����M�`L4ý��wJ�ʶl��6Z����^�D��CG4�_� AH3��&"��s��n�Hd�V#fЬMS�zP_>A=�L%#i]�*T.�xW����&%������]��a� L9�tށh��׋�������������O�Cn�q#���^1>�jK�v�N+�foi����_;��$h�zpPmL�؋��BD�M;���P���B�q�ߤ����4vJUE��e�p�k�8ӗp�B��?�^s<�
'`ϣe팃?`�����4Z�;�>+��W�Р��˟oi]�O���K��g��B؇����	�U�Cj�����}X�k��,�h^�c����r�I�e(�@JПg��tQ�	�@ҕ�곻������=c�.�t��=��vFA�t���f�h���iO&�o9gn�^�V�Y�0���Kd��n�I9[�1(X��Q�^�t�2l[����� 흕��0�o�t����B�Άn�wQ��E���O�u�RD��씥���*��5Ϯ9}_�� ��s�(ՙ&�G�>ڊ�y�,���G�j���?�Dt=`PU[q�{��9i]���b��EE��*����h	�G����K���N�`fu�����~�f�_�kJ����1
P��} ���������ݓ���#"�넳uW7��
�����L����������i���gχ�@��0 "�7Y��O�ۻP��%��� �7M�R��4;G
wzM�'���<�e"D��s���,(�&�qt%��J�b�V��m�	Uk�f�<@��ڀ�"YN���5L� ݝ�6�U�`�B|pT�`s?X����?𚳕�\Z^a�s@S�ydQ%wz���uBE��{�ҹ}*�h���݉]��=*��B��$��I&��a7�%ħ�[��rSC�?�vV�΢��Q�VW#V�s�-�=�(�E��7��E��	�l������0�o�.|)���\��4j��1%d`,YJޡ<�`¸�X >�,e����=ϡ�z�D�8u���b�����L@�("A�|6��������2����B'��v��e(�	�>}�@I
NZ���N�4'[U;�Dzh[�0\��{ܭ�r�b���U����C��f�̯�T5d�i]Gߒ*g>���E�u�R Gp�R��+���)1�_�c����<K5*$��~���Ww�RgK����-R���v���Ċ�%�J� ��ZGF�D=����� ��y� ,#4��+em���R~.�,�pW���䖒�  [ϋ�ᗵ/]��I>]�ܶ
S����:�?u�+�]x��T�<�4�P����&�ֆTI �T�Y�_���;/��Ӟ�oGW!������ ���v<Y��n5Ǔܫ��d�r(�F0�u��*�t�8;���!y� A
lQ~̕�,n��Yz���+�0�C3�E�y�I���t��6�ۧ2Io�a%sq�t_��*h��Vj=)���>����P�*�R���`���*#��(�4ɷcs_��<Af��.?B���0ݸ���ՙ���ibBl�^�na�ן�
�K��U8��%捹/`_���2���`UeOq���MO�QL0�[�r�s�M~��ӳ������=G��qP���H�Y�]-C�v�ҥύ�=�|u_W�-s�f\"Ϧ�6�0�[{�$�aŃD�U7~�ɾ�w�6W+���U���P�ghh���xMj�e����u�'�
��F�`�Uޖ�ʃ]� N�n��z��|������OAv�JUO��]N�����$Ǭ�:e�ēb섡A�s�"��ph�M�"#�ꍉ��&Ǹ�
�%��	�Ռh�M6�h��a�j�r���x�˝hO��gBO+�R����,�!	,wa7d�T����KF{{'�l����'�WC�t�@�H��i#�Vd�L�o���Go�~Icȷ���8b[�ڂ���"�nIT��@��y�+b��P���;Ռ�R�(�ɔܷ?��8 ix����lT�C�N\��D���2��rߏMQ~��/OV$i��Eu�k�}���ގq}�
=�M�DQc� y}hX��K45�:U?���,�9�g�md�=L�~��-�UJ��9S'��s6�	�!�?��Oǹ��..�)�7rw��T<��zBǙ�w��h��d�j���'���0����y	��VW��4cTb� ޑ	B.��%F��%/ŞL�894�γ��pF��?�����aR�t�gm�0���w�>�;1�7+��R�QB_DR�>���t	��&a�lխ� DO�m\	�4� �/r�y�)��|���es_Ў�s����5��H�j5$ʄ��Lڳ@��耪�6��8��7<[����ÊJ(�]=���	1f��d"�6�Ƈo!���eA�oPذ�C�������me՘#�[FE}:���U�G\��V��P,A��+m=4��.�"ߓ�fM�f��?���H|��2��LhY��yǳ�%l�A�l-�,�Vq��*\�bȎ�w�o,8d痝_Glu��Y{C���,�aѷ���n�Z[~P�����u����u����D��Yկ����d�W�;��V�6��Ok~0e��N�VR�9���Lذ���ۘ�"��|�<I�J9GLﱫ��s8�'�:#6Y�b��J��_
*ce��
僑�ǳ�N9ƋGv�����n���;�bl�sϊ�����Y�c�P�O�g�6yr|��-���J$�Ok}�z�['�tP����	��)�7�ι��®<���ٷ��U�*\v.nx9L������m/�U�m+kƆ$�f��z�v�ۧ�2�
[X�l)f-?Ӕ�̏�������s�'࿶�x������8S���hz鏛���%c���f�}�d����K��cؠ��d..m{��Cb,Ԗ�:w&�~ ;h]�F�qn�mT<�1���˺�J��n3���r���m�#[�`,Z�j)��s	�M��y�ʄe���U�5���� b�w�u9?Fr���4?�-0̫<s��V�YJ��c�
��SiA{���7O(��ꚍp�'�7j,͒��G	����h��z��ޑ�8�k�u�m@�tW��X($�`��A�� ��6r��D�e��]����Q�=�v�)'�b���.܀ć�cBL ����q	���3��c��g���S�T �C<I���;��K��ɤ� �NM%\��\\�'R�B	8�ۓ$a�JX,��Wyi�f�Å@f_�B���J�~��j(�u��_ʄF�s�Au����u�JK�� M��!F��{�hx銔)��3���XQk���J:ܞ��?nw(0�?/�&(��@B�)m]�H�2K���s��_/�T�v;�!�G�Ah�V�SLȇoj�Dqrx��a>��iڑb���r��߭N�Z;P����px�YY�\��Kd����i�� ��C�d�d���X�HU,M�@0�b�[�uÀ�G�hw~ ��e��Zx�&����	R&O���R|�w��n���J:$3ɻ��y�Ӓ�F ��ϛ�^�p���N�_].B���.�;�ǭ��饡Z��1D�l�脝 ����C��F�B}�H����)=����}AV �W�E����i�'(7_������\h6���crl�G,Mϻ�5!@�D�bK�P&�A������i� �
h�T����*h7��&;�	4l���ĵ�!�nJ
�Y�a��mj5 E���\N����OT�qv]0����#�JS��I:J��
�X��s|�u��p����3?P���¨�,�`sDG|�%pqbS&�&y��k)�J���0��ѐ��O>���gmi<��ڥ!gJ�8V����z��B��t9�6q#&�9����T��J�����Sf�����դ^U�	=~��2iu=�-�hg1x4�]�8}P��FS:Z��!�IM7:�1��	�Z��95^�b�I���=��.�lVʊkM�i=��no��'�`�8�LW�~鐮WI*��g���쯴�r��aD���w��j������Gj���"���Bm2����ޤ��Ï/�����4Z<v�oy��@��a��E'��JsL�Mf��DR0���ן~�+c4����:[�7:"Xr��� ��앾��t|U�z��V�v:d(�[Y;o���`�Ʉ������같^�D��T�i�Υ�S�2�4h6����0�� ��+lLP0O���7��i�;�:Q��pt='�O�8WtNf�y�����P��d�Y�Ͽ�#*�{�f��l����S��yI��:c�[T?v��uL�������{���O8�Y*v
��0��������K}�JmO)0ώS��I6���qY�0q�/f�����oy��e����S��7z2tiA�fU��L-nU��ZI&u�<�Μ	��qI��^t��E�c��<L@W��X�8r�1�oe=
[?{j��T�Y��' @i�Y3���o9T�p!{\�U�w�o�M�����1�h^�P(���F�����W���ٶ2n���J�l����)���HP����� �UϗN� 5�3d�s�s�������Hx���dOЋ��ψW*�-�^��Sb ���æ�&֢z��ha�e�De�{�S����x̏c�lC��
�Jȝg�,N����S0�F^�W�ߡ���!����YAY���z2�Ga�����5GJ�B�u��עo$	2�lGry!�55�_���9�2NN+�wt
ܲ�v�՛P�1Xd ���Ŧ�8��)8��>�L=4j"55����d3�QP�r�Yc��͟j(���o%��t	?���9�_���$�����}
��&n�hnP����1I}���I���)��̘(q��݂�K��bفe�����Ձ�ȁ�򌇸P��No|Tzv�+��d�+��E����A E����8�쑢$n�6Ő�8�)��iS�F.�X�6�ˮ����k=^�ߢI3�4uw�9H�X� �E"�(�:�1y�[}� ���[)P�)LM��e��j����w)�^����N��ն3�.a�oK��A����_�?~��F�2�.G������R��M���$#�u��"�Lݤ��Ѓ/(��q��t�� /[HHV�bkЏR}�4S!M6Ah�������.)b\�L�-��T�a�8U_��\d�K����-��Q����*����E�Z�o�y�U����J�*6��P�B��Q�D�?O�����1S�^��^�7��M��O�5����3v ��r���g����?
=:�T�!O�0�3V"iz&CE�y���<n�;���n�]��[���_���F�߱��}c¨�4*�N�H+Q����)٩��6{����r*�=3����N4ɱ{�Yz�����/�i�!>�a%|:!�Q ��[zW8^l�-j�	�i�\��ه�P~^�E}�:D߯�W�q����ө.�ͮ\�������$@B�{`��O�e��C��6��谟f���Cv״��Dh'�-��!n�X�uJl�O��A�w�u#�@',^|X�R��_�_f����'J�-
r��8͈��%��9�U��(�5�����G��t�i'X`+Z�C
�}>~�kDS�ڂ�;���.��C�������X��j+u��=Px-��u+�)�<�]�[��4Hzup�����XD�#��p/�㱨b����ß�B�~%�P�f�r�I4�����͓�Oxo��j)R_��UF���߂���%֙E��G�m���%��F��Cm<g���>ț��)o���PB>�F����@�E�@>/P�34Q1C`3b�Jw��b'�Th���0������z�(�P���W3��$E)�����;���xm-����X�V9������2��^�h�,(5��`���WN�{���/����=�P�.B�H���(黜!�o2�(�����XBO�]i'�l)uLѷ��S�Nc��E�	��v%.�X���{�7�w��*����M/x.��G��¬�q`�d/d�ύ5u?w�գ�n�I��	��}����ĕM��w ����6\7j3D�;2 Fb ���u����(�p��߿�*h�j:�n4��*s?���}�O�� ��>,q�B��숦������+�'�>MV>1�	����E<r�"|%z��w�Aܑ�PH�?x�]����.��Z�57��~`w}�b�\F|��fcX�t��>�:v�����r�i��<%U@$��D�N���y͍W�DY`]!E��MX߻��[l�8��a���U	�@x{	hR�]�\���q[
F����=* )���.�1���R����܉�ʌɭۥa��k���\�-B�LP�m�km��݆r�3��&&1�#���
��L��dP��?R�٧ ֩O
z�׿���e���v*���0����9�!Q.�K'L]e�\7����t�������aN?��ҋPd�9"�_k�^��[�=+rv��1`^I>�)��x��|��1N�p� �}��q#xe���R�g�ގ��}��\��ACu9�;��� ݡZ��#{]=�t�;{j먺}Z���qD�y�D-����*r{N�V4�@��!6�j�ԍ(�������;}r#���B�����7�T��:����"�;!���kd����#�S�쨒���bx�Gʽ�8��P׍����=��Ē�\��ԕ��F�́���|iwc��*5ۭr]y���ض����0\�����fӥ�����ؑ�v�b ��wpd���~'|�?��E�tz���0z��B�-`ҩh,��#��Ҏ�}H��{{�/t��wY�\rb�ږ.Q}�~dȶAr�a��/Ct�l�OR-̡��5�#�&a������i0l+@���So���b�N�Y�0Q�&�ʩmMT�&&��T�YG��V�Ղ��SW�)@����,�$<�GAwLbN�_�nAܭ�%��k�`&ݙ���(&)"ۭ|XQ�9��&���"A�o�PW��dL�јM�0���U�z�=��,�pPcVip$ln�i�O�^{j��.]3��VM� ��d��egO.m�;���Z\e��.����d��2b_Q���	tVJ���C���!��g;�s�~��ұ���Ϯ����U�8 ˮ|��[:g�p����)��X440�˥���mE�k�o�_�!بtk��
�$�7֠K	��/�ΙoYލ,�i�Y�Y=�"�I0|�8���c����FY]8����� ♃)��,�>'PJ��١n@w�*����Ha�>��X0'��9ѮOܦ��TayI�A��Xi�e��v+M8�;�qy˭��$�'��ʦ.q�C�Ql҈o'��'�#��`v|Se�Ք��p�E.��ǡ�*�H���6�e	��r���uem�8T�Th�AK_=������]���쁖�+��8������~���Y����8���R���)Ū,4	�0n�|Mi����I��ܭ�<ެu���x���`�nȭ�o� �gM|ym�4��4&wK�)�z��kV�<<=��]�@�غ���ǝG��Ѫ�����0�zS@M�Q/"���"	f�׀0/a.>�D�X��6��zv�c�+&/����$0�G��:��qHVG�b��/����=p&��tm�ͥl������(5 �XȆ� ��J���Ҩ���f�ʈR2�g��" ��э.�D�,���"���W�	ß���9%6­�U"�rU��|t�r�A�-�8�p��?�#�=�V�P,���Q����� Q�W���t�F2K0�NA�Q	?ޣSI��y뻠xբW-�anJ����U< �9��)��Rw�WD�~�7�E�ӂP��Fd8�M�pޓD�˥��D{�T`�2O>MM��L�}��O0��<�=Mm��:z�*�S��-~=N�a��M�TB,��X�{��#j��*G�&��w��$JI(�����4���"u���]���WZ�S�݄Z���66և�`(�Yi�R�!�ȴ��nM5#$�����&��'j��s�y{g�=�x���o���Q	���ꪂ�)Z�[2��AXz���O�R��ث����΋\�,O{Rr����J��:�h��#�|��������`<�8��\	e	5$��>SG1r�"T���/P��񝼖j,��kס���]���b�{�L*���Z��ª/����.`:�D�q:�xX��:"��~j�����#t%����V"�G[��E�UČ�8#7��q��H���%w���p�(�}�YB�
�6=�<2�G�y��*�����XH�\�$���9\`)Mm!�{/��q_�J�K/2/V ��,��ioO�{lO���t��a�g��_-���dy�6�D��D4��
�+�¼yNV�re�GZ��R���U��j�R�}�# ]���p-h��^W��W#	AR�f�ǯ��nP���^nǸ��W�E��@�k����1W�T�ӧ���:�����Q"�6 �� TN�H���`���''���x����a��o�19�<��1�~
��M�Q�<�BU4�!��u � d��}>S<?
#h�$&�cl��"�P��d΂��םx��j�<H�3��x�:��NKNӃ�;�-U�n��L���U�Wn0>�u���쁾T8�R��kH�ݑ-r��3>��Ct5N92E��̟��=?�xi7a�0�9���ڟ��iA+�W�7ኳe8 �b7.�[�@wIB� ��(���-9���-pv΄�F؈lH}����f�+�G�X\[�ڍ�E�@���N�!�����2��j��_r�����쒣�S}ф�T���' _�v2� ���x;��Z����Z�{��r�Q(2zI��."4T�􄘄��m�Bg��C�v�(��8�񾒢V齀ҁ(�ݯ��o|lLH��&����j^�o���ɺZ�I�T�C�7�������_�c�Zvg]���i5�	�	 �d:���W�.�T���o��{!��FG$�o����>�$*'��uP�ۤy���J�*��(K�!l�NA_&��}�PF�I�h��q���(u��|b���)Λ�ez�!H��'�̩�kߥ���B����]I����;,���?���T�����f:���h�,�UN�V�]@�\a۠[D�^�)�f.��_&�,�����kt� �r���w�-Z��0*� �x|X�.R���-ɻ��TB�C���ҋI4XN}Zm��gԉ�I�j$SϮ�<%	n{Ù���*5�HH8u�K����
(ӧGвs @{8�w>�+�4ٺQ-�<������1z�͇%a'W7�wqD�jF�ʊ�Nh�n�jG�((�]yV-s��ǧ$k��<`?�`�#�XG>.���=�_��`} ��ȨZھA�r�.?:}�n�G���""VdЦYtmA���H`���1E���d¶��;E�=�G)w��eY_͗���Q���Qa�G&�퐴ݰ(j�H�6���?5��f�KI'�Q�Q�������4.��%�?O�Hu���t���Ӭ�␏\�fͯv�:e�viq���9C�ޢ�SB(�pu,�k��DX�9T��j�&�i�z�
|d�W�<P����ϖ��%6���Mx��łp��΋uѕa���e��1�+�sw�{�^����c�4�N3+�|��T�f;���� ��Һo�&*vY8Ü��}�;j����G���9�*�$�̼��o�_
F���M!��o���[����;ǳE���I�֒)B0쫳�	������o��/i�p�q���{9\��0�0U2S�T1������J�0v��fc� ����D'F{��=�)�Eu�������x��Z�xl{����6d2�Li?�l�J��̜0�ƤRkpm�D3�yc�}��Dh9��Oz��	�t�a��K:����&m����*�=��o �������%��, �1s S*!d ����.���0UuO5Ҫӓ��Y��
��Q�(̮��$7�"��Z/��ny���p����Nത޵�{|f�c�aG�>J���Rl&>pd�� �"�g��l�QsV�V�X�v�C)b���8�5�\��SܮM(�w/��V<H�TWrm�E���5�mJ1X.�p4�^�iD=�U+�AN_?�
��E����^B�@�S�c��-4�{�c��a�I�d�"����K/Yp7�C]܀{
3�؋6�xn
�N�h\���ٖ0r�c��&��ح�����_�6����k��g��<g��,��?��B�D���1lHPZ�	+ 0���=�qM���K�&C�	��B1_�������z[w��ʑ�P��6�2� :��N��Ӥ�"�>���`�g9�X�a����eѦ��o�+�^�䱒U
,���;�3M_� �^��[���c�8�]3z� B�J�ЇrHh�C��w���A��N��LBz����~#�\�W�:s�E��2�� �)�o\����4A	S���7=��6�@�h+�������"���F��s���sM Q	�̖�Ӥ�3��`Jg
~����ej�^Pf�OڿѮ�� ���k�U��f=��׫鴙��}�v:T٩r�P�ѿ9LJt�����g��9�{UD�(��Խ��ǲ����$
�z�r��ۛV��,�+|�,����B����o!��ʠ��V3����8�-��	���c1q�2S�Z�����8��( �zhc���e��ƣW-tp},���)�x�2�>�(���"��h�"4��49�>�83;�f�Q!��Y��$"�(���X��_��x �_�#�r�xu<�+��m���>-9:����L�u�����r���b�c�4n)����r3�O���P*�o��{cM��fʬ|V��Y�H
�
}�fǩ�^7���pA/��Gp����5|�-�k�~�V֪�c_����~�P�6�T�8̞۪댝���8�Ǿ�	�R?��p���i����S��Th��s=�c�/MR�L�!�O��t��y� �i���x^;H_[��$���8�M�1tzy�$�>�{�e��Y��n9fGW?%sб�����쟥�CN3�_��dXc-�k�2�f��<GyM7(H���F�+82��X���# ������C�B}�%��g�����?z��p�r3B<5b2*R��Χq���ό�I����9j�*H���T��Vs���3�1�m�(��3���7��`Ka�Zj��S�sKޝ��C��ʳ�\�4�Q�H����U1W��˳���)�&]�"��v[~��8�����1򿖯;�,���4�J7�R�F)P�r�?�*k� R0��쒥)���h<Z������M���Q��L�s��WI(��ٱ =�`���ٲR�P�RqCsRe{��o�Q$=P��c1q�ϊ¶����?��G�Ti��'s`T.�(���d���>:��am�Kc�sÕ��z�K+!˝�:A�&�Fz�U9ȥ� �(C�hzZ�����G3���0���ً��mB������`*�xlJ^��8>��a�(�ӰES��McU&��hsҦ�`�����$��6�p5C	�o��ָ���i�����,\Ø��=<u�EW�)����k$U2���ofvKR�u��~-��^wl�+]/��>E�)z�Orw�r��D�
�儉d_�8_䴽E�~4{�����q|�-�����2��D&0�*�s| P�fv��\�ZMs��Vg�����{+Zs=�7EkZM=����s0�y0�6���_I�y�,�!@�xI��+��)Ϩ]=�v������b�V��� {d18�ئ/Ņ���	h�X��k�/\������}��Ĕ:_�Ь�AY@�a7�*�!I����A��m�Br �W�#v����߂Z���f+49����TD)�QgF�P��+��ɩ�~� ��2�J���&ZuI��˛�����$����M%���L%D��QE"Â�GC�����<n�3d�D�]���0u�x%�?o*����e���G���+�yn$@`�@�S�n[���$zc7����[LƇ�)�e�
!_���n��S.l��ÉXB�f��ZKH�`�j��YpD���h�	�	�Ѱ-�˖(m�O�����i�/eaѽ�S�i]�>Ѧ> �@����ziH�<�#&��t\�Lm8@4hH�����2���Ę tS�,��uv�)K;4{��)�������ۇ+��Q�%H�;f���%%�P\��0���l,�ڲG�V��	�1�{Ĥ��� ��P�c��rq��1w,�l��`�8tںu c�B��_�'v,�멫�ϋc�����}Nl�\�	�ȍ:��I�{�mR7��RoY�
x#��t�#�
�
��q���8WW��G�W\���[�e��"Zqe�
�2>B1Ǫ[d�SM��.�w|�>��B�sy��FH��,}<1��`@H��JԆ����%l���8F�6��R�&xOĖ[�����b�zc���s��sq�N#��aMbUGi&�zM��,f���MO"��"�q���Uߘ��*���0��?8�ǌ�	���q�&��X��r�cR���&���we垂+E��X�ca�,��2�/���i�x)-��.V��a7����3��nPl���͌�oź�y��o�y&��``m�<�?�X<�����Ztq4c��CBJ�d���y.�3NB�w�hL��ȓ��:�2���]u3�ϧ�+���}[
D6�Ba:)v�P�ʰ{�����.�_�S90JGC����9!>L�9X�=�=39tMY�H}AQ�5��矹�`�w9Óij�XbW=��q�^"�����q��xb���'����ZX����@*?K{�(�J:�"kN�e��yl���v0S&OPŻ��'����0FI��V�	�6�]nP�&ci�F4S���ܑ?�L���j�7�F�el�����)�\�S�6(r����6�IZ���D!nL��К� 0�q=5 6���-��g������Cv��-���`��$�9n!��	��ԂVK�._�^�/Em=ϱ\"z�I��i��ޛ"�ʕ��
��U��/j{����q�e�DU�}�b*r��;*��8���P�A����e�YE'�䪈�|��|��[���%��W2�� ��2��R/Ck����f��!tA�]a�.�6܈X�"[���;E>ҍl� ��66'A��u�>~R����3���~�2Ł9��-ģ-k7/_�׺�OBPXb��o]�&l*:q��/+Bņ�ϡ/���t�s�h�O��J$^I��Z/V�'M�3"T�u5�r��b��_M���W�O|2����Q~$��qT�L$�*Ч�T��F��8�ru���ul~^�7>k(��U=�$�a^��LϚ���B֞1���%�U��!�.�Y,t��V@���]I����.���Q�Z{��"�$<�=���ݥ�v��P�2V�Q�[�W[�\��c"���wL]�o������p���/���6VC�����f�ˇ��uQL�L�0�c��팄btogxH�S��j���L�&�l�������L�4Hmr�����ۯ����7ޔ.%	���,�����D�}tߛ�7Vrw�z��ʫ��V� ��膮�""�֚��oD,�����}��xNw1�T�MbF��gԥ�}�w�@�v�np=���\�-آPN��� �-�^Q��o�r@Z��ME�E�-��� k`���W¸��?R�
�s��dвg����V	������ eQ���fĎ����|�')`������#	d����H��Q�-��6:�u�Z7���*З������f�����ٕ(���D�	�9a����g)B[y��r�G�.�씎�̀�o�=��Ux��ρ-��R�q���#G	�8��-N���*�F����3�kb�E$URBD�Ga$ƛێE��r��8�4��!~������E��̣~�m�T��N�:~�ؠ��E���H^���|�O �oX(hst./w����:�>
ܺy7�f���S�>��ct�ۅ���5��b�������q��^N�풇"�b��6�V�
��u�_���K���oBQ�!��]Ʃ�|�lA�7n/%DI"��&i԰��T�А9�u�	�F\�;���ZHB����F$�z�'Z*��N�k}J��NڇЃ%e`}���m��[4nu2��͔6��zs.
�`O&�=����RHWN_���O'��UM�~y&��H͗u�V\������,�?mc��}������Ugj��e�����(�nر|�$��|E�I�&�+m���?��k���%�O���>v�9�+6x���>�)�5C��be�>5�\x'd�8p�4��q��?]�2��U>�te��H�ޟ��D�M��69�
1�^�K�w��&�i��X��CN���A���?��h��J������;X{��W�a�=G5����Z��lu����,��8�4�Z,��9���k���+�Sj$��f�h�C4���d��]��V�~���!�e���*�A�k2mEfx}�+�媅DR�q�s��y�&���3"&*�7��W��i�bЭ�:(�~}63�ŵT0�Z$O�V��S��_F�rqEty�_ۊ~v��c�t;ؘŊ;����Qţ[ƚ���Vx��/<�r�2�7��^D��x7�h�P���>R��^"����[�� KW�C̙g��.�^ּeT?�UZ��Fsh� W�A ��	�U�_�����.��ް.�+�����y��S���<�8�}m1��d6�!Â�(�m�\0TR�k�_�KTF�����ȵH��d�L�Ԇ����Of]��V��1W1$��D� Q,Ukq>\&H��Ŝ"�����|�����up3�����ٙ�h�������un|i�SY�����#P'B��Ƭ�绯���k �0O��	JSN}��ίL*�`�� �Dh�F��j|��}���v.�&�d#��*�l"��ƂU&IH�Y�l�f�.R������Ake?רl��}�`�:�0:.Ga[���qE*w� Wj�ƽZ�NJV�<��v�'�L+��e1t��7'��xv����.�������,����zn�x����u��#)���./I��9��{���ـ����]:�z�~�����mG��a4~����h�zgR�흙�V���iq	�����+�5嬝���\sN�A��+@�8���+
k����0�?�ז.�*�����A�;y�`���2�*D�3U�N�}��'�L��p0�Yv5��n.ߘ'��Pc��hM�s��pA;����L�@q��X��vT�g"DW+Z�Q���@}|���;�V�Qs��5���6��g1��[&���[O[VS�ܸ4�%�����G�w�<S�ՠϠG������l<��`c�<�<w���{�q"���b�ڷ�^1?��̄Y��:��7�L�˘�~�vas���Ԓs�(�
ӆc����N��A/m��T��]�l�I����ً�|������k��I�l�#|��;k1؏ �	7�ʂ��v\�&������S@�M�Ok�h	Lz*g<چ��n>b�3B�o�d��_�pv^,���� 2�S���f)��Vw{�s�1Q������J���3w����`��z�N_���mLI),�(|�������'�K1���Q'%�by�Ѝ[������Y�SZs�q6���{�G1���D�_!�J��T����7�w���.\h��� �#e��F�@���\V�S-y�R�x�RN��K��N���AwUТ���*�eq'��X�v˲�`(��y���G��P#O������}��e�qHL�3@�5�8T�ϨX��|��T�v�"�k�u�1�~y�ʇ'�t����f�����v�cM�3.�d�Y��WO_�-��E����昍���b��]���1�6�V�)��J�ޱ�`�E3Ix��q����<�-�����;w�?� M��̱���7>:)�֔�	�(^,KW?8������{λb���[&���O7�%;'����gCא��GX�*����z�����1$n�m��Դa�[��dp�����V~����-���Wv\|@BM�̪ܞ͆Z�p��χD,d�Kl���O��8��1ԣK�>4��;G�.��m���0u��~&�U����ͳb�K��U���]-rY3�
�'w�Mg��_"����Q���,ۊؔ`R�բP��D���J�TG$$CNm���W�l{�F��VJ៚O�#��2F|�/?�����g���j�|����z�!��nv���7j
u�������XqӪ��'��q-b��+�����7�k����-[̋�>��ɚxG%��M9��R A�9�P~�&��j�'��Q��דˢ���kJ���D���������(=�;���n����5O5%���= C�*'V��c�Y��l�j`̱b�wwz�h��a��9|�\�>�֓FݼSq�l����#�N�y۬�*�2V�8�g�Ӎc�4?B���M�%�x<�g"h#B��#�YJ�G�_��_���������#,S'� �����mJZ�|j<5ҋ�ـ���Ź�h��P�ӆ���{���8��ܹ��cԇ*Z�qҠ�ñ�OX,Z�t�N*�]Q��$zN?���n�����r�f�.��g�k!>@{�	V�Z�=7���R�IxU&�M�������Ѽ b����C�A�Ii��5�Q�P+2`�P� ��p�G/2a���&�x��)=�B<g⁯<>)�<�@c��1(�����Y��[V���C��F���6�t�A:Q���ŦG\�I���!i���=�q��mB�"+>YhM?ɽg�R��7T�d�rUH�	����U�,���7%�|:N�����/�G/���&�%?��E�uAW�j��c<�6�f�W�.�zvd���#�Tb���Ĝ �>��#G����o�@>�(c��4����Z�H㐐�x����]�Wl��/ǀ��zlQ  >�0�t�q�UK��_���Q�img�g*Tz�o� �;�]59�+Z����[�9Cj���eD;�i�k�C�<5y/,F��Z$!�A(��V*N2���V:ar��G��ǣ�� ������aͅ���۳hVp�S�� 0��s]]Dݭ�8Z7i��k^�A/{���Q�[�cW�;,�5�G?��A���	3��
aG�	0���m����'�G���~��F��c���?��q�=r$�3�7�_Y�� �6���I���wG�������ɘ5~ंN��� �"n��y�r瘽x�ĝ����S;p���rv���S�@��3�_��|]# _�Y!�(��^��Qg9�p�΍3��k����q�t��M���f��qI�y���Ίk+Z/��1�Z]b�M�P,����k'�1P3E�C�/6�?W�K�9̶�R7Rm��T�t�Q��MX��mX�������m�a��h^,Ն�C�_�,��':W��?���YgxAt���ZDz�LXc,�V��x�~��ʬ����iӦ���i,������4�l�s�ȅ}���0M#-p��%�h�>@��v$*�Hom�l�`d}�����{���s�*n��Uly�nP2�e�Pz�G��'�b{?�!���bA�4�X�VT<Gn.�9��0�d���-ra�����T�+f�1��:��伋
 �c�Bnu�,��t�Ϙ��N�`�%�%!(��c����\}N�v�w�������vj{G��c&�W�Xm
W!��^�W7&@�/��Ћ��fH�Mk��n��o0���n���k�;����
����av)
*�ɂ$%A�=П�ZZ4VIrUkO��3�����q�ȭ4sw"��*�.d)��;V>?T榀v+4!u���^�v]���u��b��
lR#6�b�~���+m$*Ϙ�\{���Ihx�O�Z.
��j��[�M�j��X4��D��^����zR��26�O�`��i��D���)��M�A��:���m�}�řZ����8Qm���#��f`�-R5��e%8	@�2���i-�����myW���_�n	y��@�-:Z��?���>�����;|ݩ
V��B����@#1h.��՞����ö>1�����Q/�Q����=-���hv�_�ϡ&���W��0d�$��̬�݈w+�������,c�{���/nD�eZ�_5��hB2;�F �69/I�HQ�� ��ޙ
�T��@Ya�Y�H��^�C�"�l���>�I�m����};��1�t�� ��up��d箍&{8)c���ɇ��:�ÿ���'oE32p,��rci�u�7��k�P�<_�oˮ �2��U�Zy&`��l����\!��@�l�)���|o�b>��l�Hl��_7�����V�fR�h��5v*Bzk.9^��_"�{�!%@�����3<�)"��9eR����~Zd��,�f]��v9�=��\~vqb13��+�^,�3�n.J�U��ӈ	����WGT:�%
�u�Ώj��$��iu��F�7o��ֹP�PerZ�-u3��9Lqd��y��^�0���T�w~.֩J�D��#؟ŉ*EQb]�q���Rt ��X�,~J�GhE�W��c7a���g��Tk��cH/|~���1Kc����=�����'��
������_ 5$'�Z�B3����e�|�/׾)�����]�M0��1A��
�k���?��Z��3���9�~Pa�ޜ�D�.w��u��f�0���'��`s��3*�{�nN��N�LL��!�,6���k��l�C��%M���cv&-�f��؍L�J�7yD���L�S�O/�Q��-+.BÙu�(��7K�YCLe�o���� kҐ�:��C�m�TrT��*��H�
P&j��r��R� 0C6�=PJ���z}���%l6�΂�1 b_���3����ƨ�
��������������^sj����0�����"v��3� �刷�d�&f�SDE�.ix�e�H��H3k���	���A���?����h�F�xr�r�$�@T4��*����B3A��u�$۝�[�1Xe�^2/ͷcv�����첈�0-Ũ�����~���l2a^�rHoa�b�([Е|M��!�4J��#��lk�/ҺQ�������M����k>%I �H�����&_j���[���a1�zM�u1'T44��v�ASAak�A��&��i$ĸ�)g*���J8��Å�C(6��!�@��sG��mW]}m_;�������� ��+vI]�T���u�rW���Ґ�;���i����u�#�Z�j�㽪���`����!�}DO����T�Ӽ>i��'��-���R�v���
�/��	���7�AX5�~4�R^��1�rgl���9�l�j���	z]��+W��6�<"J?ȴ{W��B&l{f�rO �o� �h�����f��1tF����G�r�&\3���g�c�٩��?)�+��KR'�����\i�;������B��s�(��h�?�/9	|��E&��l*���x���ЗǏ��S�{�
j;?�ҥ��*�-�Z�I��.��!ư��p[\�g8��j�����"�+]ӭ�g�WK�A��aC&3�U�
�k9$�?a��\y0gq�,7�J �4^��rPa�A��٦TPݢ:�����Yy�z䑰)�U�41�:%4�H������d�K47Bڿ�N�A�Ɵj��*�R� ugB���_�Mx���VUiҌ�!�~��n�ܕ�c�$n}��H�"�G�q��>���)A]Cr�hM�wg��\�W6"���!CŃ�`!��Y
);_��,�~ߞ��	O�\� ��T�t�Ǜl��vG��N����ƌoZ����ƿv�@I:v�w&��(?��I�E�o�VP�� pN�U�_�unn�R�����B��(�Zd�x�V't�ܺ��J=@���v�2r
�)`�)���w��y޳J�� _v��i�|�Y�s� �;�b���{�O�x>>Ǳ��'���9��^a=�]=#��EE+�=cOv�� 5�$$�2#f}��	?�[���M2�Ѯ} ";���e3@���
8v�po}��5��<��֞��9�hs�D�/��I�s��nE`Z\mT?�\�q	Ú����ŏO�Ƙ|�S��Ae�R����ȶ]�`�K��(RŌA�qR�_��FO�y�%�G ��~�|@|K�^��ȷ�U���u��K��AV���]�H�׋�	��8h��Wˢ�n���o&��em?qc��9��yf�R�O��WX�@�r�D6����NHIvE���q1I��������(e˄�q%$�!;�v}t��EKl4p���.oO`�}���Rj��߶a;i�x �jr'�mr|�G6;4��y"�p�tR1KT���Qc(=DA��q1,����Ҭ�ض��&!�<��+-0����Tg���)�p*$�d�q2�)���a�	p��UX��
�H�Y�ZYv8���Z�+R���'M8b���:��A#S5��A�G1\����f��W
����+F�3�E1����2�#OY7r>[�}�}�k	�x�|��D�x�2Aa���OH��2n܏@k �T���L���RS8i10�m���9c���!���M��� Hm|�C����G�_�A�UZ���fc^���E�|64��p�;�J�Q�/��Fݘ�k��AB���c�1�j��͟�W�J��p�\��,�Nt��f�#��n]_'D�k�O����ҁ�;�S�Sǝ:\�$� �i*T�����{ҿ!&"��I�[_���]��6P>ϰ���Î���<�v��^�O����������L[����
��T4"}ɱ]�; �v����U�6�	��Ծ�q����vP��%uG	���q<�\��/��yc5�o��'�G�K+.�z
���+?;U1$�H��e�X���)�ɘ�L���%y���xsDT[fo��v��u��3 :Ww(@?��|���\���CEMA}�� k����͊6����V��F?�,R�̒�#Rny>W��(Zܡ���'E�tl�\ݰ����	���ii4RP�f��D���*���U�(�7ʥ�$��_`��H�w�x8�}�6�Ni/\���Aa��]�6"�B���ɏk�8j��
}�B�2��7%BV�@�����S���u��8�G1Q�Ƈ+&���� e؛&  N�iD��kP-�V�ɢ�$L���B�<��aQ�>o�c�v�Կ����aSwr�.h��`RE��Dzg�:A�9$6�\�Y�g_W����-�Ȳ�2M&��<Xb�uD, �EN�:3%П��]zI�f?�~F�8+�,��6�!v/���H���1g�0�j�R�2l_N����˱��1��z��6�x�v&�0�]��7r�s̫,���Jz�-�'Ǯ*���"�,)�]r{ھ���j��}s���؈��P���#�\��!��B[3V�ǥ���E��C]�O�������B��R��RWQ�q���
���H{4�U{r�M��H��: VR�d6x:.��\�Q��P.�,w:M��1*���O)8%Og֭Hñ��}���7�+>�}�b��MOC#{�r���AM�-HB�+v�7�sHgm���q���E7���:�F��#���ip_1rT�T*XՌ�E�-��$A��PN��x��	G��'��"���|<3�kٓT-�"Vr"��]�q9G��N���͂�����q�=&�S��&<��y�� ��Afܭ�  ����* �����/���|y�)�VOƌ���i�����qEdE	�J�u�I\>N�/��$<�)��$�3>L��Vt�v�-!ٴL:{�U�.	���\wV��~�:�|��.c��O�m�Q48���|u�kLSB��Z�S��]�6��r�/8@`�򀳛����6��8���#QV| ������| �ݟ�#�W���@�m��C�'I0��ٌL�YD�����+�4O߮�����<��߷P�W9nJ�Ŗ ��=�O�L��ԹK�\���O#S�8'T��:����!u��zE��ٯ[l�K��B{1H�58���0c����W��H�}$k���E�+*jhz�^��z�x~K��R\_w�Y͂U�G�l#'�񓽐�ˑ���0�F��J�1��~}�h�J�&�5b�E�#3e�2��ȯ+.^�)/�4Px�~�T<�16_*LY�Mb����`�Zjn��N��3&��AY(�B)R��;J�E!��d0,'3͟���E�-����,6��Q�y�I����ilDb�������x�`�e�g	�P�f�u;J�)F)T$��T��K�"q�/������ABU{�A��H)v'�;��^�W������VX�D[���Λ=a~�/PSI<�W�{�thx�|��������������Ev{σ��
�@�/��ջω ��>+���^�:1]��YT���"��"������j��q�u!gw7�}�h��{���RD%];��� GQv�k�I��RPM0��"T�T�ם��|�>�&����U����$�S��'h���+�����=�-/u�}�ڜh�Ӿ�\sy�dO=���`�9U�;q���ZJ < ��o�	ǢD,��B������%[H����)E��L���ĕ�����O�i���l���r:�˴���^3�8�yȂ�e��>W���BE�vYh����x$�`_�'K����qh�H��	�P���sWz�H��}���F���������S��Z�:~���,�r}GHH�d��舭���,T�r���%a3��{D"ȷ���y?��P�o퐍&�V89I�X�����	ug�F݌�'��T�
ļo�{2�)����[���ј�}���N�?6X�Pޙ%?��*�ܑ�[�w�?�|Xپ���ڭ�7n6�������2�� ?�7�#�}��2*ͮg��y�MK��c�k:B��+7�S��o�1�p�D,�<�}���H;�R�*��C�O�Rg�e�b�v��G�����%,e�%�Ѐ;�R��U���=^勒m����E/dF����B�����]�W��d���Y��D|�d'����{n��E@+i΄K�n����΀I�
Q�܍����X�����d7%�^"�7��!�8�S:*��u�ڵ���/.}����^��=��ȋ���ז0�j���$VXsr:�zQ������Q�e:C�y�L\ʐ�T�[�%�}e�cIf�{?LE�l/����:ǫ��/#Y���`�̞⏷���I6�j}_$����Μ�qG�,
o�˾�0�q4;_�{㮫"wk�X�M3���P��A۝���H���`h�"� �`��m?��Ħ~ݦ���#0�0�'J�qV0o���H�:=2_���d�'��� ou�H�=$�͞J.@�r�����W��s�����#�ϖ�o�?tZd\�C;��8	����l�8�q��LH���\���ux��w";�`�nc�������Ӭ�_(,�8���Ie]�c��U2$�^xm�$�������g�@��5Q��JW�b�T�q�I�fiw�t�u�*)����T�|�7��sT�f�H+#���
1.6�� !{y�!��v�@><#���0H��O)��P�iS�
{�����o:�)�U�6P,����9GR�H�L�l�ca�=�5��w�Y�&x���WDv��P���s6Z<؄�T���z��/~�h�̫2��{�:J���q}���+� z~!�"��a=���C���Y���x-���+]G��X��6��� n�C�����9tI�:����cꎆ)��Ti-�2w/����v>_dYGk��+]��&��?�7��H�jJK��'���|2:X��y���f���*�Q�CB�-YKXl�Sd�,d���<�w|���a�N�u#�d�?Bu�Jo�bLeB�X�����i����)h�;�
����^5J�2���=4��wX�����Ш�P��څ��kx,I ��N̓�^9u#:�@ɒ�Tywz���h��Q��[���(Ɋ��������R߶�ht!�"�t�n�O�z���{@M2���[?;���w�`�S��-��*����*	�,q�D���`�6b��='�댳7� ����Ss�o/:���<�i���#w���R�����edIg�&��J��k�js�{�)���(; p��PKF�c��K{�2P6�N�=LF��8�I���C��]��{LS�f��B��eY��a�������qR4韘 ��X7t!9|��B3<Z����u0�&�����:�%�0�RRp�7��`��Hߐӂ��]����?!~4e�[�/��ަ�b���p��WTl>)r[z���x�ȗ���Ʊ�s��@[uѻ���%A
G ��t+6ϓ��e���܄
������.q[�VP�����"i8�1J���ǥIhS������
C\�G\齯�VZ�Hhr�p�u�V�*8]1��fg}S�l;Γ��.��4(<?|�#a���*'�~v��$��q](�qiT�<0�b���7Kݸ��7RuC���-	oTn�[��8����A�^����ŴQ�Ho:BE{'^c((?�Svӌ�\���"7�>�yj�2^�̓�ڬ����dX7"���m�$�%6�Y�h�p�&���B�uk�g��]3d6�׏��F��lZ� ��v�c�f|5*�]�/^�PaBJ���n��q�+eF��있	s��|�3G0��7|�x{c5f�l"`�jx|'��.��:_+YQ�q��J��&x�K�J�ߊ�c�(W�3�M���v)���	�Ɨ.Q�vx���;9�Ck�Y��\){��v�I�s܎��x0>��p[-�Hw��c��>Ok����O�Z
��Wd��ir�
����9(�C���AE5��g�XG��qZ�Q!�Xc��O��h#�!X0^f���;��Ef�n��J냼v" �XU%��6�@���?�5���K�kOY�������D&��Gzs0�L4'��5�y[0����};�e/��U��E����3��'��NgbΠe�c�l*P+�f���I�Z�*�S�sq ��dG<�����'�JSƕ}�@",i�H/��!i�U��tj����k]��sM�v�p��$Wf��_2�l�:nY�L�Ut!�I����!�`$K<1�� ����yw&?D�pn�&��|;K؞�_�a�q$���}�T�� �g��qņH��5�Ԉ�2E�%:�bH�?��G����LJv��WԞ�ūMb�G�)m�M^��@���l��~߰��^u��:����፱@���jz����T �^Q�$`̭���XS/E�[$��{�S���?�ʋ�w��|�����R��x�'���$>\]�X����KJ��&ِ���/�@0x��%�R�vm*�ݒ�Ѡ��7N���D
�󓿎�sCU�W��[C�KKw�S���B���tVT� �k�w藥u�oa���l<gR�&a-Ҝ����K��'���F��6��;��)l�S~o�?8�Y
e��U��DEDr��ς�1NRC�gv͕�&��9)4�.k�L Ur�{�`�Az�=��{)�1)����Bf�>)�I�ז��az/!�ȆLóZg��]����Sw�	�W��A�+�Ā��ĩ�SO1k�}j��:<᲼��V�4�O���W� �0dW�*�H�|�;�S-�)��:o&�h��bU���`0�[-mâ�& |}��6v~����I�*b���7�i��S��%<�A�m�Hl������3}��b�G	,.$K�.�ز� ��^95�gy���a }7U�);�7[�N����K�<�nҨ>W��B�J�^���Uh32�E��%�.n��=`����}=����ym��r�닛����=��{%��nNR���?L��6(bzc�N��73
�.�s��v����Q��]�~��P������6�	�e/YC�w	3�֌F��VB�P������*�_����ۅ6���h���E޴d�`B�M��񠨨�^�v����PV����`����*%�	���Wإ�BUW��Ɔr�.�`͐E�|�u��~�[�rh�����D�S�f�����Ә�lk�"ü5%�A�
8��ۤ�k:�j�isS�?wA��:���*�ڷ[��%HppS7�t��^�AC�#d�h�]<T�Z9�� ��S��'1#���ۺL�:������!�EL�ۍ���!Q���wA�)�N��W.��	N�qOQ��O��@��� e��狳�%K�Oo�d%\2�;+]�-V�� L��+,��¦7,	�4^/��u��A����"��<T�_�ogn[�f�is�~�>�V�!���e&�Q��40h��L5�G �ǓZ76�zI��J�a�|ď���rҲ#���]�T@�ܣ�h^7ޖza��1��\�0�g�0�}~�O�C�qt���K�x�� o��Z�vp�r}4m
t��n��)�K�s�����շ)9���;)�^�a�ug3]L�wL�#�a	�J�� ��|�
"�zo��hָ���� �uN�s*� �.^2�'r���Qq�2�gZ`� YJ5��<n[��O���y��w@e�W�
Y����J��B�v�ux��"������q(�ӻ�ڵT���Xk��E �4�,���ʜj:6K�$���f�0�~�h>�?�tbS�x��Q#T8�E�4�Ӯ���4׎� ]X��#�����J�vϕ'ܻ��(L���L���E��v�0X�i���2�ڋ�z>��ٰ��S�`�i�B�f����een��`N'C��X���7Ttɞ�?,<37`�p�y��٫���B>� OT��<w�������� S�lJ?V��]��}DI���U8�+�G�[_˦G�@*���G�q��g�,�[����Cˌ�r���kjwX�x��Vu*;aɊ
����7'����lzLS��������È>餖(ff( �0*`�~(��(US��k����� G��Z&�E2TY��#w)��^��&�5p�5K�+tm��\1.Æ��'J�)� �����!����R`�bv���S�\ 5��J���s6��}H�W���b�H�o��c�d��8!�Zh��S�����o�fhz�6l���uA?Yhܺ*�Q���io_��쵯o��$S��+�(p�	�">S�ᳯ��s4����%o
�K�-H8���j���W�a��(,iG����y	ȿ��S<f���:7׿�}��%V�#Lz꧂�y���Q�k.]P?��:E�|?7O@+�l.f ٭^8J��d�>�v����#�Qy%O�|H��wR>}�u�	� #�C'q��LA��S�#��sm.�:Xhӫ !����eQR,��r��*ː_ͻA��Qz��L�����/S�.W:(M������Ȱ��&�F���T�sc��#���q����J�������b]�ː'[X)��-����=��>j��|�&���Y�� ���R>x��`�|�E���:T0�,�.]��'�ƳIN ���r�v2?�.�	6�S���b�Px�K�k��R��<D������q���>����U��k���lL��ɾOPU�~���z�#�N	nh���"z�#�9�bŘ�ϒ`q~�-A+��W�(��aD��+���x>�'P'2`�st���ho�T����q��/{�C���V[�'��u�97%�'^���zӜ�,�Iw��׏�F���˨l�h��r*~FDB��}o�fΦ��*g1��59Ea�2K�}�.�h����SC�����+c��	���C���.��g�ͯZ1���M:�Nt8ޖ�y�qQ�vW���7Vό2�����DR��p����koP�h#wvH�AL��F�8�A�]k���w隿��L��:63�v`�s�S�Bj���*P�����e��%�ބ�a��̸�!�*�J^���&�i�͇1��:��=PS���Sv��d5'̀/��)6���||:�)?������	�~i�SUa<����v�2�_x 1�	�/�qL ZN{	�K}.K����xl�0\���2q�ea"S��ݝ�pt	-{�a:x��.�}q��覉�T����?L�t�\��%y#����
�?��=��AƲ{�8�_$2O�8o����V�U�X�,�՜(( ���ɲ5��=��
c&?���RA�x]mB�E���a�ΰ��m$k�G9���y�S >s6ؓ�6�L��U���I�я+�M�C��G��W7��f�ڰ����,c� �P?f�X &JӎO!������p^�v}���~�ğ���؎� ��L�B5�Z��0�̾g�F�"���1;����4$Y��,�3wc�ج�����^��m�շOm��A���۫�T6��=�N�����!�i��
=h�G�BФ�N�ޕ�������E�-8�������砹�K�.J.lA�Y0�,���dX�5�ˋ&�.�>��d����iX���h�9�+ 5D���s�r������i�*S�a�y[ Β����s���PR�4i���9���g�q�}����L�SZF������Ͱ	��ќR�XO���e�'�޴�,n�GdX�\�:��,^��L�G�cu�����p%�rg%���_B�g�;�
p��O�������;[��!p~<��-Iz��P'oR�ͱ�;�\�ű�H& �+-0ݟ��3�.�2��yʿ�J���9���3����Uȱ�1�	����FY=�Vj�W�����:o��/�7e������L��M��v :4����H����X�ay��-�7�c�7��DW��Y��^�'ɶpl�x�X	�EԺ9��e��Í�(�
:�}no^i�6L�����|m�;�h��_�ym���Қ҉H��/����7�UzM�pc�&h�T��W!FG� ?k�-�pՂ����<<Y#���Ѭ�zvQ�q(���."�qQ���RvdRp����O/���KiB��Ȣ hI�8+�Ƣ��A�I�}������ӧ웕:+{O7E���M�����)!d�*�����LK*�7�b1�!��^+����?\�(�)^G2�̔<rz�ݏ�n1�V�Z�P�A�����fs����vl�C0�*ňh��'v����x2�<!�ػ�/�4�>7Ș��`��:7Ή�{�9<I@��r�6h�=�@� ��à��6��5c�$-��[�o��[ ���A	�
���{9��Yޥ55�eoc�bH�1�������[�����z��H��[|�O�D���J(�� 	�Jt/#��꺇�%;c4�2e!UM�蘆|���;�S%A�:Uk��Y�|�9�4�p�	���% A��Ud�UE�'����6��N�@3��K��NQ��`�	Ľ����n�Lmf��%V��������W���T*���4�΋�䌨a�૆c�T4���5x�a�;,)2T�U�o{3�#���8��.KIE��z}}P(C���_޿Yv˱d�^��M_ �Pj�{PMfĪZ!�Ѹ��T8���d=:������,}�"��$�I������wM���♏Юx{�h�s����	��(�9ZL`�5	N�G6sJ���\@l��7�' {L�������Q���).�����r(��&N�n�)�	
��d����X��/�j�1�6�P��ܜ��L!��{#*��1጑���ވ�q4��d�|��t,c�$���?�C�<���	��9U�m,"����fk��EaT�m��t*�B������=߿�B6L�aӮ��P���_0�]=[T�:'-'���Yk�OP-�*�]Iq(�@��։�Sr	 ��E3eD��&��ժ ���B#]|��i�<��4��h|!��Ƀ��RP�Ӫ�Jì�j�/`�Z'��3p�v�ǣ�6 T���U\ܴ|i��w����V��|�4�f�C��AA�B��R-wV�N;��7�v��C�s7�z�@�:'o��1���6?{�Θ������_{p
�lC�f�C��9Wb:
���ț7�UY��61qH���jNP��ơA�F������(n��_l:�H̔8�G�YLɈ�.�y�`�SVF�/���Ɲ��$^v	�h/�S5(��r7K�[B�r��W������I��v��ا�X��<R,^U8�z��4L���f��ܽ��A��vr��X�Ė��|�R�dg_Uw���������(į��}GX����L�Q�s����-ݻSg��Q��O�r������������*�C,���8���3h,��D�'�<\���F<�	b�j�*1�$�V;�̀�L+aajh�g�Lyɴqe�g����o��p>�5<Z�H�r�������U-{i�>�Ӟj�1RN����*�����r�t��^Ic7��z��`�P���~�T��>�v�8V�_�y�V�c�~fte���%Ư8cD�1~Ŋ}���{�*-�6;�>r�4A� ��mx��	�N%����T��ٸ)1m���� u�E�N�C��z �r$���ӼP���R����/��"�Ҭ��8�W@��-�oZ��@�&�����%�2�4��]�kCY4�q�����$:v���Ou�@�����!�\8��^&̱R��Щ��{��6]k-���ę0~������8eƃ�m���k�"�~<2��m_/�v���B�!je��gQ���7��*�*p�!j���������S�ܑ�.���¶w`B��Z~K���Y�dpA���/6���d{�ٕ��	h3�s������.\��r�	^����&��&�l���e�5�CI�p��d<�]*�����b ������kv�%Ftx6��1A<�&�{�p���!U7���Nt�����2c7l��E7�C��1��Ų�6ˠ�Z6��s��ث4�Z�4�R��>YeI��x ��ZX��3U2��'�fqK�n�)�9 (l�?�~ˠ��>G�$�Q~�K�h��eB��଱�m&��L<��"�K�����Y�ujґ��[?]./��l��gq��ʓ�ʥ	���3��C�Z�9��/4ɤ���B�˞��NO�ST+�@[GM���@���e��J��ytvԍ�����+���=�b�(���[G/'�I�Qt�c�m�ճ�A��m�%��mȢ��w�f*�@?��'F\��%��
���x��F�����V�d�o�\�e��D��(�D�X�k�{k�"^�
��G���1�����ml|��s��輆�����Y+6�"�O��*ܝ�E�k��hY�hy7Zy_�D��x�"
u��͛u	hu�����wb����o��xL�T(-�f�BDeN�}jNEQ� ي̌U��1� �6�K������DG�v��Tqs�Pc��"bF|����"��X�۴i�!�*A��@�P��{jS�q5�
aOd6^R=�f��9� b����I�%���u�K'���rcZ�[�1�3��� �ާu�W����ffǰ����nx�KKC!�҅��Ѩ!��[��u�\J�sC�>b��~��)
���v��Og�N��^.v��bɊ	���/Og���v#�-�X�F��;�8����8���7�@����|5~4�ӕ$՚�6���BQ�6f� �Y ��q���Sb�9�0�e�e�J�=խ+~��dܬJ��À��1�]Z��͆�7�- ()�����5�4l4�)a#�!��ڔ眆*]B���!oE��8���)X?/��^u_����.ڎ{���x�k R���0#xĢ/�����-VV��P�m�a6's�����P$����C٭�&����)��K�"a�k�v��ƄS �;?�)�ߕꣂ\$������%W謹��朸�0'+��RS2�M�� OQBN�%����E����������fO}ᮓ=���f���Sζ���,>f���ҍ\�u����Su���\d��b��k�u��קv����6��D�j��B
��h�P�`��Hn���Q���5kv�W���sA�yol�k.���� |t�DqӤn��]n�s�����(\�r������\�� s����y�Ǘ�W�XN y ���`S�f�q�y��o�EQ�c�6�4' �c������l>|K��4r�AA������J#�5N����E,[�:��k�-� �BuE������9��+UZ�ZKG�^��2�r�}�&������W>Gx3����d�^�bo�d���1S,1�$f���G�)R%s����Q�_P�`�#o��X��o��L~���L���FTø��rNb�eZ��tQ�\�	I��oNL�8ٲ8gϟd&Ha�6���u�W�=١�"	�&3��?j鞳 *�}9��n<xL�5��	@���Ilѹ�$3X���yQo�w^C��!r�v�E�	�d&�%2o?�DC1��OP���Yyeلc'��Yd;�F0]\�� )���S��3� ��=�-�|~~�t�3'Bh^M�rsiG���Ĳ��8�f��U�osF�W�ѵ�����Q�Vi����h@�u�kP�W�|���EJ�x�N�B���֞^Q6� }�0���v s���Q	ẟ�4�D���Ǜ��?'(%`�g��I�g�/�k ��OF,�Dq�ۨ�G��i'��G��;C���9e��o�#��,0��� Ԓ��6����!fT���߷�#ϓK��l����$�I��~I�y��Kd7�Нy�H�&�qO �\�p_1(d�k�rP'��-����X (6дzG����x�rWW�N3�:�E�:����ì���ᔕm���pLYV?M)9�,�dNr�nn�1eyM:�l����Sܠ� }��%AE����ֵ���=e��I�:��D���m�j,3U�{�5�E��9�q�����t�}	p���%���e�����Gy@w㭿O#��DR!�:x�d��1�%n\�Q6�����=���ZVc�g�)���7�}���4���>{&vF�V܊��s��������3����E�,��s0��^���C���Ƨf���,Vq��������5����.�w,&�5ڢ��@�+�`�"��ja�k�2�ӏE8�:��;���֩�[��4F�NB��DZ���^2��hhU�;:���Rv1���s��E\�f��B#㛔*��x� IR$��D��������T��e�M��֒����QC(:�B�D�$��$����H>�����nK�YG�#�m��,���ɮgO�U��), N�w�h�5�U��T���I�lf:�$���{���s�Y�\iK�c1ʅ�����^��>ۆ�OҼfH$��=�8a!G�^ M鷪:��4�b�ܑ�\yC��f����qm�4-"�-8���L/�C���ё��	�N� ��e �!?fb�a*pXјb���H�(b�G�p˸���FL��h���؀���s�M�ܱ��.��֊�1R!�'{4WeinMV��x�Q-�I����2Z�5a�Jd��� �w0�d����?1���O�b��]7�%kf�}��z���W�Z�<#l�zz�5�!b� �R�sŵY���Ќ K'孶:-{�{��C�P�� x��_�=>��%]���2�����RY� Vz1��ou0~�4�rTc��N�R����U'~�1��}����,6����e���8��lu�̂@��hu����8�@$�Dc��2Ҍ/Ddp���ļ�W�%��.B`��I��,�;��0⦯4�P8����5��3ɞ��@�( o+�P�w7��P[�ܒ-#�����G')X��X-�{��{�əX����kz��0�ݝͯ�ֆ|�[MᔠK�i8��`��o��ZV�V!�%Jխ��qɆV�.nE��6� �I�DYqS�TT�i}ϖ]�M)߈C1i]�'V �І�*(�����	�����s}���2��U��n�%�6H��UR�c�>?��>�z(,��Q�F|�Ӕ'��XL0���ޅ��G�t����;�o]!����v;��5p�(���?��Ź#����*Yg^dJ���dB<=u��0�&�M��n&�k4F+�N�y���tSjT�3��?+wh�Ա	�jGSrw�o���J�g�K�j��M:�UgBO¨J #\@�*Ŵ\�X�J�\�g�����2��"z����b���)�_^��G ���+�����ѥ>�Ƚ �C���%��g".F���^�)0[��YU)F!(��"�U���M9٬m��@�}���x��?D]#{}�%�	pɾ���^X
>g;&+�~e��֝��ը�� a�SX�K�	��X��g��驛�s��g.�1�>�W�r����ė��]ˌZ���K�s,f�oF�=�=�v0T���8| �Lr�6�%pm�`k��~TY�\7"�)r���{s2�n%(r��U�����g�A5Nxh@8�woY�q=��E֌�P'�G:4q���M&����U�.�Z��4ݑ�.��D�&}�8������o4-뫒���D���WP�}����c�G�=�
I���?n��;��y�`��
,4r����T�4ۙv���ъ���5�J�i�p�<�>��JA��`��XL���%��@�woq��S��\�L:LE2v���h/���U��ʦ�e��QC�_�!����k]��` p�ϝ�*����Z������k:6"Mcҧᯆ�S�5 �����/0;��o�	ޛ��^�*�%�Q�g*�4�����b���F�����G8�/1���#I�bX��R\�f�WnL�]��v;�}�W;o�M��! �8$��@�c�/R�����a�������0���xwI�����Fq�>�!0����4��>���r?~��"�a]��:����ۑ|�-�T��.�$�#MgiU��uT�����q�<�.��[ꢋ��,z2������'p[��mu8a��"8�t��� 7��J���E�����F=Eԙ���!	����@Z>*6E�� {�c��Wy���.M	�FbQ��]����3�.����F��Rt�IVO����*A6r��0�a͹���[��^�$<�h�1�H+���o�.⫶K8b�bS9Do"&�Q��/φ�F��{{<��<�l��4��d[.����a�g��}�"��$g�h�}{ ��x�`�#C�8�Z���iP�Ne��`��a�N��QS��&n/���(��;�sX���:�l-�{�
wG�~�*�rr����j'0���+����pd��f��t����!������p01XE�%tU�kB�/�S1��;��?��՟��/^J�$:P�ј)%@o	ދ��D$~�����f ������3�(���o6n]2$�IIR~0@���^>B����4`]��T���PD�u�=�L�E���s}���8GA	��ۨ��p\J�EJ�)�,���]�/E�{`���e*@"��r�S��R�ٸ�&q�B�|�jv�����|7E[��?��6Pm��<�s��C�S`ͅ�a��a^�
#Yo܃�6���a�����m�ni�@lQ��W���W^(��J�j\W\�/E����5� ��A�_�h����=�G�2Mw�/RM�mIRD��(��lx1�s���J���}��OE��a��W����<5S�ń��n�*ZF�8O��]��J�L��_�-(d?~@�{��S�h�W�=X�g&��+�v��6�ć��6�Ҳb3�� �aٳ�'C��f�FN�Ѥ��� ���VF��{�8���nu�0�
U {��N2+"J�S���/Ĵ' mf6��Z�Yfq�?~������5E���g�?���6�s����m�Kñj�ί�50��8�Ȋ�-���M⇭IYO�cw��
=-�5���M{�UG�T�-^}��'��R�T7q��Bv{����4��2���M̤��\��V4¤��;�9��t����`��o�1o�4�y�0cX����.��,��WM�M�^	�X)ax��;Z��� ������ĺ��n�����''�"5����JC�rmu���~��X���B���/�k(-Ǎs[z�$pG+M�f�N��a'W��D�{�5R�[���R�K�M���W��{���H���D�7�fA�d����!�%�.D�+�e$P�9#<��T= ��w5�	F'��K�P�;(c,F>/)@�g��'�VZ�Ȏ��������w"�^C�,�}�6& S�]����[c�־���nJO3��~���x=�<�J��������Y�*������������a铵Xl��:�����S(v���[���]���,�E�r�@��y�M>���G��0�P^�T<3���`��(I�E�X��F���9nF̈́���h�ɚ���;-�W�� E��s�n���~Ǖ�	�`\efQ�����$�׉l;{�} �us:ؔa��c#�"T��AB"����9��rX��h�5D?k����2�v���2]n��OW���\��ǙX8x���Z[m�lr�Ʉ��VPPr;~n��]�:��^<0�ʡIA��#Y\m���[����d>���1��[p���?.@N����-���H f��i��Z��q��+"�8��Y��`X��'��11����,��짫�'78�$,�V��R�
�u��nɖs��7�IͰ�B���#���01̙��8�8<�պ�/���,Ž7B�J��=��9��3��L�Ce���-�P�ܜ��'�#H@-z��4���V�bO&<�<?,�j%����O�Ĥ�������E �1߱�&zP��E!1�Ɩ���s�g F�d�W��
�@��oVsd>H���0��,���+	�A�0�/����<���ڡ ��@��|�qe�. 	�� �n�T�{�|�r\ҧ�9֖wh�6`�#]/l+���lJ�E�>,�:^�6�m�*�xע{����2|�͸ܢ1Ɲ�@h���T�e�E@b 8F&���`|��s/aoG,�����epNm��ܽU�ZƇnE�jгZ�(�`A������S�A�\IZ;8��"t�$����eC���s�*✄y�ѱ�r���W�rTN���������P榒挓�<�c�na�O-��,HDy�[`����g��AQ�j|���/7�p9���Z��jN���z?�~�����p��(�	K�����{�
(5G�ZK
��k�|>}��m�y�����ȦX�C�
�R2]��i�8����C�T�6�ש_�,� ��gQ��C ��Fu�J�/��t���W�:��?7�e��&�7i;$�̎ns���4?W*�xE��~���])�R���7�3J�A��*E��f/$���,j�ʅGC�!�}�sY���(A�6p+�¼�"�s|�k�Ɍqv��]wȃ#��p��;���W���8���DD��W� ;��\U>Q�j�U���ʉ��5'�:�~~׆u1}��|D�7�*r��k����j���]������p���!D�t-INS��F�EN��5������7�p3/'
�+\l�'�W��M��
'�^�C%#&8���z��w�د��H�0ΰ��E]w��O"~��U������,��3)l���r�O���e����o�����E�f,�jw��_n��33X��A,>���ك;5���`��^~�`�	�����5U�lL�_�����i�`�V3i���住17J�o����o��	�)�:��{�ik���G?L<�FBP�Ygzf���m���.-�pQ��@�v$ cO�����1z ����C �}���[�w����nkO�~&�1>��`�֤�D��"� ��
S�R����8��{�ӊ�:��a�7ˌ"���V+����͊�$�̦H�پ�c1;��]ׅ,��-5�3`���F�'�J���W������R"6��.���� u�cTz^kU�[�l�?��o��o�n��eJ)Kz�|��n��s{j#;�rɜ�P'ap�$ɍ:vz"�o��� Km+�}hX�{���%�W�#{#,��$��ɺ4�)�/Je ���cW�Ј�7v���D����%n��q�,
KvI��v��M�s��+@' N��׿�1�]�V-(�A��@j|-|oܾ��󐝴�˲� ��*����ռ��9`�ϥ��1|=������GhHHJ�o������Z ����D(f~�M2�$��_"�3/Mϕѝ�l�]���3Xdp���� ,͸+A$�9o7\j�G	��A{g����?�x��"��m����V)Riu|�� ��/�ܸ
�k�0����ԅ���ª�����{̈́�L�^2ᙑ�R=�{_kk�_����h�3��d��3��ּ|1n�Ա����8���KL>� _�c#��^)��?�-��Wo�f�]kI�H�]�|�����b�b��x"L&8��([&�����c@�F�o !�Џh��0�I��d�ppb俬�cƎ�U�������<�	BC���Xe�a��W��?|��Lv2U	=�8e�k�y�C��#�,g��[���+�޴�X1�y�}���Ħ0��v-�z�d��c��Ҫw��ig�C�5>?/��{D{�9D��i����I��Á�@F'��O�m��Sr��y+����D,�eϼ0�ل�R�^�wA�,���3��ƙ��̿N�P�<�l����/�`�K6�N��W[XNL���M
�b_���/����'�{��c�O�H(L�����D�a�	8FoO���em��B��n�9�<`,seMᵹ7H�4tȬ�[����+dm@�P+as�����`B��A�E̽�Z���`?�G�0*�$�v��U�ӯ����;���W#@�Ś9��Ok��<�DT�f�`�r��+�� =H����G���F��� �0(�{7@7ב�d<x�J}� ��S!/&cbK�ը���¯O��Fe-��_a����#����l�X�r��j��SDE	�&i|�Cu�*�Sj��`#K�gi�wb�'MU�+J���2�D��R`�O?�_pxkh�i�>ЗV��s��h���J�b�������ѝ�O�q������A�(� ���'�Ԙ��
�ݬ"H�����;����qq��M�z��ѱ=���Sj���G�l�q�1�+�"�:���|Q��C�����¸�dFI��z4�hVP�O�j^��#�d�K�|O���䊒��<M�Oϔ�> ��q|z��_�v/���n���b�{J��[�ӟ��U^�1�?:�E	 |��6fP����q���:O��ָa��ՑF�ܠb���D�u�/c�:�)�l̘��g'�wlRZ��j���B�i@z|��Ft�K�A��{y��QR�r�|�����^s��b�u¨'�'��v�?nM�8��z��ծIqA���jN�!�w��,�2]P��
��9�bq��y_��<���m�Fa�T8*��s����S^���c.!�4��i�_�x%�0M�;���2%8��?m/��Ou���d.������yL�,i�����������r�(¸p5�5�E�"?�5�ksI�{�@:�0h{���Tg�YX����*��9%	!*Q^-�EDeb/{����)�M`��P�a����Ȕ�#���O��i y(a{�Ǣ���vi�DÔ���[��7Ct?�9"E�̒y�( ��jѻL g�{GXrt~���a^������s"ӢiT��6�
�?�\o%~¼����ůJ�p�T2_�RP��i�8B8"ԯ�&k&� #P�Id���^�ym����ư�"�*Vs��B�$6����u/З62�Q�
R��ɏL˛�0
��� �5�s�>����1��֋:h���S_b����{TU����:1l_H&��R�Sv�v��D���N�u�v���Ra���W/z <aj������O��C������`�J@|��ã	�˱�!ϓɵ�&9{�Ed$�O�9�wc���e#nc;�Cp�Fh/�bj���R�9��:�չX�o� �oz�9��q�@(�K�����LׇO��4.�ѭ)T��o�hc�xRզ@"o��dR�J,�f�3k^��d.AP���4$�)�R�����E
C���Nw�=��X�:��{%%�Ǭ��-�=��4{�J˶{��fɝ��cxPRTv�HQ��5��Gp��bЇ�8�D�]�.��ի�ǥ6�f���QS�:1�?XNv�T�@�
&1"�p@rW}?r%��χ����A�`�_�U�@(kp=s �~�>h��J�(m8�Κ�`��a��S�:�X�Y��@j�[i�%U�S��Ч",+��!�؁�'�L��^ސ�K�"��L8��H���_�+�%䔢�"ݲ��8KV	6�)�わ�0�����uA��]@��G��o�>�S5x��䣙C�~x���~#P�eI`�׼�� 5f5\+r��ô���+�q�� ���4��M֣V���L����E2v���o���k�y��×μ�d�X��8`9�&�»
u�܋ ʑe�|�T�?�Z|��^}���I�ܹ�����=�7=�8�,Q���/#��棓r|�g�NR���?و�����c��T=ʰ���\l�$�}�}�\u���3�bic����W��T����z�9/�٥7J��0 �:7�Sˋj����m]g4���]�Z��wS��6�w��U٥ŉb��%*�:�}R�N�r�oԌM��џX�m��=�̛	[B��#���_����gX��l���3�%9Q�Y��r�����w�XL�N���(-��Lcsw.��IH[��s��z��A�]q�'��{;ǂN����m�q�T��,��r�kw����Nǹ������D����N���$���W����M�!�L �Ɛ�:������;7,�O4��=E��g��ؿ��;�g��W�ݠ����BC�RT}ڭt��m�=ݓ:�����n�4�f��e�����pƖ�,:S�.ɫ��]eJ�{c�J���wSpE���dF�����~�K#���ʮ":z�����|����ѱe]U�Ϛ���2�d���92w���c�L��+2���p���də݊侕ͮH�i��r�f��a���K(Ͷ�C��� )Xh�r����+�aG�;piHP���"��3)?v.���G����ю(��+Q�I}:�[AW4���bw�O��$&h�W�I�8��;2G�5���8�{��$�d`&����/�'\��:A.�=vL_�ur8��g�2���o��c0���8T��A��ª
��!��b�^��d��x�1ʮJ��sB;������ךR7)�-�o��F�}�;��c=�5���#i�����̚h8ӹQ��ˇp�:�Q����ۢ�/RL��&���>��m���p1�$V��/�c'��^��G�d6[T���<v�����1<�{�Kz��n.�V�8�lT�a�}.W3������$C��aOrjac�ܿ؅�U?OX;}=9Wӻ\9�ki�)Y�Rj�6�sA�r�,��}�{���'���6 El�3rӶ�̇��bbm�֍go�с�e����\h,$�_ۗ �"u`�a����t`G�hN8֋%���l	؛������C�إ�e�ù¿ԣ�ө�:d�m�8C�e�O=O�<�[[k[t[1��fjj.�x�ttPQ�������;<T۶׺DS��3�4���t��S ���$���O�Cz�+o�Q�?
���'�	�y/I9��FC=�X�wy�s,ڦ��6�g<ó�4Jɕ�m{1�ܫ���|����
j(��:&	�������S���_إIk�'w��h'yOz2��P/���1�N��\A����E�0p	�mxtAO�a����y����A+
�n��dBO]nh���W��Q�{W[�d��J�0�yQ�("�hr���aI@XSB���3��ۡg�⽧��`�m�ToCܾ��C9�>�𦣪Ԣ)dG�y��Z�<�A���cc��I� 9�R�m�U����d�*�K9�g���rw%��|3�����.�0P��t�k���'ڪ"�h(��B�L[MJ�:�95Q�o�*둸�(���+��a�����.���V��Y7�O<�j-���3��7D"�X" h�>1����K���������;W����]=�M[����36�c����Em�����%��Q�����JܛP�{v�Kѣ�md��w���I`�&������D�+�j�0�~)G �I�
�8�d`���1M`f<��;I����"갈�+�z��b�qڑ��P2Cc��7\V���jP_uV��i1h0���Q���}�t0�{5��%ՙM���~��n��2���ûY_��M�M���Ė��cy�}��q�Si�7,a�A_�}�m�t�"V�<�2��+��A���v����-xd9/V4������b�ލ�|�Q�l�!��6����'EC>�5�u<l�y��k5)Џ�}�g ��"��b>�h�qs����{(�&c^0(��[yj�KJ����Hk` YDiP�NBc]�2G���l���c|9qFh�cB'�(��F�ۻ�}�3���`��ߔ[|��$jl��Ĵ�������8Mvv�E��x/#�k��i�fy������U2�[�@��p������"cl,/k��%���<�@2�ߠ���BK��a����0صۯЋ�m���~c���(b���<t1l��ٜ��<X�5nDD��5 7qp@���$��q�O�n��������PZf�n��YU��\�s>�`S_�Bَ�Y���#q��Ȉ��N<�����U�ok����V��x쑜.y�����J������(�����3����1 o�?"M��*$w<����1���M4G�E����x��_���y:�ٵ��Z�&���?�CE߄���L;{����ؙ��9�'>A��1{�m�L�6�Ӳ��u��#X1�.��S|`~P�ػu(�N�Nt�[q���N�ć�/�0O%8�%D-��g/�����D9�-}�>��k�Zb�GQ��8�}OK����;{�𬽘��
�$�/�xE,o���t~ �HՉ�@d��p�s�ܫtx��;��d����T�YO�[��r�}�*w봅�b�-�E'�l� φè'L��G���!,�'x�qH���6$��*v�d�q��ߵN��Y�m���{�ЛMˡpR��tQ�����VaA��#J����A���y[�VcZ�Q7N���H��A `,AE�i�5Q6����;�#R�q�G�>�Z*�i� w��dj�hu���ߌ��	�͇�?�)BXK�<�����U#�xB����(���6I�4������ӵ�@cg#�XI}L�v~��6�l�֛w�q¿#\6��?P7M��S@p+B�T�*5D��W *�Ǳ���z��p�w9����3�0ᱱ��˻��_��g�g�������@�?�yJ6�L�Iezf��s������/q�����s�geMz�t /������(c���z<�
�R�'�L˥����J�1�p=��>ݥ��
=B	�7��=�_>\��l�{���>��I�0�Vߦ�(��w���Q�{�Hx�K��d�<d�ix���
�"㫨5��4)���RȾP�@ň�&�$B�ڹy����0�p� �����k��F�-q�x�>�a����pV�Z�&@�*	p��'���]������<8��SW+�@EJ/*�T���<M��˺1,�X�܎�oa���bEs�ϛ���w�Oo��<�K6Ai����LEe�ê��r�r��}3��s�TN��%��c��������/�ߑ��~>K�o(��Ij�/W(*�#XԌ��j�q����`3�!���r?=!������=�1H�DH��xf+F~����+�Z×�k�	����\�<#>���Ɩ��t��ԣ�
��H%��xR��	�o| ��z�n����zN�?p��@!��!�b��,�MǪ�X?��G_'���<�D�v� ێ�q��&��g�����n�J9���Xp��SQ�ز�ʀg%��P�
�����|~�S$��ޜ�T��^�v���w��V��@���L�}��]�>6��>t(ã� f��,�8����I���1_`�T^Q��_;�����%���.	(�1�\6��_��\�)��bJ99�,��h���lF�D慦�������a�on�L �n�I��m�As!W��N[��fɋ�@�q^����|� д��'��G�S���y��أ�}�Weī	�T�ꄯ�^�t�����<Ãޥ��	��`��&�� �10�v��t�E�W�#w\y4/WSo;���˙|�=��	�F^8���%΁�����
�=5:g�ת�㫞W�%D\j�9q���<U���t��ڛ�Oޅ苗Zq��ux��7��o�i2QM�N9����W]�UIW�ԋ�j�ty��2�4\�dU�U��(�Z��X�I���Yh��5=�?��8�B�|�Xa
"�i�rkv7R�ı~?%���?g�I.�rx����N�w���
�����i����}N�W8�F��D�˰�0��{Z#��7-%lu���v�3b�F�#Mi���}dO`!3�#F��ߩ~ی��SU#y��q�Z�x]:�!.{cd��e����Y<oR9�ڲsw�����ӫ���+r��f9��"�Y�vx�RO������S��<��0�$Fq~�������4��z�`]M8�gEP]��T��7ŷ�`�!�ޒo���:�E�5�Ϯj�Mߐc�Bڏ�4��M�x#��r�\u#����P�[]c^N7�o�x�h�v��AM��ڶ19��s���8�}�t<�E��x�y�[�<y�5
1����넾R���s�{狈��`t,d[�o���1�M����c��'Y���Rc�C#�]���)�[�;�Z;�w.wV�a�K& 0�!����XP,knY4�kʱ3I�
c�9C�'X�(Hf-f����
��c֠�(���[�F��,�L��gP��sc��ա�N�7�BJ�n�ōbG��Xw��M*����wl�J��Z_p]"�΁�WW���h��5H��{�[���Vm�K0��졼�Β�p�!~�sy����$l[��"��2���1�n��j�d>pM%����}gj�<#�+�E���4���A��Ь�p9����E	Zy�D�����C�x�~i�~/T	"�o9N�U6%�*�H^��?�n��.1�
�m��`������(l4�|'-����^�6��}��J;��f*���F����T�|�ģ�Q���q�f�A��%�B`�I�E��Vө�[�[Ek��=�8αF�X��ҼQ1�B���J��$px�#����6M"H<��<&�{)ic
P��̼�O@le��최��H�q,]w���=L�
��sSs����aCL�D�xDSf�g~򭵙˚��tzD�E�y1J�r1�Y=����	�#�rR3���Ze����Y����+O�!:�������:Oў�c� �n1��5�D~A�H�d`����lrк���Hv��I���Wi���0B�}�s�h7�	]�쓙o1L(�����p?1�O�K��|wI�9s&���w`��F�9�٧c�ur4olҺw_/t�cT6��DR���W�����yu�n^,���Jg3S���-3֧"}�l0䵫a�:W�9���~�6���P�T�%��'1��S�'��sY��;�)k�˛�R�]��c���͠�yP��,$�ی���=�"�#iMh�����^Z��80�{�>q��������C{�ӟ���wD�6��/�Es�&R7�2�4���OS%sb͆@�!�`A�}�k�uN��g(��g������^�HpQȈ����2�	%���Sg$<en/d�r�~t9�K:�Q�pJp���S]MZ������R�*��D�g�,��h�ab,߫eih8L�I�=(����s�W)q�~��vIS�����U��VuC4���*,d60����{t%\�y��}�Z���"�aC�8#��<< �Z�\��K��qt�~���ܸ����`+���m������|���	>��>ڎδ����Z[��VZS�]$�1o*Y�U����d�����AΕ�3�)�]��)�g��'�)`}�e�����>U��[OC��!)���-<=$' �/�ci��)�%P"+�c̂�Q����ؼ��}J��-��n�\���Ǚ�k���_J5�������XY�� ���au�6Lwbn.���l�O�uha$���s+Fm�>,�n���b�^7~R�{�m�-��
 
�=絲�	:@���aeE𾱜�R0E/������
pe�z�N��i��tMW��y���9�g�ۉd���<@N�S����8ɀ&����Ea'�\�(ޅ<5nJ�xlbʍ 1�Éf�������h$@ԏk|\��wPL  IZ�\q֙$cܬ�4���&�Y4(����_��}D�( �w/?Վ�ѿr�6{�x8�)�ə��\8v����Ev����{�j���#T��GY�Ubj������j�`Gd�z�����c7��ʶ��_!��H.�%}�%>0Si�c�sP�p�V���B05�}����ɣ�m���J�H�(q i8��8�"�ǽº�;��w˖o�C��v
k]η��ηfzw�N|�լU;��W�l�.�!��bM`Y)���	��z��9P.�����{�9{�V�2�1���v�ƋfC���3�r��/�i{�u���Γ���tR@j8G7�[�oZI��֑�uZЉwD��K�}�����<@�=�ܝ"r��ݯ;����h�������c�>�ϙ:��3���b��M�Ns��דbt%��i���3�;et��	���sT7�qVs�5���D���F������s݂���8(?J���A�1��6�h�<�|f�)BM�1�`����D��:z��iS��V1��%']21�!a���Y���x�J�#�9&�c�Hh^(��]lz�\����%V�du���8X�2��D����ǭ>ܺ���=��eF�����T���1n�A#�]�T�`�%�3z�|�[����ˍ���*����+�r�E��a��׹������l���f3{C�5v�l<{�2�-Z���Ыv���嬧�F���*����\^�E�'I1�G��B����!�	 �\�'��h��~f�BQ��%r��[�d6&h�(�2�T��@2��� ��^�F������l�ޝ��Db����Ď���E���!&'�%}E��,��e��I��EШL���Z�Y�� C�����4�"�J1S�W�vBӢs��C6���j8�ے;y%�G����8M�a�q'�Q`�����;&���Ξ�L��������X��Z��<o���KF93�['T�T�fq�����s*T���&�.�_'ȼX�	f@2���O��"�s�8�սް�]7A�����k��R��l�l�y�%���0�=��;���p�A��M���둟Ѿ~��$�G��w�>�uo�>6`�Q�c��[aP�F�4�q5���|�Q�PJ: zڋ	��!�\�q�w��Aܬ��ӵ5
�T���Fy�m��A#[Q�F�d���wvˣ�*�����I4a�p^��ҙ�e�#�?j<;&�<��|1��a�%j�o��Hj�C�O�]$�
`� 2z	'��>J��?�kNf��)�4����7 ,�Ʋ#a9F�g�'� 5������g��F:�;����VqÑ;���8CZ:���[���kY�M�l-SD�[�m��vR<$�S%��3��r �����4��Yi^j#1@�0ߖ�񼌙�dh�O��h�J�/���q���z�Þm?�;�{���/��4�@�ۭRg��q��1�|0�1�}GEi�zc��S��bO����0']o�-	v۬�3
��7�/�]�[!_�҆�K�'�b0��=u�����9��fL�\b��kiE�];���bhb��M�þ�y�vୈ@�y-D*��?Ǎ�ؤ�6�F�P�b��^k/��w�R˗�v�U���.w�de�v�^�O�>�D�>�o6e+�D�km���P�y�#^6���~.���!$�P�?ʶ�(�������9��9��_2|r�8G��s/^"����k��<�/�K��a$��z�Y���R�,�b�S�9�=��-�)\��@+P��G�|�}�C��TY��s��ڦ��A=}�s��}u2 Vʩi�}-�]�D��o�s�#��� O���J-)����}��������
G�
��n�%]���~�G�º:0������p���e߼A��#	 B� 6i�B�p(-�|�妐~��>�'�ݥ��%��&��aɶ��3
����ɐQ���5�N=�����?�Np����G	]3�.s,������W�v�MP�I��!x��p�i�7���'��$��KK�f�D�vի����S��ʶ�����C��
9*���1H�H|,E��{��L	�˃!N)��E"D��zsv�	��x뇾��F��ӻsP�����H,wOU�g��t&�#L�/����3@*�W�ug�t��p*j|�6�wtY���Z�r�x�l23��.`�+��0�*ݗx�*��A������3����G�z�T;�[:'^��,^*w�����Pr�	�Ni3wsd+�إye��knfK��/��?��8��Gғ��z��L����߮�y�X!����g�g��� C�'Ǟ���C����~�9�1�����-r?�}��D�ݼ�r*B8�5�)�V�ͯ��L{:���oP�tYX��r����n������M�Z����pl0� �Y�5s���kH��R���w8�!����X��<�J��nzg��q?��t���q�pd�ڞ�r�~�u���z���q��[sע�Ĝ�tO�%��\��R;~}����KK��c	��NϺ�B���ŨO�F�X�6��ڑ<r�#)�u�)�:;��cx�6q��ɫ������Թb5�6��#qͣ8w�� �,����}5����L-������?'�?j��h�c�l" �b%n~�t��˜r���>���� ��y݋WM����]jl�ۆ.i�B�T5��h��w���sؒ4��-����[*s���Y��(�|�t�g$=/)��O�����}4�����l�"�TS�Μ"�0�#m%$��W�E��&cP�t1�&B[�*�X-H���^�'2B1���<q�r�O
#X�/t��Ь�+)�[�q������}��k�C%��5Zk���g����W�������^Zݑ�ݗJ^g��{�E���'B;����oN�|�7=�*ԋ�� 3��W}"�.��Nׄ��F�h�;�ހ>*�|<L7��]d���G���ޓs��RP<�b�Թ��|ZZS:��ޥ��JJZ	��hQ����l.	�h�P��R��4l��up��`g��α�sY�Ƅ�}SZ2��D����j��,�R�s�R?ubD���3O)�J��y5�O�#h�K'�n�7<���e�_u#M[��B'z�M��bQ�$�)vQ�q�mJ� ���Bl���\�(��8�=|�z{ķepuU�/f3�A7�;I���8OT��ى"F�V��0^�	�O<��I:�,����2�b4Lz�����o�K�!CdpO���1;	�g�vD�ÿ�XLo�����_��\�O'����Y�����
i �J�(A_۪�7���pk���}�DZ��aa%���Eޣ
t�����/G��=�����!<$�4h�"�
��M�� �TY�-�)��z��/n_����zNyv���F��M�U�q����a�����<�!��ĭ5\���9�L�K�o�Z.C"��	��L�¶�{��v� 6 [�|C�E��1H�x2	��Uf�8H�g�N��Иb*�������{th`aϭ���g6Q�q�@���٥�W�s2p>�oq⳵hǝ��WO���$�7�]����{"��3	�\+���d_#�}��q/nX� ˲�ܷ���(o{��~d������{b�M z��xIsK���_)�Cg��A&�o�Rq��@p�����M�f�!�yΘ��E���+*�Q�K��}�"^��#J�vf,��Tf�o��c��O�u�߉�~>6j`{��G�c�:����;���p�v�ƥB�Bў�7+j�.Pf�UR����c;NHR{��}�u}
:	'�{~ʜ�N���g3R�P�hpa�j	�їR}��7���S�D�%�&�)���(�ԉb˹Ȏh�d5e��o�>�J�N倭>�IU%��)lԂ>���v+���x0'v�"���!h�}��|v¯j��;Z�	1�S_�{-��7_vͻc�ߏ�]V��\ؠ��ٽ�� �Cc��LU��ud��n��)+!D{���>��L�q{�=j��Ζk��d�I���m��棾1T��L�}2�DWj������+�@������b�X�)Z!����n�]a8St��!���WVo������:;���c��i ��O��5ВS�&B
 P�,J�Y�]��'(��X.�:����~�����b�����EE���~&���S�� �T��dq�	-��0�<�zфj�'/��+�MD��ئJ���_IP�CY#�W�(��M`��1qq��R��
~�.Y�_?���DI0=K�?���N�:�\���n����L�Q�3WG"����yKC�z*�*_ܖ#��*SPz(ĉD�唳�#���e^�^_�Š)���f	(U�l.�%�Q[g?_2,�Қ��yn�{���e#�[W��=�LJ����^�k��^��<��n��^��P��~�-�7@6�M:�Z=�wL�;e�v�ϗw��.�J k�v� �QHˆ��rb0�#�ۍ��eØ��ezw�"4�0�!Z�<�؞�S^;��T�{I8�Z�[���!	4�>����\Ŧ �����A�ӟWN#l��j��@�a��OM6)���P�:����a�{��=Q��UǛ�h�_��9c���ں�m�.�8���pn�U�{D%�U���d�;�S̬Q=$���:�!l��cu��GU��|�=ꍦ����'#s���v}w	�i<4'<ˢ,�Ӄ��>�F�W�v��T8�)�]��f� ,��� $.4L���kN>�zk�]�.Rf�N������whD��I�M�V.�[�}H���D���>�z]��Ǩ�!�8��}і�"o�����X�Uo�R�ا�tcv���R^�d�U{�z_�xGS���=�|b���M�����1�"@��s<j���u��ӓ���/P�s��Dy���.��`�zz�qUd��)�� j�
����O�k�� ����B$�y{�9 ��{��h$Mt}e3�N���l��j gw[�)�X�a��!���л��l�2 eQ�a�h�U��:D+"�霝.�Fɣ�J�ʳ!m�����&҄�J�����jʽ�SV;��l�,��	��u/���'o=~<�bG��8�n����2�٤�T ��Ӗ��@�k�;�_�{��ha��Xd)�Ű�j���s�>(�v�[v�؆,i����(�J�g�,��R�G�+�}ԟ�qD��?�DY<A���_���?|�N��Y�ݫ�Y��y�Y�Cn�H�b4(����S)����H�*��M��]
X���oȇ���W���[1q���)>b��r��3�,�,�
�����|
�U�t�mG��U&��z3f �C��LAV�Ӄ�%�"{Q�B��|�T���-���;Hd�<d�,rB+K�|՞6Pa�t���QR���?o|O/���S����҅A�iM�b�Ͳ�-6|'�B����ǳP����N����h%�E_��/��#��Ia�FWF��Y�`ۘ�7��D���Qr%��#�t�Uz1� ��9O����D�B�Rf�%�f���c�Z4��K���$\Ϳ���!�\P���?�ٯ(Ս��-�����̓u5��Óeg\�!�������y�홿q	��������颵��r �8�O��0 b0Q�(ś�f�A��_�V f��IrU	e����t߫��m�H�7o�uIc�����2 �؞_+����<`�T�L��s�)�Yt�s�-w��>�ϩe~�[QtU�d���"�X(�Oj���u��m�ánI�Pm�@��{�ug����C��I!�lX�`���/4����o�F�=\���P�|��v?����j���J���LW؟�¦����:zX�DT�F���Ъ͛��(24��5�o��'�&�_��ӭ SS�efx�]F��oPa��ۏ��u(�-j\�����W��(�,p���#cLkd�"@: Y f��%�_οx)9'�>	i����XFk����8D��0֦���/_Ͽ�Tf��
B�s,����`�3�sլ���bu�J�4ڗ�q4U%��Al����~8{_�+2b��C��T�\��~�/)���}���-��FA沂��Cd��hY?�=�	���#���6�����'z?��	2���Eǅ:�afC�X�����v��N;o���G�(���r��g��煁F�g�!a2^�u�I�kD���v�l��I�=���L��k�\M�N6g@N��X� eyfO��R�a�ys��q�%E�t�_�fq��2��"VNѰ�7���,��۔I`�
���Zc�V#x�i��P	@�DM����z(҄�*�=�u~��;���΢�4ۇ-n��>���-�q�r^;I�]������%P��^��]h�y�dcr"�bh&b�Q�`�l��pn���	A��Z2�T��|�VL#O�����8�U�@��C��~�s�ڏ`�'���[�D������Xu1S!*������爱�lủ���Q�q,�mv�# ��/nEW����Υ-gC���5��*�2L�������fI�[r�/����P(LU���/%֦��b��;}1�$�ʻ��p�`�eD�_��6p�ŏ�� 
��h�UFn�Tq�O����r
��>�C�tthCE��e�qH��e��BZ����&�<���0��dA�(��*s�\��uM��!�N�p�ON���l�4(Hb���e$6��M�l&����c>	.DA�t�s��{x(-�iL���@vt4L�@��
[蠡�m�4���8�"�wV�E��(��!ja�5R'���2c���r@�������ꩫs!�'���ӓm���g?hmZ�\qOl�4���H��)������(��3�[�M7��u�p��㻇b�Բ���D�E�.�yǉ���j�n�u�����Z����Y^������M�}h�O�j	ȟ���{�a4
��64[>�;��{���NO��������7A�[�
[u����Z����s�����R}@�u�W<�3�}=�_��XCo�`yuj�Luz/{�� }�J4��8^rkC��Y��a�os��N.�Ktu��R+l�䏩T!��A��O�P���{@F��p\$�Y����ewc�	�s�@=�߾�K�=l[r�O$�� ;�O?sUk�$|Y�0���M ��a����^'��>�H�������N��H���a �����dXs��p� &�&�>�:���.9��M$�������J����-
��ҋ��\���>jM�Ql�)�8m.l*aH�;�Is�4v+	���!�"tG��/$Jc�-��L\/KHV��� �G�����L�X��bKwu��(�yD�܍��۹�ħ}Ĭ�~*.o��E{(;�Q�F!�C�E���XJt�8�tg���vX��-�7��z�\�W�~�a�"3l�	|��\�t��t���Enϙ��50/��٪���K��i
=.:�1~𶄫&^#)����9�������@�������`�7�	�9/X��} �>�4�	b'?��:�S��.yj:�Y�����ۜK3���!8��q�\�M�jj�1�B��� ��G��u���x:&���� ��f d��Wз/@M�p�y� 1O��*���^|�'�>R�r �%��>���J�fG����m��z�N2L�b ��Lug��=�����	��y�<%�^AN)��{6cV����]�0���ġ\�r!8��T�N�W�N}�7�NB0���0g�?��c=-�K�=����s&�ϳ�Ȫ2"�FC|7�t�eU�H�Y���1�p��K+l�t����K�I�I��-\�Tr?~�o��=�MM�)���K�2��n����9ײ�a�*�P�,Q�\	/-M�w�,�&���>68	����?6Hm��xr�2r��VgN;9��%̌�r���n,�O�'Зupn�X1gZ�X͸Z�KԜ�l�������m����s^5��Ǉz����5���:�$��V�ł*YPX�;w�Ys���v�M%�4�೉ejG��Kv��	y���9~0H��@9{dJ<��1�>���;
�ԊFX7j:U�|�\��k�!����o��'s7�������x"�;���E��r�)?p,z��Lx8����q�)��v��5��R(F����<�{!8�$�c<̣X�v�`ڬ���Vr�x�(��N$=íe���B���.v��c�"��8��$-��I�F��P�<��^.\Q��4�pO�~�i�!��JK*�&�˔�r
¹j�C\���=���zjL�g�y�ue�u"�>�z��4���Y�8�^�������k������P��j� �H�a�J�@E!�aO�JR0�ypbOkn"E,ۧ��G��u�Ⱌyz�k�v�(�'������r���$�k�g`��6��
c=p;�|X�~."<�62~�#�/����=���3х}l�����J���ף��Q�;0#`Uc#�Q����=�rp�H;��ƣ�]м!�qk����Qyi�����'�k��5)Qs��O);?z�h�1X�W���,J������}߱��A�-�PX���3hW�&��{Y%.W���:�K:����J��k8q�he��/��;
Y����F��mh+hO��I��!����� �B��%���������#�͝��H)����D�;~�N��$��p�h��.�nh�h(��Cu��ƌ�\�Y�ƌ�~��1Χ�7��bm��x��[���Et�k_v�ޅ�$�kQ�s@�Ǹ�u[�@�5-�T/��)�+��D=��=gj�y�F��oRL�n�"�m�*�Xw?Ҋ�[�T��bP���h���r�A~�~�r<�!~c�!��X#�:��+�³ʊX>�h0�����o?#�څ,���E1��,%��������>�;��^�����1��C�Z���5ut	�>�c�ݯ����kf�c�[���p�'��~�/9�=����%i�Z������C�u��� �tR'$�s��ɚ���p�2����9׬eA	�����Z��޲Py��]z<I][6�񘳅��;ȫ~� ��5G���#t0BNa埣���x�|� &'����`R�<^GኼX8�9{�y�҂3c�����M@S�	L&"��8��p
���2JbT��{�ia��v�)Lb�ʽ�'���	bO�-�j1��T�\�/������MtNZO��!����J�8�f� �p��ćlnR����*�q5s���w=��DG�rl�,׬�6�~��G��f��X�ϑQK �m��c5B��д��o�>�L5$<3�L��5�h2�Z[�!�z�4`E?��+�Bu|6iڱMIm��F&����iP�|�ae<u_jl�fxý߽�<d �1��e�{���-fm�d���kK�Q��o�}i����,��r%���5_F��os<�E�ף�<˻�?�1dK>Z��n������!(�8�l�1}��ѡ��<��e	6�ܧ!=f�������\���(��cH��&�4�*��l��m;�J��e���J4X���2+�u@��D�)�������H]�5d
r@�>�E�$���I�Hr$�����A��}�T���&��������U `���_3❤��7W�� ]��H�Ϗ9ѳN+�$�����G�
0XC���(���d�-^ʅi�?A]�&�����b!���_E=�1���b�S��
�ڼ�*q�%d��(�3B�.�T��M�gd~qG{�b���x��ͱ�����Ţ�m�������AG���x.�
�"]��m@���@�-i���q�Q���_D%2���H7pz~�u�$F�6�����]��xZ�g��vSLC�W��t�I^��<��!{�L���������v�ⵝ����Д*xu�{����6	K�P����\�>ج��^�o���k�O�y{��8O#�!�Q�"�؞�97��%��="��d�n�dC%������oh�P���d�$�E�U57��ך>S�rK�I���'��.���1M0Tݜ��E���q���\8~��wb҈�S��k�?���=��J�8e�]�_�.�T���␇�w�t�.8�*Lpݷ#2��)�5r)��_�G�+�ϋ`w��h=��G_�\��� �1��{�J��7.r��4�S��-��BI�wԤ{�@#�Mwk7c>�vy��48��D�,�t��e�sH��h6Jb/�VksL@����b���q
�5<If	����if�9���~P��g`$�L��m�z+x1@���{�m���ʻbbZ�J��3u[j�����C�V?��R4]8�g�7���M��ѻj��ˣ�N��Ýh�Nn�h<�rǓR�S)��Lfn:�
�+���C��)���c`I gdm\q��߮�Ÿ]����*���2���V�:�m�+����͏ń���J&�DPY�\���t�a�rF� ��"|oc�����Q��^����0���
���h��5��	�-A���$*+�Aۚh	h5V]��:�DB|M5��%A����0�_{}�ޅ��mA!^!��_m�<w��9بD��s�<+��!�H( ��lbh��5g *���j���|{����@=wJgIY��9E0�+3=�KI-�}�:_�ߵ�0Ɵ�z���}E�����B���j�[W2�����_c�aM����闛j�Ci�K=�/�R�Vq$��:��n��䛪*[P5ҧ�����nɠ%���:FS#�#���A�]�}��/�T�d��[1{��7�K�@�o*g��Y����U�f��9�S�*J��U+����#���']�+�������k��Vy�$�R�M��]E��B�-I�}��X�t�L^���
����%9K�ZN0z"�S�j!�����twAf�;uqփ���6}�=��"�))��p���/���Jt�\�gO��taӁO��dId����\�8��%�AȬ��?>��Pajc�m��V�Z�X�������4o)��跅��j��/.E�D�i�erĎ�-d�6u��#{p��@��CcpQ����	�a��r�L9�V�w�*q��L<����O^|7Fq ��a�Q:�6�S)�sK�\�k��e��17y�@�ͣ�8��3EKGHސ&��^&7�#�i���6��1dx|!6[{�:o�J�3V��8[�����_S��{х������򐚥�-A�zJI)��4���g�)�=�T�:e���
�ӁO�8����$��Ӆ'����̳[Z������$������)p�5Y�^9�}9��S����}�uz5���}���;����V鲯%�
5��ea�z�r��/�B�}_�z�ZB6�]��Wi��FH=�H���ꭜv��iI&��+b�q�����⤮l33�9�.Ak<���$Me�s�U�2Z�p�ܧ��5����x�-�榓	���ywM��Z�Y$�Ii���
3$�3�7�1����Ȟ���B�þMp��0�ؗ�tZ�G�|�%��~˿�;/����I�T�Q��-o�Ֆ�Z�|A$��c!����^�'+� S��·��ւm9�j���T�3#.��Sj��K�ل0e�&���1�M孮�pi�C�Μ�~"�F�@y���y���!��<�Q�E�d�3���d�3�J)S��F�q�v�%dgJ�!y��~�����O�
�m 8hR �m��zė���F� ̥Ư�}-��U��S���Oq�zx
G�&�W��a&����x{��1����l����
%�F�#�XǷ��dZKe��[-=Z
�����*���G�����^��:cT�*�������9��F\���p�N�N�B+#���_V�7ܿ��ǻ������X���:F���G)_� ��ȸ�3�����0�e07�j~ �Y��_i������#��Rk���>���c�(d�4�\`[�����_M���a�<��HQ��S/!��' ��f Q��!�JY�[s�w��?2Q�9,�x�K]Uod��Db���C�ܗ@1�*�[�/Uwj0K�c��A]kA���Ze�F>�?�H�%bn�TQ:s��MtfL�*���h���Փp+Ćj�����-J��^?�rU\�BW�F^/;��P���] ��ێ���b'v�ڙ������ ��eL�Pj�Tq:��@F^�B���B�r�K��I�i��ˢw�ŉ�s���`�����5|��fM��4*�yD�ޙ��i�
u��.���?!�X)�u}?# �3|5�2�@���X���]����U� H
hrO�6\,�_�{S���F�Fg��T��Lݢ�PI8cC�\������h>�:}%5����H�ℐRbb^�
�� �Q������k������b�� �õ=���b��Z�d���F�^]�YJ����J�I��w���x���9�
V��vJ�$��4��2�4�����+�J�8}�*4�n��%�6���n��6�ye�h�x6���M;Gr�'8EPz[n�N�2�����X�q�M��u�����L�bI�o"�+�N�Rk�7�3Ȝ=<3��z[`bD��C�E���l[������b��(`�����t',����7]3�4��mc��l�����Pa��^/�����詴t3#��jX�c�%�2�0z^L��L�8kFO���~u.)�ۄQQ��)�gG���F
yqyG������	�I���E�|���օ�a+r������6|@_����"��B� #ǎ��j�{7�(�>�ފ�7&'^�/��
�*įz�0MSC�	ׅ\�r���1�~o]
���T��KjJSce�8*#;��}��Mֶ��FF|x��3�r�E�N�-Δ/OHdF����o�0z���x��� ����3Wx��<��%,Z%�k�}����{����!�A � ����&��bT���R�qs]��rkQ���<�=iŷCV��Qk�0�Qo�F�o�������c�5�뚖�|�4���{�:\gb��0����}O���U%�{\�3J�(�d��%)"�ok5�`ߊ�C�e���D飊2L6n�s��Y| ���8.IOt��x���'UH�7�ǧ{?����j�w9�ά�� *��q��W'x3DZ���Lȼ�_6�))��ŵK���p�z�ƭ3,Ũ�Z:7��ce��	o�(�	1c2���CA=�iQ����"2�`��\a'Zێ���֏�i�x������0;'�� O�x\��
܍a�KhHI�cLT��e3J�I�FLDDߝxD�>�]B>+�XrRq���^��F�{��k -$(o��q��/.dO�3CP�yov�����^�Vb��j��dq%{��&?nG��|����t+x�U07#�?����	����i���])a��@��O��{Q֫�,��5��kڿ���W�"V1��/{��%���ۗ�񚋦J���b�>#�lP�%�����䏛6Bf|F���w�R�Lv�u����G��)�P�!�{RT�!����|2W�HK���}��:���>�d��B�2,�֤ڟm��h)n䏿:��Q3�段"3�up��ޜ��9�p�(�J�+4�u��(��rŘaA��Y5aέ��祤u��μ%^7]y�@��b>��\��Z�-Nø��ed�2���� 螔��a�^qM$Clc�(Q銿�1"!�ѵ�a�1lm�%ㆹ��]"]oomõ�#J��`)o��a"n|E%"Aє�>�+XQ�x^�]���H���<��22 ��r쌾��qq=_{TgC̿�I�?;�"��څ|̎ 1�Z 0���p��@Ɗ��O�h��k��.⇪�4�ui����|/!���95fE���͇?ƿ����	�vT��Lm���Z��N�!��m��4!�Ռ�a��=��Op�/���)� !�?���$�cX�¸����Eu�|�]�H��;3Hq�/�#\1�
���L��+���ƿ����冐�I0�f�]�>�3�E�f0�;��L�͸7�d�oy�(�9�|�č:~�;QgW��m�}'z�`5	ťNa�yU�����0<mۖBTX��n�R�VA[C���_H�FY��I�,JS��>G}�k�7T(�[&m�tҿ�5���}��W���a��x..W�齡!��\�Vu��!J���>;b�K���¶g�k�^\�����^2��y�ו��K������8.�\t�Ӧ2������/@f	����נ���� �jvD{�I�����q}�e��z�cv���oz��l",���v��"�v����2��8�Q����e�>��'�P��):da���FM,��W����&-a-��.=��m��u�n�(�w��]$I��W�C���s�`�%w�N����f��H�q�~s����$�ι
L��DDVۿ��ޮ�Nȑ{EX==�k�ه	���#��ҩ��}c���D)7����?ބW�b���B��9��g��87]�F�SE(!� [���{�sKe��v��%�s�z�:k%�"*�S a�F����u�	�CJ�����i��m}_�QG�o�.D�f3�cD/�=G�{�ǹg�>@E2�C;���yh����0�w 6��^���(1����%q4�D5��C�y	w3t���Rv�{�(�@��9Q,/�M�|a���d�~]{�G��|\,n$�!F�8�__���w��������3}��2�^�����6՗BL�>���qZA��p}�xȁ�|����x9������ &S4!��f�r U�b�r��O,��y
��!������aB�U���5z�h�]��{�R��A��&ͻ����W7t��S��Xz�(��V��f�
��P����m�|�U��tMyoz��d?�Q�
�"����]#�uo?`���젵!�#��i��0Ƣ=[b^� ��q�J.o�9�t�Piw)�!�C&��'�Uy�fMm4Tu3CX�6�@��S�NP�	4�����H4: }�g,��PӉIb�����x��}���.�kKD!y��Ɠ�mB/u � ��������]@�ԫ���T���7u=:�:��)e��-�oiT�?��e��ǵ��Q�p�%�~��#�#Nob�_���ػ(�[h���6Ȋ�(i7�t?M��.��+X{���RѠ�ֱV�Ov�!#X[%�CL�2����,zmT��]��.����AnL��gt��ED�Mi1��0��/;X�w��%LE������u�����[~�����w��&2�<Z�@C̩���Q���'�����DdѠ�w^�uN�O�Q��_�1��ޢM���?�8��S�|�F>�IZlZ%+ɪ%^��k����x�$��T����1�,��S��2�he��T
��,r�PSy�oZ�Cd���!U[��o/<�	�hЧb���$���Nr�8RM6U�k"�va���݋��H%A����m
�k�p�ї�~�#�&�(;k� $��p-�_�a_B�C`q���eMx�����Fa�K��=!��mG��yM9`AMݍ���FS\n�@�|��v��W��yCV�^:�$�L���c���u��%�r/����x���;�3$�)6h�Y˭�H�<6ޣe�%I��8��y7�i��Dr��2���av/ۣ"�Q��XZ�^	
u�'=�@�@ತd�=�r��1,�m"�z��]��:��]��up~�^ɐ<��-��l��o���XH�V�$\v�&e��\��v��p�w�R<.V����o�v��v��S�V\���IPL0��d�_z���#�>�}�=�e����i��h��8JZ���I�������N]�Ml��
ޒ�G`�t[���YN��X)G�݇�`* �C��6���M|�2fMB���f�F˅ �c��6��;t6
-t�\�AEεe s���z!��t� {ȼ�i���R�OS�у��9�8�{��ui]�jjd�@�	�˷E��el{q�h��ir�"����B�"[� g�W86m���<�2������rS<�G��4Lm]�?�]I��:#�����
D�\j8�*E�&�Y�`5`>���ՄfO�mי��3�I�8���5H�~dXU#H�������˒:De��mV�z��缗#�vD�8�~$�(U~��A���՝yD�X�5���P�K{0	G��C_3v��/��k�}�����;��?ܣG�_`B�>_�\��ar͜�t�ƑL�]�����G��6���@��Tzg�����%�sW$]YA��e�(CX��	f6	��",ŽqU7VJA� 3E�ta]��d?ܗ�^��/��f�,�@�/Sy.O)�!�~�5��:�,��
W�����M1�tQ;�����.b��e���^���?5�� �nN HM&AH�������Y����SH@f0J�Sj/淠���
~n���Wb��Q�$\՟�m8�t��G�<+.]�?_�۞�?��R���э�k��Y�V�7������^/��2-���A a�})�ճ��ɛBk��o�:+��F/�E.N��{�f�)n4����&�'~�c��9 �n+@ۣ�|Wx.�/E}n��I�w
[�׀�~8�(�c���8��6#I���]Y�h�@n���Xy��]kB����H�\,Dkc3�i�V��H8��Ѳn���gsׄ�*���y-P�iʹ��:���w`�ti����7I
F��:�E�6��h�C�N�^hb0���yt�������)Đ��ǝ���sx48Z#�؍9tj*��t��ƓVz#U�L�"@��/7n��7_�G!���q�2���:�`9�ƿX�ִ�$�C-����O�x�lK�%���움�r��B�{޿b.{�����_z����.�5�ф�W51+���.����h�&��\|}��\��4�q���剦�w�C�����g"h �WM��:�`)��!*���DV�$O��a����X��j�6�WG��'��K0ik�S�uj@GhE�e�ך�A����j��`�h�|a��!��V�]r)��H�Ѯ峩�/�J����QKPVΣ�����>�W;�N�--ev�0���4D{`��d��.,���`sz^��M�q�5麬��_{^~�y�+m�F��] �����&��HL��9�LXX��{�]�����2�aʥy��3�s+�A�p��=���W}�"]�~'���Լ��`>LA���.\�M��
�d�6}�F�ܒ�@��ocx�f�L_ph�֌G-�lL�~ %�#N�5�Oj�:x�����2�&��uu������<�t��*�BD�4�	!���`�׷�풱�1���q�� f�k�5�=������^`�ף��*��E�#˗
?K[r @�!s���=�}?��h��t)!�g+��!��+��M�RP�I��t���|�ӝE�ɐ����^���������I���>L��"/�q(-?���WU�X�����	�P8��%��=��~5��;b�L��.�ͭqLpI����߶#SͰ��!���0����b�ڨ&ZO&H�X@�~��a30b�r���(�O�İBǟz�Ϧ0N6�v�)�r�jM� �@;S�	mQ��ȯ=��\U�y�%��Y� n���*B�{�q9�=�Z���c�W������Bb�z�/�������p􉓩`�y��	άs�1���$�]j��/C�ҵ��4�x�k��.�@l��8�)�|���S��٘�jR�a���E�,qi� �U���cq�0��吽�n�s��#7�u�'��� ���:���~F��aF���:���������|+ՄJ��Րj�q�#�����@p����;_�8�i�' 3�aYg���t�<dyj�������'��aKޡ	Q	� �K�O�O��J��s9�P?��Jg�-���JM]��1���g��������);X۬B���Xqh�A>|ݖr��h��5���-�%֊�:��7CS��M����)��鋬��̱��#���W��� b���b��Hmՠ"CN�V�?.�B�2����A�ԣN=m��@zv��)q����. �����X����ul��V�l�ֈ;��K���ԟg��+�ż�ɨʛyk����K=8D��D�~!�A��K�o
 �@��n9?@��}�gz�Zd�I�˙�  ��>P��\��L�+�[_�n���
������)P�j���HA�t7��=���~�e��}��JH�y|	ϰD��B�N<�O�[*D��/���2]�.�Sy�ʣ�+,�H$��i�'#N)>�8�s��óХ]��P��-،��+K�7qco"�`k4��<,;r�w�Xs�L��ُ��5�l8�tb�>SS��S�;6��"P�Z��7�I�%�1�pJ����b�io6��ĦCC�E�Q��3�tR��ș����^�g�/���փ�f��D҄��	s�.pmz�ۃ��%��sN;��Y�h��T����,S2�A=Mb\�����fc��1�U"��O�ݝ7����Bb��	��Z������K+�7�1L2ߌlw�#�*�3���;z���H�F��6#�؃�<�Ew��L/4��p5U,�vb�7q �K�[ucZ�蟓��ˆ3�.���*X�-G~_f��oe�����r&k_�\'�|��� L&�J��v� �LIt0�o��LQ]�eӉ�(Թ��z5d�ߍ��A4__�>\]��'fF��%�~���a�j?\d|��'H�A��B�N��˵��s��L:(e�dG�|�e?��M�x�xp���v�	�-����Q8�]l��~nw���$�f?ϟ$	z�o��f�� ��,i�R��=5�Qj=�F���⵼%�V��z�A��3�2�N��.l�Ԇs�3��z��,�Y��N{�Di��}�J��D���l���\�u�m�r�έ@͚� ��LGU�/�Y_��
v�L��ʹ�:���pc5��s�R�_��;��=�@L��6�XaV��j���`.?ƾ�s�8�
��i�f5�h�(�c�}wol
�+L�ፀ�4v�8���4z'dE��JC�Ʊ��h���9�w~�q�S],�X�h�����	��%�����V�J�Ӷ�ԤQpq��J�&��Ԑ��xu��	�*�-'������f�t�0�I8���9(�t����i��/-��0!�z.�U��+�U��$m�1AN�=J����FB���}A����r������;L�������edq�6�4� �ZO/�T�Ѣ��B��9���@���>o�?S�6/�f@"�����I�V�pS�iՌ��:�8����?�ʬp�W��,m�0)}hc��hnX0�7c�RP�_�΍�Goj���Z�s(��b��{���NK�}�8���v�\��fKH�����e_%Z��k��.�+YOK��+1~=���k�]L= :���ty�c�W 7}s�u�M>ׁ�,R��YU	6�(��b�t����;5����������ܼ��n�5��0���gv��T���k�Z���a���:Ic2���N�os���I�S
���"8�~/ݘ���^��g�z)���ԋaj-[��Ln��]��,��6���m���M�$�@��%g
�E�>͂�9��Y�󦛲Ȫ�/��R�̜?��!e�<N��m�ob��(��o�T�ܷ�FZ��r8�i%)��zE�S�G5�A`�㜁~3L�T��� �Ɋt�幺�S"%�;0�����m��E��6��qZ�?�'<�N�}���|S�eu������O-0SB��%��QQf~�tYx~�+6��>�3 �	����Os(�p}^�8������D�a.��Tz .%�F	�n�{��l{��^��8�u4y/[���R.��od����xr���{j$5�/��wR΍�D�ۋ�>�ӣe�Ve֊�L�#����Z��ݝP�y OK�(������bCؽ����g"�̴h��F��H8�����X�UpK}��� ��䙵Jj@-�~�	N��l�3�5��'�ĕ#l��vI�9���7����һ�Շ�8�X�D�"����+��,t��D�1���Y�07��tz���)MlG&�k�λ5�A����s!�9�Yο	hR$��u�����u�R�b����1P�F��@�p�Ɗ=d������e9��&�=(��p�3�����Z�]P=6/
N�NgQ6���u���[FV�d�Vx,�B�4���������Ou�Z<#��
��{�aځl���p<:�ک;.��B#���Q/n�3�XA��VT�I~��=����dՃ7$7�9��EG�4�u��@ı�����Z���բD@�.V���,�6U$̼����R��3�OT}��u�3���D �ٯ�ɵ�Z�ͮ�R�	:RI���Ç��� ����,�(�؈w���e�3�c��-F�@�W�6����W�OG��r�bl�������~5I��H��~p���{�z�a%R3��3����X����O�Se�4�JB�c܍o�
�#�:{�
���5�H��P���nz�(8�a���}��wk=p�T��}7��4������6 M�Jʋ��:k&�f$�i�i;ʝvA�F��H
�Ҩ�ϋ��D��̑��?J �uL]����� 6� #p�E��q�<ob/�A��:j�f(�a���~�����dw�C��!`v�h���\N�x,]�c����. ��$��LEDY��Y�T6Ǣ��c��JK��%̋���pr���	�a�̍�yb��0]eU��kҐҗ}Z%�gN�j�E�Οۅ_S�����k���g%]c��L��b���q$R�W��?�9C~(.��c$�>�^=�Ո�өV���S7&���J5G�<���ɾ҆�%�bwx�e�|�<O�"����rj�� �)�e.ɢ��<�g�?��kp�A�'iQAQs���t�~Fi�D7�=��a���fԥ�Y��y]�D� P��1��VM澰$N5�ӿ)2�ݛ#����V�B��ټ����#pz��οO9'�����=�}1�1�k��?F^~��U������)�r3U�����F��K�I��6RA➼��^��������DX0.���k'�
�������r7�����}��T��0�]wP��[֩}���Nq���|�����������5������g���>3�v�"M�7ы����ʰ����������e�c���v�g2kTJj_>"����Q�z3�MY=H$4p�>l$�]�$��5���@����['b��8�u�L��Dl�TA��z�4�{?���^�w�i�w:�}��4����`�O$DK�5���7ɈgM<�� �A����E�%�N?��FEu����Z|oH\l(��[Y�6����N��rj��zH��.�I=�)Q�\������Z��%Y��{ȩ*�o�w��Gy��x�]�T0<	��3�5�D6M��k��R��6��r���&�'��>v9������@ �W�5̫�jj�U�����v����\��<�ΰU��o����m�Rq����g�u������F��N-�ɏ�uU��x���H�a��� |u�"�]�-������z���w����>Ke�	�<� f%��a$Z�E7�B!�e=��������V<��,�&~p�-�����z��惘@/,�����,fd��>4����Q�gs@ܖ��#�����������*v	���H��p��s�0�[UQ��tE����=�>��*�B�5��U�Z~xRA+~�%�(]N�9�������
�?ś�d���@���2`l9��t]e�=� s��p�j�&3E/�����LZ�i!̃�eyf�>+�;xD���w6�j�
o�5�0
W�U�A������* �7o��-����2�̻�m��lZ�3�Yç�R���&�2�6W�r��b�>I���Cݼ�BD���S��SF��2��b"��NO3�U��r���a��'�>߯��o���UJ�!��Bz2�. ���=�Ms��s6��R�S�����R�C/����a�9�/����BÒt�Y_�x���W��9[����Ηw�v��b�[��FLj�x��j����୓�&�'�mI���ȥ����0�iY�=�V�22Z��}s�U���aE �
}��<�ܵ:��% ������O����Էzn� }2�b�,+y%b��j����а����St�x��h�*a�g�JQ�H�E���g:�Z�}���b#�x���>��ܛ)��m3M�t뫈�� ���?�C�{\�8�X+[6ˀ��򞱛�n�*�"�����f��qŎ�%E�b��L�J(���.2̒��������v�Dʺ�����I$���Ii%	P��B'J��u�~�V��d՗;�owu��p�7{%��΅�tp�i]0���%��-֨����EO�m�8Yl-��5_���u�ME����\��|�����mQ%�{��e���0�A��
� �ThD]�׆!0]+�N��/�+�򲳸eB9��q��sI�Ą$�%e�+�L�|Z�Q��u�1v#(���C���+��O�"t�t��(��L5\���� Aߟ_6�c�N��V�ͫ����F"�h��q<"8aZ�w�s�g�b�X��cҏ�-��a��*��UV4��&}]؍	���h���(ڟ�����<��i��Ԗ	c~�N �]�Y���˽�����I�Iu�k�$����)���WPmLƪ��yk8� �j��4#V`��֥�	��^Tk�{AguD��$$')ޭ��\�������j�v����u'�CwjK����7>�E߭_�^��G��>���蘸�	�����= ģVF���E�"���/l']\���;�>�pYύk]w�:���]�po`�`�Y^HQ1k������x6��Ѭ�����
���T ��Q�4��� ̀�Ff�
N
Y�l����K�)���>��w�Y��<o6಼-����?�,�1S:ou5�}��v�
�J1Dy��S��t�9�I��]e*��t}����b��o9���Iܦ��x	�;�D{=�n҂d����{)Oh�{��E��Ε�A�c����MZ˶�)���6>�E��F=>���t�Zx6�J7Ŷ!J+$�Zg���R�i������N�N�,WQ����SJ�^�F�>��y�-�zrX��*�M��n�ΡP.�7�q�E��
m8��'B��Q�j<��&޺d�����T�t�TUt���j�3�O�Q�̀��N�״7rDqF���=4�*W���3(=��rT)驌}iP	��L�ݞ<#�o^�v3L��L�fN����f��0�"-�w\��Q1�O�z�S�(]#�#}���}I�ך��	���j�B>w�Rh��ۘ?~��=��r'�p�ː�t�f�B	�|��j�h�|�i��+H���B�o0�&�`orj��Kp�eֻh�C)]���]�� GA��)�=?��i��\B��b�}��ީ�vܲ�>TR��ו8C*�z�����!:
 �=]�fB�m�"��e���$���)��e����FN���N��.�bq+)����Ѐ>I����3�yM�7
��%�ʛ'J��o�8�O�b��_�������p( �"p0���45{�J����u���`X	%Ѵ�o�'�7�*�V�xOt��3��-�"�Ydv�8:3�o���M(���Rk���F��I_v������1m?o�ƅ�M(m���Ec���6@h,xj���E�@�ݍ[���3B�\�	�B����d$^!�K"<�wl~F����M��sQ�Ƕ�E��H��l)zKU8N�y����M��6��Ⱥ��w���~q�'"ȮȯτU���ս�C=4��n�Z��:��eQ��� �k�[���udM����΁'���J��_��a��1?Li �LEH���nN7�>b$L�}��M��tՋ�Q�1�"��k����-/`h6*�A�6�>(��+��O��n0�p��v^�C!����\ѾϿש
*��k�%�0IQ۸d�;�;bM���kR&��/s�y3�ߊ�ئ�-mXv���Rs뤧�f���0��L܈'��ɬ����H��99�Hl��r�W�����u��"o&$�4D������w�����D�f��D�������Q<��{�q������ɾ�)=��т�Q��sC6��v��/�& 5ܾ�L#P�8s1'��^UWg�U�_�F [�_w�<%ע.�?S<k~=�K���QV�UR�p䲦Q��r�^7ld�:!��q�m��nF����(h����9����el��"e q>������x����������Ƅ�Oc	�������;c�*��O ~rk(�s<��_�Z�q�ם�E_MB�sPYy?�{3�5�G���=#���n�z�
����l\�QƏ��-�\4k���w^��������B��0�g���sp�u�,���䒷����I � B���X���PkB�&(^�:艂��w%�RИ�	VB��%�UH�5ӱ*��[l"�ȗ�
@wda���{��hTHҢ�\�
�o��>�`�:�i�}�������u�!����@'E��MZ�!����{�=��Q����?��:��I�ҝ'-�w�@��_y���B���ӈ�Ċ�;PY�7���=�����	�a�s�P��8���B4���
���3�#������2�'�Id�0߀󿷡D�cО����Bvz`˪?l���孝��6f��|}*�lLɕ �h�����g\?^�%���$7v�DT�O����:���M 8�^,�,�(lbV����(�>.��᡾�|[3
bI5aC4��?��Ռ�F������� �R�y�7&��(�С����Լ(i'���ϲ���i�#1��V/�F�*Z�)�B�}�*�ۻr���$��)9�k}�E-aK�_���JjѿS��yn�B���ߝ�)��7j�|�K�yb7c�V`}0o>��-�o��յ65��b�w[���S{��z�:,e�+��n`i�X�@v@ⵎ%�׹k���VV85���a���̏���nP�i@Kl�;,���g�,��i�m��W��V`6���@�$���3\�1A
3(��"d�$v���bp��`�鈄EqOoẵ!L���0���hLY�o���P5�m��k��S`}(LK����@',�7��=.9�%��#�x^�='��Q�O��q4�|<i��r�uߙ��� �t��*��+�=!i^W�1ρ�<�>�Jِ����#�KN������A���A��M����Y�����b�yC
?�Hq��� R�^ )p卼.F��8d�e`E�V�q�6.���m�î�J��EU���E? #���'�M!����4cɵ;�C��%!�����5�H{��r�M�VQ�*�������'��_�����eK��@�W���.��
"��2f�<M��ʘ�6�P�����ϿV5��W�\f�U���s��s�uO�Df�>˙N?y���e
Z�C�)Ρ)!�m
�!b�vJB��W�3�l/
C�jf��6�4(�wE�B!��cF��|��j>��9����rA�'խ�y�|����w��?�O�F��К˒=�*R� 8�V2S�wd���c��v�=����
��G*Yz/���խ4�ClJ?��h�������n�t���n��l֊P
	8!��x�����Տ���;�52����*���9���ߗ��MbCi��
�&i"� ����N�f:|�r�N���c0�m8��q�"Tm�,<O����/���p�x6i>7�k�^������/{�h|��C{l󫽬�f��t��,I�_9|�+*@�ܚM�O�F
r-��Q���B^t����t���xG�e��k��Q��'��n�Y"�vM@r����,׶�W�S���Z'2�K�w���T�%u��	K���NY��|������(=��`[�1����@�Z@!9݋j�`C�8�8@�P�a����>���<�٦Ny�$�"��-%.�I���2���������v֨FrSV��K�Zy�`��<�8���Qvov�\J�ߨ�K�L-�è0i�*�<nOrT��.���Pw������&�C�9g������Z�m�;6ʢ�R����KcǼJ�I�����	�W�����f���~j�e�B�0���a-e����"-H<��yf�n�?5(�iɽ�$��O�w��e������_�9�K\(h��ϧ�,)��5Z�8��\CR$��^�EvE�V-+}�t��C �������2E�J>V�,u��{��"aePf��*A��U�<>ٽ~l���> b�j/�pJ��'0x�{���^�Ə��u�t��]�P��Z���"~i_�dQ�'���a�D�-�FX�I�n(�On3M��J�����_�����z�ʔ�Ś=kzi�%�bf�d���0��$���������/~u�X9 X��_e��~�	w_O��;��,.���MW��9���>�!$�!��
�	�C>���Ӽ����|�1��&��̬v�b�a)�#�2Ǧ�^9��6t�D�k����U�I�k�+M�Ͷ��*¦��40��m����~�C�3�ɐf��c����P��B�^�2&8����Gb���ʏ�کep	N��䶸�n����|8�>�Π��o}����~�$����|(�څ@�θ�34�!��+E�rzKS���~��3$�l�%�
����?�k�SA��Ѡ}`��9���zIQ�J����L?0�X�7���F�7B�cO��c����PK�D��p�&+_��G���k�=55�ѭ9��`]�1\6�"�[�-�KXߴ�<=Q��ή�	�����U�a4H~܃l�8���*~FV���DS5J���=�Uv�J	j��dx��%�i��p���|R�I� ���[�m��h��Ш���E�T�@�!jR����9�՗���d�q#^���~�0�q��ox��|IRÓ�½�	-<�]���I��B��5�T_��V���x�$j����~��0�3��)������Y�/=^����3�c�ʧ�$!`=��������Oޭ�`�ٱ�U�pNl���@�ZH�|K�����0��{nJM,
ە9�JnK�ۉe&�3�л�1��,��]�~)�"��>9>�X�S�Q��a=*�3�)/-G%��>w�zUR�!��A��Fz�c	�0��hB <}��AjgE�7�"g������ڽ��X ���j�f�@�JG����:����;Z"���Fn�m��˯�I��������d�{u�A���:w �ǼcT���C݄Q�"3���g�lkĵ��Ҿ^C��.+=ai�*�
~ �RI��"d�j?Y���&	�/�w_TR�V�/H9�@�����H��wgv��ba�O�kȷ��;F�L�Nˬ,�ިC�Y.�{��6��:e���{5�uFʁ�Z����~���<Z6(�i�]�I��N��k��(5����������=C�d�Y8�����I-߂ҋ[�fP�[��1�T�ؘ�b�U�'j˅�j���dI��zC��y7;��c���i6�>�k13��qC�ꖘ���{�X�"cF4�@m�4�'�I��̦�,��!vȫ���5:�kfԴ�Jm!��9D������aV詡����N5m�n���cQu+#��F
�����DS��3��W[�QP�^��o����O+<�
[D�}$���u�<N���Of�/��E=�Ĝ�wm�16�|��.'F�Bzg�Ͱ\Wo��h��1�A[��>H^%�B�F�kJ��F�.�M�Zlx�X�h��DHI�����4\�������PeA�lx�a�S��~ƙ�v���V�Q�2>'���Hq�Kt�b������,*1)�p��vy֣���W�O�,�T��K�^7����>����XB�.�Q�*�:�>�)��V�a�A�����"�Q��zaʒ��e$Cs��;QO�E��d=en����\i�2nie_���%k�7_�Y	�0=�X}�,b���W��X�΍�F{&�%�<Z��dI��e)Bᾳ�?z�n:�7�xI�����\�:B��BnL��i�����h��9��W�I
���+f�We�6F�}8�o*��,�i"�y>/9���)▫@I(������Γ�Ɍ7�h�V�6ndZ���i-�ě�S��C�``އSC��mkÆ�_ΐ
�Iֱr䈂N��U,o�E�Bm��5+�&!"�.-2_��J�0�2,�':���,T�������^���%��X��
�N�I�&hbo��gM���/�5�ɫDő�:�����A�-y��;fQ�p�H4����p�.ԑ�.�)�^�ݒw�m:N�������� ��F�4"0!oŨ��D]�pa��xw`l4��}wK�PP3�loH�	!d1�j2?8���J�.A��'@�ͪ��yy��Os�'^К�25Xq���}��u�x�2��9�i�5qVsr|��� ����ʴ�H�#ѣ��	ˍ�@����n�r�qQI:��8'%"�>��g�va�?K��㘞���;(+{ "6��;%p4m�Ѱ����\(-3;�z�C��_��Q�
e��e�&�/���#š�H����92t�fw77l7Q�D{��S:,e��o=*^(�g�_��B:�nf�m���r��$���ѿT�V/�,o�Lˣ-lu�.(k���6���B���; ����`U ��Ի�sxx@����K`�m$��A<q��|�� �=�Zӯ��	{�Y(���s�y)����J��PHe���lG�:ӨP}g�*ƺ1Q�t+/Y�T �>�"0�}	=�Ƿ�}��z���"&�������EcD:n���(��^��fӴ�D��P��B���QͰ�����z�wGf��"��v��uC�u�A�����Ĩ>8����� 9�E�����M���ߪ����$\���P[�n��P���ä���?S)���2�Lp]u0>⮃3���[b'��'B�a����}Q����S�bu�
�
����Xd��rm�sh[��3hk���ؿ4�ج�ϔ'؞dL൐��U���s�Yx������b��A'rV��bj�D���d���у�#�烃��?kn��P-1��n|�� �����,�
; �2�][bMg,�M�Y+Lm#	��#%�@i�e�X�5����vGO��z P]O��6TH�s����R�B�_���F7��>�n�Y����9jmDj6��6J�OZ�6�	'+��5?/�jޓ ]Dk0�몄�J!5\"��N9�	6sy���ELF9r�R/4�@�j�%���P��F�'�'�ƾ	�2����c�=ʩ�]p~����������+9�F�g��bnſ3�@�~��žR|Or��)��7���V�A���F/wI ;,I���W�kfV#�V �@��ȥ�#���TF�{y��YXH�������U0�����Kv8<$bM	�}-����r}�O�D)a�oeT��������if
��b,Zgw�;���B��j��wte�u�-l1C^_<��P�#$ZS������"��,u"{�#t)�uHΓ����U��x��
� ��xw��ƵG\t�4{D� O"�u%$�Y�o #����Jp�y�R��'��s�.F���eq2c���`�p.�v�Y��Y�Z���C=��"�?�aC#:c��O��F�f��0�@:,x�H{��_A���s�����$�E�<��m���Z��ѫW��"�S�n1�mxI�dH8�$;�/��Hf5m�_�;2$�;#�r	IT�M�)_!`���-�����4�UM�v�X²? 1���ZFnND�\+�xe�4".��Xe#r�a����q��«�d�%Ձ����+L�q�ͱ���n�]S��	^���^�a����-,@��*'��@{\��Qo�+�v(��/r"�@�I��b-ВE���<���9�Q��Q�k���]=jĜ�<�G�8�[��gF��u_���$/˯D
='n	n�r3�e]���B��@q o��16k���h�1Xu���5�O͒�y4k�Ws3Q+��܆F���_�j�����
���m*}8n�/V{�.�;;��NG���M�{�r F���l节l�l�©��i�7��|�ȑ���z��MF�6S4�0��	��YU���vZ|b~�)��"V:|>ﯧs�����:o
�H���(�Z��Ć���%B�~�@Z���B$R��R]��}6�<�՜U��@���!k�O���5��ꩍ� U,��5F��O�6���b}Oɶ@a?yC�"A5��F�q��V��-j%g,^�U��H1��,Y^,�.��8���d��l�n~e��>]���c|�ˡ!�ÌAjd�N{E!� 2P�o'B����27n�%% /����?i�>g,l���g�w�O^���~~�����*ݣ��D ���$[s�J��M*�O������A=El�9�GA�0Dl�Ph��U +�?�I,�г;�����qb��E�Z9db
�+�wi�ޢ�p�[;(�������l,~�qT�����#,,�{�n�,�}��d
�5?�u�΃2���Q�!����1U��N^����?��1�$���M��p-js(�����KD�8.X�)���)�����6���;��P��@����n�,��ɭ�!*�:a�d�d(���q2(���ݳ����EMM>>�`�!���l���B�a~�tJ۬1�w���(��N���y�މ�iJi���pv@���U�p�btGG����ц��[�vy̓K���{��O�m��]f�O�:SMˈE1^�p�X-�L�����M!῿��rJr��`L��c�VKj��?{&"��5��{��kgI�wD�W��ڠ������j84�ԥ���D��Y2��81� �wxT��,@]��	�R$�Ǆ�|�Er�J���ёN*՛a���[ �o�_
?���鶏�����t���ם^�h�*x�`@���\���Q̤(T3���ȳD=L{����}�	p���q�C.j�;3,:g\�Ӂi�:���f��u����M�ŔPM���X)H4��f�9Ni�D;�0�ܯ1��0��>(x7�IcS�`#�ww\}}��>k���8.�ۆ��p�ˊ�������� Y�(�A�א<OkHNc�2�$��7���8@Z�ʍ�wX��^߶MŊ.�r�ꚁj�8�'������ȧ�
r�6yr�u���cCd�
C�G�wb&m�D�\ �+Z ��m	�����$�A�٦���W3���o4�*�Tf�6U(��p�p�����8�^� K(K��B�s'â���,:u�Rߗ,T���8�Ё�t��+�
@x~N��/����v3���]�ZC+$���K��2 9o����$l���?�l���۝׭Wo��/-�rҭ/�jې�� 9<��X �;S�t_F
��@�T���D)-k&?F!#�h���K���ճd;m��¦�2�=�0E��#�yI��-Y2�����l(5����
� ��7��Q�(�7Er�r�( �l����d�h�o����Q6�������_�~��<P��U�z}�=�K
j�^B���0�_t~m��yV��-eC*y�5v���Ԩ�R��
_��R��6��ux�
}w֙��AtR�K;�8:GOb �-���Fxr�0��#̹m_C~
�LJԢ9���lʡ�@] )���ۖ�0LJ�C7����oWmh�'h�v �u�)8��pvr4fo�W���L�&��SOs��q�w�ZP�~a��zz���ǭ�#����5_�$9WX��=�n�k8����xMt{�W�0%{�`��`�o�����2'��K$������ޓ1R��O�(Ƕ�]�1��x�/������W�g�[�o��� ٍ��O�v+4�.�Ĺ��?��r��u�Ů��"���������`;Rx��J0?��uVT�Yy�М�<����in����ו5���*�uХ5��D=6��7q�}���X�(�+Ad�E�V�D�s'J�����
��)�=9{���
<�4 /E���%O��Q[���w�C���X��w��V���tB4k$3������V}LZ�s�	�Pאd|h]9�k�0S��G��RT���5�5�d�n���_a��ն�>��DL��=���i?�V�e1�ڼ�8R\�����(���6P�5��]jd���X����h���˕.�U�z@����e�V[VO�]mѭ��ArJ�fzP/��;�$v�PD����Q�3y�4J�jW;�1I�>:d�5��/��R�����q�V^3��9d���1�[�,�,��9�Ӕ��+{B{��:��H���=�+��PTF#(�g�=z�c�$V
-���>��?�T;Hn9�˦&��x`+U=0r���2�kc��_R	�SI�UoT%{�A�^�]L��j�)"���Uװ�H�7�>�@�#Ai�Z�{3�� ���.l
���~�B]	A���c:��I��2u����=/	Q�J�m��ug�'u����T`��We��5+4�m(��O[�F��u'k�uA�;9�ǋ�Dmr��C������n�~L*ل%�d��PΏG����^V�6��d����f�@��WSq��w�3Jj΋40P���+V��P�	l�Μϱ~�G�"")Ϩg&������x���Y	�B��}poi �f��R2kt����6#\'��>��,��sL��O����8�y�7�D�޾|blS	y�C��"�3vq;��Ģ�ۛ�hX�p�3n: �+�O�a6`� l�fM6�� ��у�<�o{�4�r38�V��T'�($7�A����k9�`��bKB_u� z�z!���TH+�Q�G�P�W:��3�w��2�LA��Co��*�)��L�c��e�R6[�L`��80L�w@#ɮ�����%�f,��75�&��N#)c�\aq+�a�<�d*�Ѱ;�қ<��C�tڀO�� ��e@}�G�|5��a@3�ҫ+�6��j`:�sĿ�5�����eD �4�n(g�J���B���qXI����H�!�C�������L����=���_�3~�})Y�{5b�=	�����[&X9����s?y��@8�̻�H�6��Š�����!ߐ����_�ű�n��In���IG�z�!wG����,&�����Oj�Ys�[�9�d<��p@�9���̐m�Zd�8}2��?��1Ln�w�����x��~0��C����]ot����\KP,:��Kp}/ݹ>�EK�5c.fR
��E
��H��ekЁ�j��R�4K&b�ԥ�k�ܮi&��b�5��Y��!x��H��O�f����Ų��.(n(n$;��p�J|�R�x��C����kg|-͘�u4J�����_`�_,�&�W��W9�Af��WrϷpM�4ġ��c	09�Ha��0�=+v�䵈z�4�g��9<��`�A�϶��_�-�� d>�9I�6��pɁ5y[��&��_�(�t!>���,�V[�
�C#d����i,G��'�ֶ�0u��Ь��l�]t�U�"�2��Xe�Rw��D�,���5sA��j�36�t��{^R�Mg��MB9y�/��z揄0�-GP��,S��?�*�닖X����$�����1�_��A�{E!�8.|Ծ~�����&2�Fe�M��ÈK����c�u���g0Y`�N�Ֆ}��N�Rt����X����N���J��R�al��1ۣ���]��ʂ�M�����g�K�S]0M<�������6����wQ���ư6c�Ƃ�/��b��ae*fi<�dˈ����3�<��#��y�8�b%�OB4kа�F�����Xs�LP�<D��x�45�>ސ��ݣ��c@B��Ѐ�F`���?�9S������	�_ס��`�w�}Z}˼(T��)�[�v�� *��s�1]:7�Pbm��=�����u��DB�T-rʵO�2h<�-�[�*i[�;�6�=yG�q��㬧�;��¨ͽ�mކ���0��ðO
J�#N3��\��Ƿd�4P���C��� k��~7��"�qmH-)$:eϩ��0"�%�d�-�OD*��팈��o�_���œu깾T�����u���Y�{�*���[+��n���!Օ���bcG5/e�����N*O�� S'EpL���(��]RB���;^.���0��*�M����z�<N�)��lگ<�a
��h���x�F��^7e�գ=����"a)U���&C(��3�Ӱ�{�h��eo�^i����v#t�6^F��3�M��m����q�UR?�݊K�P����m�[^�̇�����"B�	Hv��@w�-��?��ƅ�<k�*i9�v4 r����p§4v�x�B�X�*)y��O�33��)8O�K�-P�_"�#R��S.7�cQgQ�Q��Z)\���ugB5��Ǥ�m)0uI�7v���ŧ��e�`��&������Ug�`�U6ik򞌀�A%�F�?s��<�	q�l=�:�
�4��)��3��,�zw5�=	�h�ٻ���E��s Q������Jb�h�{��ugw�S��
i�H�^S���#?1`/�#�{� c୽��f!��$]�|����^j��	.�O9+�����r��/�Y��[��|o�ܕn��렾�M��F/ .�.�����Q��Z��S6"�ƣ#�c-j���,H�@���k�KZ0�>~j��Ptz�o�"4��|�	�R�ky����Ǭ��p=5Jaw�*��IL���k�Aܦ��n���A� $"ID� ��Ѩ�&�G�ѷǗ�4bs��z����F�_����;���JW��uS)��`�����s�8���Gfٞ�1�4�~��e.��ݮ��2�xC�~c�md����ir�ҭ�X>�J�LUM�Y_�7��W^��m͢Y�{L���p��`�>��o3R�Қ�/��UNI�qWL`��8!/�+4G��-9lg�Ql1V�6o�0�2l�%6�+��)�m�!6��)l�Ǘ*TP�7����}�,0ڝ:�9
�-����x����(-�#ɀ�zWXQ3��5j�`�MUk.�n�.��������9�g�=>��A��YG|�F�	��C�bm�nGQ�P2S�"u����`�-+����4yN�7��n�=(iG����qQ�*�"B��������_��v��M�f�=I�I�!d�	���B��x�9��_e$��f���RC,�{l���\���,��&�����Y�q�]��:��n9r��MM�pU��%
�$à���z�	��(V���+��E9]0�)��g�l7�s_���!�h�����ʡ������I�H������ٸ=5ظ𭨙������"/�WX ��`��&��g��Tw�sF�*��ա�+���%}�{����+t�/���z� ў�kTi#�uPP���Vy��!�}bN���t�+�kZ#�d�%�n&��]�X�Mcb�++���>�_s.(x<e=	N3z=Ho4��E.��z?�7g�Dl_K���-ΰ��G�$*~VF����Gv��]�߭_^\�)KC��եC�|:�'�81
R!���U�x�@SK��w8�/���=0��V���b�����n����V#���/%��� ZCI��k�f���e(j���TP��F5���.NZ=x>;h7�R(�@�wkJ�G��o��$�-ň\�?ig�ÔDɉ�ˡ=7�+	�k�W¬��a[i�@=���B��MSӈ��$�5�p�3����Ln�f��� �D�ar{��wn�~(�0L��0�ٙ�^6>q7�w�x��~1..�#�NUg�a>�#_�I����t�~��,26��]�NP~=�P+%��Q���ㄛ�y�?�Kzu�����FX��_6F�J/}�s�4�Ә^���8�6KX�x|���"
�G�z�)3�Al�=�^m��}�'�W�ҵ7gTG�_�7�e�܀��:B�Ϙ��y+,�����"���dl�]��m����̹��䥻F��%�5�Dy)+��8��-&���=�ry��I�{�"�os!�d�<�������榢�۱����+�Pņ��FC�q;�tٙ�x�ַ���(ݣq!w֮@��8k#:�e�d�I@F�tF��U
�&��w�M�h0&!����&��l��vX�T�����-��օ�I86��R�L�żU�=��LSC����U�Y�p��^T��Q�]�k�ݒ��T��Q�|�Ґο�95���"A�A�xT�},3o u�i��ǉH�L�����u�ė��(�6r�a���m��E���!���1�l�L ��Itһ��V*�X*ɂం?<�;�PQ� �q�Vk�q��M=�tj])�?�ZɲИ�j�c.ͫf~�j�܈,%��1&��l];]��)�S� ���M������-�ޭ� ����Y"��<H	����5V�@�Ug��j�^]j?,I�&Wm1�u�=��?�;��j9���US���Kl".r�tk��,;a����TO�E{��ݨ}ɺ��@X�����USE 'W��o�m��!�b��)2#��^�[��E�9�?g��O�~Z]����M�u��m�Q�>��#��H��=����Cp�:�fZO��~A�z�d�73��ڍ	Z8!��[v�L���m{U����j��I����jw4ȊJNk�Q�yG1 �9Y��rv�.��k����cgk�s��Έ"b�hW5�
��Mx�,����"=@87��T�e�l�P��T@��te9�2�G�*�*�ěrۮ���+�Cc}��l�B��mJE��^�"Ug5��v���w�mj+�\�P�{�X�a
��������N��dL������LF�����*������2��U5g�b�I�������md`!�`���'|��J�ՊK,�)� A�!���lE�y{��B,��e�g�W�����x1���Rl��W*��$�<�����`%�^��g��Ǡ�� ��߁F�����B����U�qk
JU
a��t����ztc��(W�mi���u	�ɹ#������]����J��f! LPA�Zq�_%��lXeX���`@�2�D�qVE_�+d����ߐ+�p���%���y8J!l=�����PN=����4k�����^���!$�:Ӝ�ʒ��{l��p��p�j�������}�wk4Ć�1��b��WD ��U��Z�����0��-��+�d��Z%�	��a/:1�N$�8Qyi+��3�~J]2k�c�ϱ�/�8��4��m/�1�W���蓉g��"�ߕ�����PR�\�xS�ֿ>ԛ� �[u{��HļH{�"�:K)�e���*DER�e�VWEΊ�rF�������8?�1��T�:���ꂦ�(�{~4B��)�1�R����Vn@�*���kz�H~_I������U�sa��������VH��*�)�
��Y	}O�~`�jǁl��W)"J)�d�%N�#���Aܷ�	5�rJ%<����j��MN�xa��j.{(şY��B��VB��Ɩ�?�O���<��9,������M@#Q���L��fCW�g�B�� q
���2�-����d<��O9iR=7�QfH����'���U����a��Oh���O7sM�'v�긨�>�rZ��'*jQ4�����k�����(�A�����&��s�^f%�(�jWs�-���8T�r�]�\ߋ�#��U�s���O	�q��f�6�H�HP�V��C�=݄H����I��-o�>ܜ�Пpy�u���嚙�_�@[�1,B�
D��T��9~zc-{C���	����;ɠ&B��)�B���$Ƒ��`q�Ѯ�7H���+����tʊ w�n�цcЏ������!�ձ��gQ �4ț��&�b�Zz����\��.qn�d���A0-��}H���)�)�����a_��f�O-���UsP�3�l:�ӗ�"��@M2@��];��h��:�1�!IL,}3�y��W{q�Zit���|�vCm�蒏sv(Kت#�]dT�e~;��TeCG���ݚ�]��!��Eyk�&n]��b{^���0� wܦ��׿A�\�/���Y��-"
BE�\@�N����lܙ��sl;���ܖl�!"����_qq)Z	��p1�v���EšJ_VA#���%"Y"�j'�/�t#~$�5f����6^�1�ue.���G��EEQ?K�j��W�����:#�K����h�SV ��L�5^-���oÚq���2�ߵ���4��r��h+�Y��9Dl�t���.�uFjx�뙵fV�wDB3����5�
�10Bs@n�b�Un��O����G����֛2qi&�O�/>Vl�@��}lA��k��|-�^�B�c�y��Q�t�6�o����4;�&e���x��e!
��K���7$z�8l�q�V*�X�Ԣ��@d�j��rVy�]տ�@�-_@j�s�T��qkӅ�S�	��~���d�ŉ��7����<տ�z�&���b:R��\n�=#y��mº��w12��T���e���_��)��oO`d�a��|j^4��y9���B	:Y{�4��h���o-�6~�)-��,�1^�E���إ��MaB5��&��+����wF�^>�>=�[@�-�(ψ�*y5� P��,R��=*_ЗѼt����z�ʌ0�	��l�F�/���KpGG�L#�������x���Hݠ6��o���,*��h�Wp�8\�����z�E�Ғ �_�f+�i�
ó�����˂ K����v� bm�
j�p+h����7,DkG4�<4 �׉�ѥp�]	�&.(p��������F�C1�#E%�L�0GP����A�z��c��r���J$ݻ�	�7����j�c�+*GL��^��xޕ@�OR�椳��Y�2Ml2��I�00::�]����p:��Y�Γ��33+�TFכ�;��.��yZ��4sށ7��b7��n�G/+!����e�
���ױE,
#��ݎ� �����Z���T&ʚ�ꓮ�1� �!'�C�`-��G5����p�[rN�-�@��C��6
j�ygt+V@��M�=�?)u�����:��"�@%9�:�|���� �^�|5Eo��
�q�h@��U$,����
>�U*����)�F�|L�<�~��,�a�!%�0���3������]�j��7f�F���}F��Z`T��'?���7n�=�7����Z�;�"ϧ���?�{�ʋy�o�̥�/O�5�u����ЭfZ�� ��J�s���͆+��U��i�,�1˜���l%�u�kC�Yd-��M/^
G�I�(��9��w.�Z�F�K�AB�h�F&��{U�����E�g��^!bq�l4�؜�A,�AH*��=tF<��e��u��d���J�����^z�Ԡ'���-sW�_{x��z�.�,�6lp�~;�Q�
�/9�66waEh1�TN�>�n5|0�h��ӏwmL)?���lcE��p��4L;�"���HB��[�j�N��6��	h)� qg��Hk���P[�R'r	}r�?�2�,y���d"�/�#��T��K<�P3�ݸ�T{;��>.�OH�0I"I9��fYstx�T�3E��5+��2p�ؙ�}�p ����_�ZF��܊�J��B���E��A�,��r1yQ7�Q��R�w]�K(���L�J�׳Q�r�F>������s
/{p�d�����p��� !�բy0��'� d�O�\�h���_�c��� �Y�M���R���i;�r���ӛՃ�+]�*߷��W'�}.^�ǼҐ1 ���>v�.x;0���D�{7���>�괁�o�����X�c<t}=�V�OKJyN�������8����pfYM�6Vچ���Q�
.���A���K���E�Ҟ�U=+R:�~i�5�ʍ�if\��B����Ke̲�.�<�E�}d�]�M��/���W��fgs���&�GEb:����?@Je���^vjP�8d�'9~���dݶ�,�@5�.���2A�+��O%m�]�Ha3���{]�=$DA]���=|��zK9M��/,�a�nI#�fBcIS��L�ū�nM�l`<���E�"�/��%"9�\w �o�zb��d��A�A�S@��I� �t
�Ae����{�$������j1Z`@���*����8�̌��˔���: #{J%�!u3��Xc��hM�Y�h�� 9�/-L���[=|�0(�;�QA;;`{�{p6n�O/yE��)����3�՚��_�w[\@t��r��֒����A~j�����8:�C�0
�� ɤ���,�0�fȩp�,\�O3� ��l\z���ps�^C��ruL�¦����u��L�d�#���Xk*\��&	� l��b��?�)���!�Ō �>��L@3�Ev~zi�q/�?pXU��5,m[���ɽZ;?�3BD`�o��*Ҿv�ª��.@Ȏ���ve�l�����$�P�8 �9y5��T��G�{��q��S�C�^L~��ǁ�-��F����3dIڡ�V�':�~2�p�C��Br�m�iϣ�!d�����w�nt~a���b�Wl��-����%uco'�����+?�����i���.�U���3����J�ү� ;�=h,G	�'���&M%�T�A�O�cI�� ��k��Ҁ�71��\c����p�ܑ[���£ՌUF@�|�_>��[��	��~cmM �	o�z���������M$���۩S�|qm���#�F?�Dv�r�^,���E�r��)嗌yȦztR��\����$�]��+b�8_��eW�-��{�x3w�5Z̖�wT�i�u�j�@T���$Q���X�巓
�eC=	��t; �jgY�B�V�&%h����!#�CHb~�eP�)���'G�W�-�Wm�(���<�<xa��2��?���E��+D�4�\�)����}�Ael�r{7���#o�����cQ}�N!�W�H|��D�e��*}q�	o3�e�� ����eU�N���b��a쟀@R��LڗK��*e,����̐��A2���o�:��Vf͛�_N6~��*�����(�Y�V̘�T��pn[�[&���iPO]���FO�]1��v>��ï|��� N���X9ƪ��I&:����S��3��ѣ2n-��ڣa�20�2[�H�+{}Kf��9��KJC�?�翵�o����I��Lj�-J�����o�����ZqyʚD��;�*��ЋR���������)K�N1r�l!�"��s�����>E���F��_�a[���XUz�˾�,��%OMS�)�_I�ʭ
�T6���Q4o/%���~�f�<_�l��dx0���b�R�0��FJ��f�/����GN��ib�qͥ���7 �6�|j��j�O�Yl�]jR��,�`c�ʮ�A����-��a�z�fK�NE��_��aЍ���W��D
��3����YW�^�-¶_q]pzf�Yqz��-�le��u�����z�j�� 3�,�3'kDKi��]����sse�r�w��N3�󫼩}��G���EU�>�I �QdN�I�!J�\�ǀ�jc.1���g�-��r1ŸY����X��L���}�S���%q�%�>y%u���JYxm��,�����ϴ�FF8��!M�&��Aї��L�;��(	�  �)��b�1��z�:(�����4��WMD�. _\��#�6fB�jce7���l0��٨"�(��5���"W��T�Ho�ٝʵ!_��Y��7��,0xk*�MZ2�y{n!O�	"����s=�����|�+/O��x,=���֛׈�O�Ŀ;X��\�#;��<�˸��[ �Bn�g��$��]f8o���l�Q�ē��%��<5!�k��@�~��o	�3�c�S�i�$�%,Kҍ�%�3�3� ��< ��`�&6գu�(��t��8�^ZƮ��f�E��B�w?s�ؓI�؆�؋7�_%0�*��cN�]`���^!�����!��齿����a�ߋ�@̔j
��3�!A6�ɮ1/�{�U��RF��$;O)b�l[���n���&���˴�$t�R�ya����i�վ �)]�f}�z�rW]�!�v��������e,�����w��x�0%�-�D5����7�4�����eѓZ�>���ݬ6�݌~O��OY�1[߀�q�\��ҧFԻ��g΍q��M�bp?O��_�`�:,�2��Ji��Y� �+�x�r�S�V���;p���Ǐ��d�-µ�1��
�ېW���pdӸ~em�T������r�ݱp�υ6����
8u�����pK40�OiZfϨ}�$�DB�h�l�4_�`�~f�]�� �y(#yJVY�DےC��7�)۹Lx#m�n�u��!+��X�mŁ����֫Y��u���HاD۾�#�|���剿B�i{K_�}E ���t�D>ߗa�fFV�cу�{�e�0�+����xJ����vV����,j�# �+�d4�Z�<TX��~b���/j���t�5�)Pr$�//���ӄ8��D��l��Q��]����G��x��<�\"i`��-leBor9�M<��~=��?<�+
qnݷ��&�H���H��ػ�Q(�)2�xAY���2*�w9Л���
E�(^���k��H�Yl�S��9����M�n�tڥ��@�#l.
��t� O-�%�����Aw���ɳ�Y	��>����*���Ѹ,�@��,��Q1��5a��r���l���WRX�w4�U��o��!w�x��Ϲ��NYV/c�C�2F��O=kWc�����a~�C�$��3z���)��ު���z=V aY��!2�*��W��f��qc�*W4�c��ٴ���7�=�L�&
 �	���yR��ə^���+���]{�/-��X�|�J,��7�F-o{X�|��$)�}F[��4����+���1��Gn��;0E��lYt��m���i9H<�Dn\l,[�繶�q -�N��.�lT�5��Z|����~�:(���֐-���^V���U!٘D9�Zu
�"܋BS���D�y�h����������V����{������]�G<�޾�r��#V6��s���mf�]�6G�(CJ��M�@`��TX���L'G�Y��R�c�5��X��+�P]f[��)��c2���%�f�Y��QGU�r��/t������T����U�GJ�Y!L��ox}n��Y�K/���������//	(e������R��Y�eL ��{��~ςو�d}�d�.ׇ��;x%d��R�~]�	L�_�3)lԢB<D�7"F� ��F�#.Y���#a��H���?ۘO�֬f�JH��x����\��`H�nMIyn�q�6���F����"S�@yN�,*�m��~X)�i�gt�H�8�\)���Q��NL�)�ƩB��p�I3��#�hK7�V��Q�����Ļ�~t�}�85|F��������-3K���NTd���;[~d��K5��f�Z��<_��.��f��a����6�P��K�ğQx�v�'��?Ȼګҡ��dOZ4���њR�,����/�m��n��L˟�G�wl�)D�xW������ܫm\h\y���L;��H��p�ˠ�����)�ЦI0�,N^UH.� ks%�������Ͼ��3u'�"SX�K�j:��e�& H��+�-V�p83�#��6"�9���`Ұ���A�aT��ٳ��:���z�˅G�������4�'�L)y-����#:&��,
��=��N4^_	,��%�ۇC�ݢ�ϒ�*��$:D�f���%A"�$K/Ā]�p�A�ƃ��k����N:x�c\�ƕ�(�����I��^�dr��j�o�#�l�����>�_����1I�My|uNE�O�XXu'mÖؼ���8	nÐ��L-�'�_�&|�,/[�\�^Y��*��l?/`2���������Q$gM(�bzr��F ��xP'}���WħB#l�p�Bi&S�l
Y�0./vb��e��	�I���%�$!(����@:	���C�W��F�`�M�����pA�2C��S��ė����HȺ.)8��흖O,K�?�g��E%3]�3�3�� w �n�d��qF�gE�}^�`�?�"p9,%��e��'�� ���W���>P
G?��3��_{��٫��?z�)/��	}#`��YX'��溽��\�dog#xN����>Ł�H�f_�e���dt�0Fm+����	�!m�HcS�r9u)։���̺�.����V�_;�G�� �΍"���8��,8q�ۢ��]��ZpO2rD�@p0�}�Y<H�����N�n�Ԑ�
<�h6��/r��9�c(J	��E�їF�.)Gsu�^���Ϭ���|��T��qao���&PGtOȩQMb����tQy~ɠch�����ܦ���ڏ3=y[c�E�F_�21��2<)PNu��j���j<0��w��ü��wғu��U�'g��3�������g�d�1��d${@괠X�ݝ�H�4�x�>��&/a���g����h�Ф���Y_=�~�Q�l���ǧŨFQ�J�}��^�]p��t�)��|Қ�-�%�7e�y�2|&D��>J����r�Di5)�~��6�>ݲ�+\� p]��AS���Ne�'��H��ѣ�G�ą��@����Sg�T@��i�K�CG'�T jᎤ�rj9�Ѿ{ay��p��O�:�8�/����Mg�g4�0å��<�)%h���e���1��7��S���G�:.�)T��3�IqO�? .��M8.6�L��s4��� �Yr�7JQ|� J��)�8�g?9M���;^�O���b
EǬ���_�Jd)g�Cg~ֽi��ޮ���KV��H3�Q�ȥ�O��6OM+[j�� �'
�{ʺ�Rߓ�;qr%\/1����\^��;^���>�# L�G�nϻ$������r�\J3 h[K��j������]M	a}��5�=}����P�}�%)��;��A��fqӠ�!E�,2�+��mpo�H%��Y�l���y���,��`���6�Ǖ��f��}P�U$���,��A�B���`^	c_ŜA�K޻�:�¦�y�R^�Vk6�7Z�X��W��g�?��{N	��(;j����|��C9"BĈ���SH�L!Pi�'h�a���]�i'��&�wz�[�$L��F�>0F0LMH_�rzR�/l�u;�'j��$�����N�\ӈ��N@?�[���_��Z�tYEꉳ����_}��?\%h��6���%`�����-5VW�Ֆ�mĲ��S��lye:�>q<>m�3o5&�������[�AΆvſ�����G=Y� �ԆZ�`j>��*�s�94���j~]k���9��/�Αũ��Gn
V��
�� ���$���Ep�"AVdFԴ�K�d��׉��
��J��+t�s��$�˛��I*~<�.V�t�SDT��g���u�&\Dc,�*�]=���K��!���H���A��0��[NM'w�D�E��Ǽ��P����E%�/Ů�������uYc��O%���������^r u=;��\�[���ȟ+%���
�i-N�W�� �ז���dzр��@��_1\��xqը��U7I�;3��z��
�x�;�>R7���i�g៩΅
�x��4���RY�+W��I%	UyU_gA8��+��BcPgn�t��`{�B.U����gUJ����u���H<1RJ�,0�7ZJ9��@�m@G]�/nT�F%d�ӗ\:�%��?�J��Ԇ˶J�O��h�	�Rʖh���]�A@\-f�2�&Q7�3�;��}U=m�K��f�T[��FXY�������qZ�Y)��=;����p!7 _�qF!k�d��@c�5�U3��+8����@��d��K��9�n�
�.�����e����4�+��yB"�}�5�
���3�6��ǘ*p���4m�׾�t�lW*.��ZlV ���EJ۾OB�.."�a��ְ�O^)b��]�����p�ݝ�<�YsՊ9;D�5]��Gj ���" w�v/�>$ 4ŝ��,8hj!��������f�C���'��R�T�f��Aa�Lx��S�u�P+�Xe�ۢհ��QH��A�ĥ��T�� # F��3g�����,6v~� ~�rA <�IN��c���{R�.����է鼴�y7ˁ~0�|�+�R�-q�+�}E�f<�����o�c�ӭ�������p�0��H $��]h�L�AF���w�_U�D؏1ծ��?Y+�A�i�`�D��)o�rTmv�Xl����f�%.!��3fF=K�|�De��q��Ni�ЙY�>ܗ���ڜLPn0u��y��N�0����	u,C�Bi���:�u
�p-��]��G0��U�G�
��:����z��g���R!i�\[���T�7^�j-�R�=��:[H+�'{۟Q�ֹ}��p�TP+�.� B ���A��>@�).�>�P���^�)��+�͜2�51�����Y0�G������(Ui�����P)"D��Ni����F�g��c�^��LnV$w����9��2�盇��58Nz���y�o����|���-O������Ԙ��*�Y�/��c���L���̳��d���AD����(t,��(A��O%T%G'O��ً%Y�B��1���V��,��`������C��J� �����t�Q[��k��ݥ�~a���K~0�xa���=:�NĜV�����֨�cW'��]:�?�bN^�� G�ך� ��|�����YOh�J�6ij��0Wx �H�9ʖ�a�0N�����>_C����p�Q���d�Eװ�z;Db�<�<I)#ĸ�IC͛<k�ؿ�r�;*(y��H��![�B3�e��2��)���>����(��C�#P~xAP�IJ	�pyh�������-���܋�*�ݜ�bS��)���>O���$���s�R�j�F��y�����Ò4~�N�Wr�h�4�e^�5 y���X��5v�Xr��06���u;��6��6M�v�B�s�M�']�B�3-�}�]��p���P\J�w��[���M�[!�����Ϝ����������q$ �6��SLW�C��z�S>K;~e�"��?�"���:�D�xn���j@�J�2��*b(\���=��w���+2f?�Lp�ĉ*%���D�� qG�١r����|�h���kP�7FI*� ��0l�-^'̽pj�&���`�S�њ�	G����>(��#�D�ĥ:a �
��y?< H�C��xN^$�k��;)��t�\����˘���om��k-2K�%�͈�W({ ��g��\��י�+1,�S��B�SA�qՐ!ɐ/���.�ц��S	�rBWs{�mr3t�c�(xQ4�}HC�酩fYOU��3 �:x�w������a	�#�Tn�%���*�.�+.���W{� �Yh���E<�������T�@�5/!T�.�!^�\E�J�-�b��m�w������ HPB/�嬖��f��@�oc��Lz���)���}`��A4�$� ���]���|Ȑ���}("1^{���Byc�hl�bo:��'��W�R	|��8�%�i�,�ۻ��؟��>�K6�Q�����
!TT!���Ny# 
�F���"<46���¥0�Y�?jnOi}t�[�O=�Pv��@Q�#x�X�! ����v�f��d�ڑj�|����D��M��R�A�U��Xo [f�]���/������;�(98}6�3TP��`,d��1�а��n���b&s���~�5����Ϟ���Č����E���\��C���W�B��- ��+>��0E�)�up�k>�u�95i��ѣ��fe�u`ዚ��>x�l d|��!��t�SM�ʻ�~
+H��&���P�ٔR��#a$J?�k�'�k!G<�&�W�����̄c����{��fE��N�c�[5�&u�	3ơeۜf��&�����KwWE0De�e�M��vۛ���~�C�U���j3�C`���9۳���8�mpps�D~���^<������/�fe8��͗�e����oʞ@[0�8uX�1�D���J��:�z�����Fk%'4:ΐ��P��@ȖL��YX�d��?��	�I�WEQ�C�t����,�9�v��fZt](͡�=5&t�����Y8�(X�\��8w.Q����X	�~\fBB"�[��7�� �k�tQtZ�W�&����������-[S����0��"l���G��PNn]I�d
l�q�`2�5���SЋG�����]�~��]��x�i1(d�Ҳ;Q��?�s�wu��q��8���
[fж�-�n�V*��~e�ٔ����?���4��)���2��HP��1��ųȳ'�
�,���D[�;΂����û�-��:���RVUJ&&�� A(����ԇ3�����D�Y�4*��j���|�D���#�-����9�_��>y��@0j�����x��8�P��)A�f�.�U���t,��@X]!M���I�#e�NAe g
� ���4���L
[�j��; �X�,/5�[S�o�i���?��h�������iT(�b�}�X}��������ui�-oc��~i �-���^����z���_�}���[I������ժÃ�jN]��JXAb�fў�^�P��0�^[��I����n?D|��>m_j(O#�K�Gw�۲�=�ݹ��B Hg�c�<����|YG�1�Z�I.��3��QƀY��>�b�Z�i��(�P�#Uc!�a,�ΒCgư L�M�P�(ѩOL\"�#y~2�U�yۑ�Y��R���i�v���z�o��Vg�����8Ǽ07�q��?����\�к"H+��{��j��ӜU<��`ӿuB@P����6W��dQ�b{��	͌H�߳��J�U,��(K�s=GaT�h`�B���^��&���k�z�C��E�jI��MǱ7�'r�OeZ��T�m�2��juq��?��]v���W)~
� ��5�@lU�Aer�4#��@,�gU� �Kx i�j��'���g0�_eC��Xm)x]�`�Ÿ����d�m�s��� �\������E eR�s�Vu�|����;����ĂGO��^/�z��^����z����7��˿�	bV�q�I���0Ӛ�C'O�}|�Zĝ�_p%vt���| y�f2o:NjO��{,X넏*R�5���B�
y_D�P�RU'��-O�M��l�[����V�o��3�V���h�6-�kW=�0=��5��]Q,�M/�;�঍��/��^,��Rg?xƛ�s���ɉ$�| |�{�R� �=c-��z6���!��m�Z7�]ޔ��v-A�B��sS!�3:O�ͅ�j�N��Ye=[�W�
�m!��"�^F�l�M"{R`�^���=fi���'�Ze}�o�Ϟ(�U�':��t��T'M�Bn��i}��<$�m�_H����ms�6��fmtM&�|�я��睿ig��LX��z�>���<�>�?x��hB��gnz����~��_9�07\��4$�״�|)SI�)'��=-k<4X6:�E��JGy^�-z�
$,�����'/d�ū�P���=�Km���P�ӷ'Q��fGh�Խ]��S�'�v���&-hu�>B9@B�h �D T9�юY��_�˸ä�3�
�k���O��F�b�`���W��>�RG�?��_ί$v N;"18V�+�&
��y�C�׭'c��Y�r�'R%i��ρ[Ea�OO-6��f������!웘�S;@�w�?*�������W �J�#[C��ǆ:������/`�@�0�=�p���d�?�KiӒ˒��]�-��^9!��~WXY}
�w�}�]�|�%���=�2F�В�K�e�W�Mn[�7Y���1o8�9`��$7��"���M�&|��zh�jyLb�K"�9��L8%y���ꛛ������W�D�;�R��{*!�x�B=x�J"���9S���"�>S����I�ܥx�uM�!���=��,m�l{F�o9�sV,�}>�$jI���D\��gC�A/����b�@a+sx�*N�ܻ��~Ǫ��zN�|+/f������� }J�:�5S�LD���l�X��E
��vdg&?��5�����lHuHw6��輿0�"�}ҡ�X�Q󥃃Cǻ,"�1F͂J�4�qz��3p���P�ǔ������6�u9�g(DN2�<%�����9���jB���'|�`0�c&�t�4��w�?f��� ���I�F�on4��E��ʫ��tl�j�>��ۍȀ�@������%JS��ԍ���E����(x�&�VoB�Vt3��re%��m�d'G%
�d�s6ߌe;��d�����z��+ap2��l�����h�!�/�:Pi��^1w8�'��5}�I��!p�_S�G��;;mR�;��h�ۗ��U(g��ĻW��)Y�1��;Kp�	�m����0W�X`b�Z<}춦���Q1LC�v�������h��&�ILpe ��������{IA���Izձ_�OU�xc�ɡs<=`\;] ���� D��?�_��o�7"	@�%�b�P�=���#�;�"�c����^�	[~T��b�D�J6����A��|`�<s|��sjR��%"���wp!���Mh�j� |k�eE���>�tڧ?i�j<�LjL�a ����԰�S �'�D��5�n������%�^�e�42T��( Ъ��x�֧d?C�&�ļ��`2W�oX�~S�v2 '�?�Cx�fKCV�i���=�-�]E��#�`^��)�eTKY�p��Ζ�O����B��c���Le�l�G�V�)��H4��7>"�_�ō��sʆO�@��j���䠅��y�5�-�ԉӻ�UN�VK�)V��e*t^%��5 ܡ�j�	���3"�*�ѷ\s�rb����?�X�"W-�m}�TY��)�䟚O����#�H�F��ڷ{؅�WD�d޲"E�~v��$ʕꞿ>�<�0���>^Osg����|����{&W��5�obA;�F�㥌N�!�兜<X�mDWzÁI{�$�|��=��$$/��w)F�_H����)=D��C$h��C��}��6�v������v�����Ȧ�s_{���|������)��|�"D�W��NP@���|��lx5�������U���o�٬���@`趨 �-wY�e�7����YD����J�E]�[��J6<��[�x��5n>V���FSP ���uʵ
:����� 'o2��ʜg6��}G[�-"y5m@�F�5�V���k:�{&L��-"Ǭ1�O�6����͔���!��L(��f���'>����z��=��SZz�*rQ�b���Ŝ����W܃>��	������knpj�V�k�� �ۚ;���b�����r� L*a�qEn���(=YN�-��r�n:�C���p}�C Z �)S�%�A��B�EU����	Y��A�E�y��cMȏ�?2���.| ��0P�y�mMe0\[>�� W�����?p�[@1�J�kȬ���7������@�jS�S�zuKV��=�9˩�H&�M^_��-��H�ǭ�Ǧ�~���H��GTu�vٳ[)R��ce�,$4#�W��/��|�+{t�%�@6Ө��NC<�s���
g'a���JN|߻��ax���p���޼Y�v*���j�nG��M됴�[ٵ�Fǲ��C`Nt���§��s��p������2q��XVGL��4?�/�����a��pD ��靰��e�L1/��J��e?���e�HR3���O���ǚٯ�l~��p炮�{���Bѱv�A�9.���<A�$�p1�Ƅڢ��ܛ��u9��R�A�"e-�m_5S���
��g:����Wt�v�懻T����+U�m��`=o�E��ǹ�a�<}�.Ic�GS`f �/��C�p���2�����`)�BN���U�YR?*9}�7ǋP�<�9]{���Tn�Or���[���Q�W�v��LH9�Ci4!��Lm���{2e�%���JfqoQ�l��"��H��fn�L"��f h�I����uG
�>3��tF9'}������y3*|Ao[�,',�)D�_V�P�-�1)�7��b�r�_"1��j����|~GaѠ�����%�\�BFw���e�'�#�\w��m-T��Rr��� �I����/)�EݬC��c�r^k>�Y�Lv9��n�"��!�1N"��,�_8�*�rO���y�l�ﻩeo:�������D�R�~DV�$z�G�pH��#��Af[(�>�a�;�+�g*�o2�$��2w�R�;ޱ�b�Z�g��.q�2�f�G�k�>B���V(��5�w\&aJ���ˁ���9�Қ��+���S�=���g<򉛪�F�:h^o��C�L_��X��"S"�2�K�TQX{�t"d�ՃGbGi2zj4|������@��QGQS��V0ZL��Hˏ��>���. `\��ݶ�����������`�-E���&�s� # H��naN����m�߲g�u��+�]��u*�"k�Ye&� �;pO���=Lc���_$�%�iz���0���>�p���1x� s���P0�t��n�B#�6����P���F4G�=��Cy6��Чpf�[�"��`��*�KG17;hI�Ó���k&Bل�t|�S5�����n���CR��l�.�?ٛ�X.=��e��	�1>��ϡ���H ,9z?4�rK�ȝ��JJ��6ȏ�m�#�L�=��4��[pߖͤ�EIn@��f�@�Yj���հ
��	����(��\�֡\��;��P«�R�����o�Q�p!�f�:E�i�a�|QLi�p�.E��k�[?Qp�6���"o5���%��L��汱K xY@>�Q��@��׋_x�<�d�r�ɋk{�e���x��� B+5tr�җ�ɿ�Y.��|��L���{����	Яv,���$�޼�M����F�a��S���@� �S��Z¯���E];k;W<m��߯&�����S��:]�ò:0�ETx���ǐ勧~Mө=�2+"#��f��ƽ:�8�C��� eQ�MɚN��W�Z� ~D�䜑�H�����g6�m�yTU}KksKY��0ĠYc{��z,���w�2��pRQ�#�1�Sa�ɀKRg m ͮO�]�tPOd7�r�@�*X�4Y��S��d"��]�hT=�q��te�c���KS:^��e���������g:���w�~��>ܳ՗��d�~;e��&���� lTPo)�]��C��1R�jfʹ�sM��Y�C�a��9Ab�[V`3��ڒ�Ȏ*D��<��Te�Z`��l�L�vT��;�@l��N��M� ��>��S�������E���Ӄ�5:��vg̣�7PNE�@�xU��F�n�b��O^��Dӏ� �v�.�[�5�߳Z$eAI:��!����`#;�S�����:�l��
BMp��M�p�-�`Ф��<Y������V]���ő\N +u�CqW}ZƤ���]<�P�g��mW�N��&�l��q
X{����<:�)Il���*����<b���$���U���gTյ�2�J�1M��i���(������G�l�{�yeXr��ӕ�y�������^2R芕�;�ϋ��AEh��>c�����F�!|P��Z���+R��+�/��79(piT�\5�&�ô'
��-.O��`\�I��K��A�:-�	�6��͏��=Q1�5�$����f�%2���C~�Q�ڪ�k�8�"K�k�M�HK<�,v�	v�"U=����,�y���L	>�6�;��C��r����cQͪ�H~t�%��h�!�<�X+$�-�f�BK�@��ؙ��s{��I�1���:�0e%���iRͯ>�e�Aw�_�&�,�jf��a�� ^��`즺��|���J� � �<3�3�]�7�j>�)�&�� ���`�r)�ΐ�dKJ�_N����U�s7�aL�xQ�)�Q�Iȼ8��RG�9�KU�,<��t|�~�I�|ujN1���98���g)�"?P�t�1}��g-�����t�on�^n8�\��Vy�s���o�&��/�\�pU}e�=�+3PH�'�j�,T6Ê�=(�fM�pi�-�F~�pB��:��0�.�_�hȁ�RQ��(�.����1{G�����FIaط^�;P�L�7U�G�\�V�	�����5�s+tMB��bvۼ���m�n�,7}�pp�v����Qq��5��Z������V_���@�V�vVDK�ԛ�/��qK��J+E�f>�h�n��������1����6�LS�����i�槖��:�,G u��e�Jm�ͻ'���ҊO5��p1ܪ�R+�@���H���S���}>��;�qG�OD�Q�^\!o�UN�{�"��ì3�r	���B�#0,�2� �q���f��a�roM��&��Ѷ8���e3�k}��/� �DZIh�b���.L=�O�'*<0�[^���~��O��DE?�-9=�e?�&���ηF�^������d��[C�2�5���ҋt��9��nP���3����Bdڮ��x�$U��	��+d��/ �t*c�D�GY{��@��E�X'2����yF��Ð���/�ȷ��h���l�a�Э��-�U�|��S���c��X�DQM�fv6Bf"џ)���)��z@��x:^R�0!6���\E���*��u��h|'�F:<���H���N/hh#+󜔲����.tM~q��Z:gN�၆�^�-i�N���a?]F�J����[��v�Oo��Q5s>��zf:�����cz���N��9y�m��7Ò���e��fB��s���Z^��]�l�C�^��~C�,�mx��D����i��n���*���}+������$���9�B���NW>O���_]8��0�^��TK�a����yiCh�_^MI��X����
�A�2��)r�N���7F�t5K
l�;3�Ւ�T��g����]��k߀�����͔�тT�qvL.C�7Ą=v0ێ,G�O0ቋ�C���9�X���F%.��������0aU���l�G�TI�;����\�{�c6�c=2�Q&<���\ʕw�l��c~����s@^y�ᨒ^����9ղ+��X9xZ�:$ޛ���� xɨ�%Q$q�m�����T9yyŃhj�s�!looX�@QS����C'��h��@D���+���� �����S����v%l�Ɨ�&��x>Eam]po���g�Y޾u���E�f�}TZsP?n�s���1@he=C|�^5��}CH�qv+�F�4g��b�d���h�� F������µ���&��Y���RCo�uZs
:����]<��j<���&H· !"z���p�81��rw�N��#�^����<-���[&[8�~d?+%�W0�3s}/��(
8�O�^�7$ �͓��':�SE�5�xQ<�qn����ZguJpS����'�p�;}�(q���^��	j ����
�yQ䠐����j |�P0kI��aP39�� �B-M8sh���%.�a�D�v6��+[et\� ��5��*]Gk�up�פ����9jh��H�m�f7���.'�����eM sÙKr);��5Aŗ4LBl�]r�h9F{t�v5^��YN� cƇ�KҎ���6[7c��۳'�H�~���O_���4.��qh$?��1 T�@J�ip9K�.���D}�і��h�;���u�z;�l)�m����#Y{.���䔇�u����O}os�0���P���r2x?k�zk�4������z������F��-I��B/��`ݖde��	Q�cp�7zU�C�)��QgT���8�\[/~#�o���wI��H��Ō�F@� 1���	�a��z���)ɘfh������0S�-�E�5�P��yE��x���#�n��f�_�/�VZ��Z�*�;���H�s���{U:7�i��&��z��W
 y�[.i�5;�+�S�-��؎��{%TE�т�(��4n4��_�x=�� A&�K`~>�?����r�T)m]"g9r����J~Ze��2�^4��,2�]��"�xk�"�)�R�eT�k���F�;�@S!R�1�c�2@�}�͹�rE����̏����.��V}�f	���r�������a���nc��~�v�v��K�Ʉ�?'�,�P۹ܐ�E����)���{}Z��*�J)�"�z�))M�4��⚊��u�-,b.KL��(2��tć�-*��x���1�ڥ'2��2_�G������#���Ǳ�F����]�Q�[�;�(��CX'N������cy1tiq��!)�Lc �c�8��>�$�V	`��od�ۙ~F8��Œ6n�v��p��Y�S��0�^n�)�e����1�G��P�r��m�)���vasݯ�_������t��������6�c��M[L��4���d�x�v���5#������|f��.%0�}�+$�Մ,��,*3���N�!{�}�H��u{1�E�0l�Hݩ���r7����	���wn[���-�(��lja��F ��_��B�/�$��Y�k�֝-��}�2�o~��Ig%��l�m�`w���]��#�޾����6?�W�� <q!@D	�'�=�0�e��J,zE��
����Tn��[��Tq���	�l�.�� b���!�ikP��~� ���Sz#Na�H��kL�Nv�x]�`��E���x���1�w���P��N�j,�[������W`Ql�8w��Ⓢ��r��2c}\	
S�����s]�ᴝ��Y�J�.�2�
f�R�,f&g��!�7�USL0�G��DYͤV���P�r8�
i-47c�x���AR�m*� �~��*�x{+��U>���5v^��=�!�΋zk� Q�8v6Myk�B61٧��QE"G��8�	�C'����V���Z1wK�]�]��(3�K$�ʾƑ�&q)���D)0V5�[r�҈�h�o�qX5��Y�G��ZS���%¨��`p��*����j��	�u�;�~�MGU(�8�1E�(hw�.A�o�p4�}��y�K��ɝx#�����+�Y��9d�����9�@�V�MQ�8&V@�d6фV3��AW��FQ�e�"!�z�����@�H$4�0��x������H���x��q��?@ۈ���z�H���7��W���ΰ����#����t��i�	'�̋C�r�� rT�O�`)���i���n�p�⭕u �Ps���icnV���~��$���-�B��Kh5(��g-aQ�S�����-�C�LS��S�)��w���-JN�!I�9���_9Ͱ�%&���q�� *���\1#��`��Aۅ9D����R�Gx�4Q4���n�����L�A�<���)K������aJ�Î�U��^.�J3���V7$o�Y�m��I�$����;����X,�'Y����7��Ŀh������BD�oޟ�\p3$�	N^�|�CV�w�"�(Cf\�?&6�FY��s�ώ���t����s!�i��؃��a��E�sJI��B�͛��u�c�	��sZZ�JqP�m9�/�d�5dB9.�d�C�G��%6�v�3����5Y���k۠���3��29�?��#R���FT���O��V�ظ��݁�k�����&s�:޼�H�*[���	�t%q��a�������K���c=cV<5� �|�p�Sm\j��t;%�aW0���[N7Q�۫)*��h�(���tL��c�٧��3����	�ʞ޲�Ax��F�d�QHF'�8�΅D�W)� �ڻ4����5�vإ2�T�\���2��(��"��L,�6�rⲕ� ��4�u6�<�K�{��7��$����b۔�w�[c���>����U��;����t��?��Ð�?/������}Qh���R��.m?�*�S|B����$b�aĞٗ�a^��j�<�� U@�vǧ���	���:�E6oX��hl�ǨU.�E�%B��г���?1
��I����
��m�>/�$�k.*x��^ ,��G�Y4]'Π>6�h,7�0���Қ��X�uƁ�
X���[o�r�ܜ�|#�ǰ���ʭ���j���h6�ޝ1�P�W�?�L|�n8��������&��ŕ<����= �i�(6���:��Q�؞�~]@.6�D��z��&�%>�Y��~�-AZK��W���wy�
 ���#<��}�2�]{ё��Ov[}.N2e�#i��qc�4B�a>��ڵ[�������t��M�\Y��c���2�ٌ�����&;�ϱ(I,�v� y�I�RUZ��#{7�e[��c��BqNЀu6������4q��*l�����y���r/^��S <0V���+���+i�o) �%���'�in?=���,0KG�ikWC:M�G����ۢ�qʭ�k���4L��H�V$ǽb�� ��!�?�w{٥�-�P*��>�x������d���ڱ���#�����eUD���C�Iz�a���p�{�l�
;pN��<烬IuI!�o%���US�~��KT\�S�s���nG^@�[� 7�_}��O�
l�c���R����d j��t�i�E�Pe�;�2K{����I�#��7�oo���`k�jhh���s?<��Op<g����XVQ[B�*��{��<�S�hm�C\�¤�K�Ki��h�6vϓ6t��u�:\)�L)NIH�QГ�3*-��D���J���L�)��a0��X7��?��-�[��d)�0Y�jc{%����E?�bA����RKX�3��-��F�]��l6Ǧ���U���ba)�=X5k����֐bJ�:Y>��c@i��#����(��I��To�V%�Ͽ��ڸ���_kX�G��������>%��
xl��IwF�
��qIC��p��4���f�4*�P���GO8�'�cf��⇏o��{5 ,*�*B]>)�N���wa]�_Kܺ�֭��Kb����m�$�r� ��nmt��[�7Ɖ��oL��E!nwC[!�c%a�>9����`�=����-M����LG���n穛�kV��L��%�[ɡJ�6�Lu?�7�`���r��K='>*=?'�Q�	_�0E�S!2�n�<�����C	��Hg���t��{�����
LQ��U�h��[R&�:
�m���O�	</����:Wv��V����Ċ��@s�ڙRU�랮�B�^��!����8��&n��>��lc2�|<¶�tg��hS����-pyQ�	������q�,�6�q�1��[H7��s�ƪl�ɛ�"�Ho��^��`���'c�*��^ò�R*A��@�	�Q]g�EC� �I�L"=��B��,� �
gX�L�%��䋨��0���E��_��\)�*@�Ki8}<��%�3����!]�����3הL��X�m,.�Q�%Y��ܜ� yO�&)�Ŵі�	�����-�������Ii5������*�?еH���|X���N���Ao����%��(�]�yH}>�q����7���ks�3�2^����ITHZ�&�.�u�8������k&����1�[K���]�Q�w[�� ���~�p�'^F맷@M�9�j�U��'�F#]H���&9!D1W9��,��1SI�k��N�٬2MȢ��0mv^n��?��Ej�)�ehu���|4�����/�Z���� �M�s�e�{2�ĕ��1�'�k�ʲP����KL}F�E�W�-�5\�^�0d�^�A�߫l:�!����7J��G��`��`⦜��"\��J���}>ѩ9�r��=a>l�Dd��Z�u����M�.����U��Té��5ʁ�>��wH�ı��v-%Nԕb��f<����PZ݆z��8�y�EGVp�+b�&n�m<�0���z���9^B�5�����`7 �}��6�4ߤ�*>���>~�.���6�)��ȹ��T`kT#?�p�[	Sۻt�_��J�w���Q-˜��-"?U��d|�#m��9�KkF��޿������a��?IY�0��CY2���>\�������K#k��6��C�K=9�a!��x��yK�<�מ8����#�G,���,ǚ�j����zd�8�io���'4Y�� dbꁖ$�a/�#=��j�XW�>��ܓ&a ��p�|��F��Y�)��MD���e�,S�	��54�������+u�g�q��Yh�s�Jiq�1z�����D`�2��\qj��{q��S<jW�2-��g���l���l��R	7���B�[9�M>��D8<�`�D��͗ȇ�hN#�$�g&.k1�����9طvr��}���XJ|������Lzy8�q1�R�0[���L��'����4�
F�Mͼʭq%R�H�O^�zP �a��7OO+�K�&r���)��)��WOY%�-0���jAJ��y�O���9�����\�Ȱ<�쵘�Ŵs�ۑ�o��,@'O���Of�p%�R[�k����!N�;а�2tk�=ba��AM��\l��X��P��,j}W0d�m��AIr���r�G�����vs������v�KY��¤�0��#mᧈ2<�'�b���BO��7���a���p�Z2�B{��
xEk	�U_x��7����p����Q�qG�<����7���K���(EY�<��T���x���K%(���+Յt e�9-�zk�������Ҁt�R����]mM�t���^Ֆ�|��r���"�I��-�����f�"��ԭ*�3�&M����� ���d/v2�36�,��`hС�O5G/��m؆A���M��A�?����e%ύ������&8������W����$�ؗ�n�B
H�&kNn�W3�>�l�80�V�U
3SdEFD��� �L=#?�Y&�#7�Sז�}�ֲ�µd��A)��5�𓩒%ӭ��0lE�<=��������
�NY��w��� ��Y�;r="[f	���������T����,�#W���V��BX����KD�P�������7K���e5_�p���n5w�Wu�<�!@M� �������a���Bd�,@n㊧mj��C !�%�]�z!L��Npۣ��� ��,�,�uV*,+\fX�ai��]�Z�uߥ	���c"�2ߚ!X;f[i(巕�T6A�9�|yХ1[aXY%���ZO���_�<�i�2jtL��;gԌ�D�[,g��h�$����N��+�	s}�/���xd�d<��d[�4�x~K���=������t6j�Գ��n�0ϤߛëY�*�=�_��$r芸�3��p��������Al�D�w��>�ޒl³�����?`�c2�էS��E��لe���ĿI�.�La0�Y2w��J�mL�.��L�)(�&b�a*��5Y.���) ���rI
Y�Ţ���݋�F$A�O
;>D捶	�b�+�����ւ�CKI���NL��e�����9�Z@XY+w�=x�|WM��uru���#�(�<�'y�G+[f�N�*!����&��8u���4�s�\�ɮ����8�
�+x&�5r�	2l�9X�����k�:.��TénW�����j���"Hi�Ӏ����m�����ťQv$��{6�!�?�]ޞ�R���M�A
��}�~_���6֧�/�4q{�*�a�N�j�2&q9><�~x6�I2y?����m�?�tv\eU�.���3a�iD���^��}��
厸t8�.rV��Qpi��f�����Z���J�ik��x3=$��a䯂��%��E�MI/����i�~s.xH��h���'��{��T������Q��]�r��1$�yt"�}s'�.�xEI�|3�f��Nx�
�yn-)�Ͷq�<*;I�ֆ]C�& �PGeϨ�8n����I�:c:��ԓ��0�B;
BL�*¢���4��W'�-o�y��'n��&���]�^�.�T��>������@=�\�4�pK���r�z�XfV讈���G�
���g�4BLDXl�
S�Yu�U�zBL��daΤ�!�;Vdآ�ſ1�L��:�$f���;��Ꜷ	��Mw>��kd]̪�6�����&�����ߎ� P!�A��4�J�*�b�Uܦ*�#��=�P53�!lS�t��@è^ä��%�q[�!��;ГŤ^<��k�TRͻ�
ߓ���WE��B�5��a��-R��>�٣온��ԁ*�H3�<H!��\*�hA!d=�h�����P�Xv�Cwg�e���`ĳ����M�iX�����>+��$+�Nɏ^�bWFf��@�K=��#��h��<W!��izC�^j �$�x����h��z�lŵm�?�X�lT"���Ѯ-�=���N�a�56釪����mm��@��J�Ա�S�?]���?į��'���C��Qj�+�t��y/�=ב����Tq�f�Uj��0��9� OĸG��� O�:�\;1Ǯp�$K4��>]���~A�����V��νS;�ġ�t}��� �n�x�
���1���y!�Ha��2%��1�^C}���§��&5�>YY��������y��F���N�2���9�/��E 2R�����e����Y�����
�du[c�)�s�.ω; -�9Jۚ��Z� �������*(��LM�Z@I8��� CK�.z ��ze⠠���4GG%H��ƽ��=ŕ����X�&ќ]:��ޔ5�g�����4��7wSZ\r#0���g����^:�{�&�h�����@9�]H-sG�=����* H�oH���ɒ�j�W���A�gz�IR�ᛃ��t�j����j-��l����ǽA �|��q���0���l�Rfv�!�+��J(���Қh�l;8�)�ڈ��y����sʼ��7f��j��(�9�n�ޛly��c,g�Xu@-!nӡ&�H��p����\��UVKz)�á�1T��G#�~�~�W��:Y�,�?R�̸~�����J�Dh��CqL��ת�E*x7AR��q׆j9@ǿ�4,������X�wX�^��N��%��l�ٍ�
n�e7�������1x���7��Q���;�n� ���@��j���1$��a�8|�l������۽R��Z۟HuмoJ0I�G9\�po�b6���۸�*Db���놥�b ņ���b*n���j4��o�;|�k�ۭ����w�3����C�{��U�������=r�۰��P-O��~�y��`:s��7���w~��Y\�0R��ȍ|7�a7a�/�9S�����8�Elnr������]�yҮ0���X���)O���"9*�b|v���k�$ ���tˊ��÷͚��{�x�{�l�h+UPy(�Ο؟h��f��� [���v2U'~G���GdX�"�zpU�M���9xW�R��^�iN�ͅ *%����t�@N;�g�4ck�Kx7����v�C����ž�b�� >6��������n̗g$��K�b˫V^ΐ���0���ܰcY<����L�����=���ܡ������lE��h�E� #�<}Q_ʼ`,�PJ�"j$�`wx??Q'V��C�?�����*fMn���/sw��=^L~g���*�X��?g�èc����G�!3�:��XDKR��H���/w�|��._U����%RrE<Ek=���}=�
HWB��~��K��B��$�r�jjh-�5����({eN�e�G�ͫ���BA�Zu��֏	;uC�������z4,�.�x�Ơ�^w��
~@Fjh��j���	�B����.��IJ!&
4��;@iAE����a��XD�{�\�_����/�c.S3E�o,�%T�@���x_*�4�)�BT����4�]�>�T�m��#��і{M�i;<U�A��t�h��������b5{��zyںI�RpR�y��˭��ѩ �:I�)�v;��`���O1�s�\��둞��I�[B��ܧ�BC
+�@	�3�O"��t$����8�>��Y>��𥇡�=p�۲�� �w�ۈ�6��k�����-{Ĕ���*6��5/iww�Ē��{wx�!�G�b0&�q��n/y_ly���}^��|)a�m����(�iO�S{����:<Q�X��m�xO"6V偕�KĽj����18���E��GL�1|,W���FT 0@p�9�����a�B���KNJ��D;�E!̾��ξ��I��I8��UKL�%�󈭕��ձ_�- 3ҩ���^�k�0�%��rr*"V]ûխ�A�4��B����E_�������*�@,�f�-��Zy�=����jd'�ټ�Zw��������_�eh�ǊѼ�{��!y���{�����IM,Nz������8^����;7=��Ҁ�|���q�Ο����~�U�����415u�=�:�=��R��~-�l6��D7���'�C��F���ֻw���:�.A}�lz���Se�-�B�<��`g*�5�h���$9���p	5�s��H!�t�F���1Z��oƌ���zv�z?��X�R[ �ҵ�&�5XBggI���3�Ewbt_�|�%N8��{�8���r9�V	A��}i�D�=����R�t"U/�A����uSž�k���ƹ���f凟�m��}P�
zx�-��fqZ0�Ob�p��K�<�g6�M�7������!���sʠb.�ۋ @�]o)�T��&v(2�J�H�ܵ�}�z�.ȕO��؊-��!I��u70 ɠ�	�Y�X^��[<Dâ�(Syr�ϊ}���QnQnJ����Y������fޯjC5�{a�%#�d����Ux�(uҶ�h��/�]R����^�(@�c�d$����ř��L͗2݈�Tn����I|���I�.�����$	���y�W��\돵���4��y���C�t-��*�sIe�y,�l�~򾅲��j��:���_;-d��UM��Y�d��h�+��D��~W2G�jm]R�_�`�� �L�H�_p��v-5�o� V�c�8�9�>�Ϝ�z)���WM�1�m�G꽸͉'��7�<-�5 Cxp7�T�Dd�p�d�̏8�So̞�oj�"���"Y��}������\�X��|�ߑ�M��CTm��� �/^Q���*��������;M ���O�8�î�a�yJV��KU�����H@0ꬩaʴ�Y�^:�I���x��FDٌX6���DM�vZ�
[֡�5�bK�2�*|����⿭kY��A/�=���zjU�h�#�kÉ3C��\V���HN��%%��6���j�3����>@u�>s/�O�`��T���_�L�k�O�@�܈uӡ���J]��o��0��c�D�UZ��C�'�d}}a��5���]���Iw��y �[��M!A�q�%�t�iZK���&��jJ6�/��\6�?��ٿĺzV�gIcsŎ���EO\nS��#l�r-��߇(�v�@�,O3#�.ǫ�AQ�gh��zb
_d�֦�B=P�A��t��k@`�G����:އ�)�n[Tܵ��n������C?R6 �I�-~5�T;�[�M�Q�aXK���7`����.f�ǘ�L��T�����-�@	H�Kį�xSs���͈��=):�cf�vK��z����;?g�g�����FtW�%���-ު�_φ����/�3��\��-�#����Zm�jZ`T����X�ӕd:8�+�>c =Z����N����,W~@�S?@:lh����µ�z��a�5�S����x��SvϷ5�J���n�	^Ne/� }�ЙvD�i��\5��Үq�w%�#���T��TM�Av&�!H�7Lm�*:�У���7��_����RX��~)�p��~2��m_�SI�gB��S~��9��]���~����B�5l?-�C��l��xw�2���%9���{�a{�>$�����p���g;�ȴ����e^�Ί���4���r�civVX`�=�������m,5G����\"�Uj)���Hv�N�19�#�=�`r��ɠW�9e��H�� �:Y�ǉ����<$�C%r0	+-/���������8�6��l�W 4������:c� ��2og;��ߕ���u=�v���A���f�[��[uM$W��u���O�%��}��~��?\ ��6�3s�ai��b)·[�O4h���ƅΊ��b���Ga(=iؕM���"/_zdB��9��v(�g�Jj����gLݭ�<:P�)�˵4o��8������xa/+}��5%�87��i�6Z_}|�`����a�eQ�_ߢ�:�o����31b��܎���f3�K�lv�r��ij��~�j� ѫ6c�Nz�� �c䏁�Jס.���%[��� L�K����Ӈ����o:�&h�ة}j��ѠKީɺ��=�����t�Ӫ��U���-��R�@��4��>rY��_߬�n�@]�y�Sg�.���a,��_�)yY4ʾU.���=c{�z�fK&���3@�{U�!@�r_��^@v��FU&�	t�±f=ڼ�\/��i3���������	�i`#y�h-��c�Nw�_�<�r�yzk��Y���f���?(��^� }���?KH��c&�;�
(n���8���z(7�}b03�-��!��ג(��:����V�������cd7Җ�4���� �_eH�L>}���׫�p��pQocF0H�|����œG���8����׀���t��y�T�듈�r�_Z�F�����|����כ`D/Am��:��C�n�>�d���\t�Bz�}*��o�c^�P�l?}H�Y&,�~����U6{(V�n���x2����dVa��\�} x(_�;�4Hm�` ���B�t[SK�����A�L}\�`o�� �kfuxs�S89ݽC��1�������[����#)�8/�hEi&gg�1ٷ�h� �o�t���l�w�vn���h̭��ОO���.u���o�w��AŻ��Vb�Kp1H:N}G��n�?��!9_����Y�&�P�l�"�Qs���f7������ʂݴ6�ur�4w�g8�W,<����/��t�%g�fA}�jl=_̵�
{�EM��)��Y7_#�>�.Y'�8���d�`���;��?.FЬ��r5x:�W�w�?i��s/� dhޥ�P>;Cw�ۓlP��^�YS����s]�1e�#ه�Ygb��zn�vO�1<����_�����lN��!U���{\+x@�0Od\ͧ�Ȋ\SZ��\�.A�M?�!XY[k\	�㫰�u�F�\�����	@�A�D�h��CL��v7�x�UdTj��	f�!���Y�х:hmu�mW��%.���r׏#o�:�*U��Ǩ.mo6�;h_�I�����Xa��,j@3>��L����|�Ew��33�tx뀪��/���������Aj��2�2c�\&����OXD��ݻ<�Dk��bm�Ku����7-�oِ{�%6��%.Q��E@�L� D�g���f=�Wj/_ O��*$�����2����Z������B�8����9 h�V��v�#���Y��S�:�5��vh(v��-�ѫ�'\��gOk �fĸ�R,�q-�ߢ�4
�Gv���8m��'� �,	&���L��̆��R���7l�5NӺ��\Dvuא`pZՆ������Ua�?-0�L=>�6�$�)�8!�w��r!���M�D�S��b�1�ٷ B@D�^�����#�����������I��p,Hʟ���� �����k�t�Ǡ��u�,��*��Dd���ptI���,�{�Ȅ�����5ț��p�L) �\Q��������	��h�ӌޙ��X�$�/�m�����Y���'Pw�������褝�:�@ˈ�_7�LpF+r4s̳�-�o��l� �{E&C(kHk�϶��td*sX#��+��k��� T+C&{�&��T8r���Tf��-Uo�4�~�2���:<Q���g�������)���N���͹��
����U�7����g�'��p]Af�.]
>l�K4d�ߢ�&X��/��km�(�SͶlC� ��3]́r�p�S��w��m�bی��à]���G�6��r���o*�hIS�#gғ����[�O��(:#3��:�A)�z�������v^ۃ���1B|x��Hɭu��zy9�؀O��
b��z~�=����&r���(�Ϫ����{y���.�Q������l���ʅ��L:Y.9F�T��s^����,��4�8�
-o�Q�n��@M˽4�=٪"�s�By�c�vA�d���Vg��N��w������}�)�d��yqI�����H�"�n�B.�S�t��\�%�\�n8��
���°����N+qI��e�M�B��[\���]U5*u���u�/D�����W^]�E^S9��-[�x�]w�9a�$��?t����Щ�M��dE�8I�i�Ⱔ%+���Hh�a����۹�S�qc,��'�]�q]�~����Z>W�0�翤��8[�Æʄ,��Y���q�C6u�G޿:+��D��}Ŕ��jn1�+; �b� �=9�_�j��w%M*�Ys��T���-l6�~�ڤ�&��V(��H�U�W�C��^�#g�)�\^S�_N�]=�M�_��.Q�l���&�����#��N��uyϕ߳����:'E��VK�lgw*���Z-�L�'���ۈ�vk��9ͬmt47D��OIS�b[�h;�f�,U�䣆�$�LM`�g2��ց�[iZ5�S~i����~�@���u:����_">G�j�:ԃ�lZ$}�n�B���,n�Y��z���b؟�sxǑ�k���)��u="��i\8����>�s�d�H����$�	��%�+�7WT{�������˾Q);�d)2����zy�
�l0�<$�Mn�6.� ��n�b�\��X�Y��~���X��:�`IO���̣R��tr�YkG����m��൬�[@��.��xkv�<��+PxOH^%�OYT��
m:�Ȭ�<�ۖ�5+���Ӄ�o��t�:ד��V���/&� �fp�oL}*nQ������: �%��hWf�l��tH��"�	���n����g��(�^��֩Ew�o�UΨ��_E͔��0؞����H� ����IZO\-FF��~?���P�݈R����n�}Yz.�xoҡS�oJ�5>I�<��ɞ`�6guӮ�>S��c$M�&Ɵl��T%�/�^3Q�����%fDʽ�L��:��S�݉bߍ^��8�a< ?5Sj~�i% �PG>͂�$�\I���DKyNtJ�'=��-�6JƲ�[�I)���9 ��C��Rj������m~:f���.�6Lۂ>�	�Oy�*��{D`�Qz�͡�:��Kߗj��OZp]~/Osϳ�ԧ���)�F��qHe��əR��a��R}T��ܬ �ҕ���|F�`f� Of�y'�
�^�c`���k%KVk�	�o4�5���<a%�ɋ����:pm,�bA&8@����H6�uq =��I�p�ll�dS�n�`{��'��~N��p:��M�o�dTa�S���Q8�M�%W���v<uP�V�-����I	X�%H�K�T\s�7��&�9
w��>rg�يP��)���Z]βn��ɋ��YK�&����Y�nXxA؂ 5B�,�ٰ}�Չ^@�N�����HN\���g�c�����Ѩ1�Th̔���!�L�:ҠTH����|�����E��J.�:�l2�(�u�D�c���z������*��/��WB0��E�&�>��Luެ���A�Uܤp&G���rݡc���ME����'����xs@�u�Ba�@e%�J��en��^1�z��Ӧ�"�~��+(��R�3��ۑ���T�˗� �1��Z_JE-.�ɹ@J ܙ/�jN�@挔/���_�)��9�wbD ����!���E8�{C�5�|_��W�sw �.QU�'R���edo"��� ԡd��?xQ5�;HJQq�N�[����[��/����z�����B��	�����Doo�M�bH� jv�^8C�m�&j�}g�Î�Ycu�r��|P�A�MX��Kd�g&�f��C{�`7Y��������G��}j�m���p�&�Q�-�C����¯А��'�r��$Z&	jCf�s4����iA�]�:�B��Lrnl�c��o�r��e�{R
v�����<DP��/������-:�c�I(��"�]~��nX���� Z�7�""�c�4���[ 2�?���}#��(����bW�	gaB�3�л�~��H�Yi�����_� 9�������t��)2l�!{b�B�vf��C[,�d>N�+R�V
��D.�+��.R�S�xd�t��%:N��qX\U,t�w����J��3�ͩ�1�L�fy�����.p'����w3�����푬ޔ�����JȜ�|�.a�.h�s��$���M�Tv�� � �id` ���U5��bE�Qme3:*Q8ԵqG�9����h����6jn�
��$lX�Aov�e9ԯ�\�u�<����`���4Pkc6:�9;�:0�c��|(M��ά��(G��}�@�h{^�c��W��T���6a}��02
-�?�y<�9/n�9���y�IС^��Uꈍ��1ccK]��dM�_s�i���C�2���4|ؔ��N�.{@��0^�����S�.\ǚ�����FT�>N4w�q}zE���y�$R$�xu^�x�0�#��"g��_�;�^6R��4l���ZUvWA˨rO�#}��++��ֈ���>^�� E�v�/���d�cw��R w2K��d�}ͯw)ʋ"��@��	i�F�N߈�K�k���������z�8
#��Z�e�KW>U �r�+�c}�6,�<�ۅ�N��l��x��Xd}d�*�Q�l�M2s���n�"L��J�ťb)BWX�o���:S�!�$��AΐU��7�s��eP&/R��@E9G�!��ڗPq�V\U��;'���{<m�D	`���ί��Hzq.5G7�}�`��9z�Tg}�0�e&�n}M0�xFP��T����\�Zy���q*&�5�D��,8 ��;�!s^CP����y�.�[�Aݻ����
r?����� Qg�Sڢ�Y��@�BE���C�vǑ-,[jT�W!q�Qjp܈�'�#,�h��9���� �:w8�v���z��X3���lN�����z�(�j�ᘢ;�@��
���f���S&��f6��d��T�y��6l��!������zA�/B���:/��΂��k�T����l+6fV6Zd�c:�Rx�����O`���h�p>a\A-M�KF9|V���vZ��:�F����#�5r�1u:D��M�z����ıU�U���1G<�k�٧���a[t{C��mo8��v}r�2�w���Uο�T��&_d��%d�m_Dz���S�pH��^Nk,*�lΓ�>�� �$��L���o�����`�c��A	�q��Я���L˃�Z��b��T�p]�0�m?~9ܐ�Υwh��^�F�7x!ANҏ|�d�o�+t��2��l��������Ә���V���nA�s��)8r�n.�ju߇�3�]q� qĠ�KA�7W	��5�&�*�^��������]�|d(�o���%s�^v���W��x)�S��~U�H�I��S�y�g;>L�9onnM]I؄0�bca՟���6�����laڇKh1�09�S��c���j�|8vU�/�Y$U����� �6�5�7�smߗe�4��.������v�������e_!w��Ȯ���.䁆�B�"���ْ ��P2pb��+~P����]0W�������nVl�+�� b��bM�1�YȈs��%��THz��{����+�U�j��M��8;R�"ֶ��/�s���Q��i3��h�X�O9*����y��`JPF�U���ZZ��ͩ�����6���`��G8��x��i�X^_37*:��?���;v��.��=	��=D}���,��zk�y
�R�҆�!�L��S�D�tvN�~������>�꾷:�X�}2����[W�
.�|J��a�]�K������}{k`�=�>�]~fc�>G��&�ۖԏ���կfC�L��__[:�x�q��ס�'�I��	{��	!֤(�D��]͒ff���HW�5 ��o0,+����p-;�o��să����}&z܅�׫K��mZ�*��[0Ӝ]��
�J��0�%�i���֠IY+�^��%^-���`ӕ��`i�(l���.ŋ�{;���Db'�<:�L/�	�� b�s�#�C����i<��H����tUQG��+Y�,.L>LP��B(�O�y�}��	ˋ��� ��-yl�/��hq�O�dD����3FS��<�R�K~�;B���
�\�L�ChK��ٔ��&�
�	Y7�������+�8��5g��D����2��\��R[F0)�XN�r7q���0
w�����]�p���H܌:���B�6p���C��*ƅg� 	��ȔƮ��ź)�N�Ho��;�0�T�p�9/=NPg�Rz�S-�3h�?�<\Y����:SK!RjS�o�*����>�(c��)�tR-?ŉ�\8�P3h���^�ͱ��>h̏ݘ@ӊ�%˛�#~d@ۣ?w5:{S=�l��t�(Eȹu}����'��cZ�C��*�)�E~O�9�D1�ڼ��*�$���>�3�NtH�Mф���d�:�	՞�S{瘋�ܮ��.6D�є��皜qZ�m���&�>ҰԹ�83ެ,���"Dn�j���x��N6�i�%� O��X�n�8�����l�T<o!p���^k�����-�Ն���%e*|\�=|���·m�2e)�'�Ηc�{H�@S�ZYf�i|�~�B�V�/ U���:��!3��j�H	�э�*��МQ�x
��d��#��e�~���JiL��7��dZ�Z��O��v�u�1�V�I��'~����ɢ�dA�TK�$������Ƿ�M�$8Zs�
��K������)�wo;Z�L�ICѷ�B�ш���1���#��2��v�@����gx�f�g��go
������z���;�N���OR��x�JI�g'�R�s���$0,��5j)�)ʛ/�
��65�M����Ԧ0��K�@@������q%?;�g��'�W��*\��K�]�C�&���<�/<�B�{g�� ʌ��*5�Z�-;t�=o8[cI�Y��F�5f�7�?z����� (��`���6ND@O(Dq���|�&fy-�#s����+�q~�� ��l��=P��8��:�)'Io���#E�̑07u��7
�-1�2����gݕ���/���
*�O%N��6��H�\vy����_4p�6����F�|9j�{4s�1�{�,|C��!G٘G1����
.��3���co�B�$P�Ǆ��D+��a@��.��@l$��1�<�tK�M�e�G�ED���G�&m��K��ߞ���0%�DX���n�~z�!�����52���.���p�R���PDG�( |��8�6W���Ĺ�ǠΖ��ZME���l����>0��ʍ���K�E�f��Q��l>1o����pwSJB�Z4�+8 �ke�>�ܑ����ݏ�Q4�R�>p������V*W�"p{�/�ru-���хZ�f�Z�O�2�9��Đ�`h&�\�Rh��kqE���5��Cɮ�=U�b�<i.�|�A񺊏oݱ/$8M$�
脕AWX�`���S�H|�AJ�.^�O�+��&������H"�������I�iy�H���	��=V(r����Z����~��]Y}���� �6ɚ-���v��65?2ѧ��l�Z1��;DrW5�*G��,>�/;~Y!5,��h�M�|�Wz�g����>�b��&~ERK�m�x�oJ��[�7�Td�_�տy�/�s˩[t*o0
w�a -�7��[��۲3vYh%�9��vM���6���q���a��iX@��-��O�L�p�T��E:I�>��q'����㍔�@����
#��%�]��O�R��m���	�z�h2�z`	��!��,��>qC�(�B*w�݇iW{��mm�ST��Ә���O9^m	���[ZA8b�~�����d�H _�U�֧uJ��YU�Wg}�ܽ��>�'�^C�|����3����)�r�� AN��gf��Ɉ��9�5���N�L���@t�1&�.h�k�"�5��m�Ȟ�وh��
@O�'6�U�mcz�ƶ
�[��Ϙ�~}�Q��?��$5k*�t	��ZWi��0��8n����	�-6�U�D}�փ��1V8Yaysf�d��>>�.o-��ó�!�<�u5�r�VoK�-��Q�C��n�N�U�R�WT�YD*��@������dξު6��5h*UF��w*�$��
)?����hoemE�}��@��ઞ�eܜ�
�� �t��G�񌍻pM��������<�2{�f� />O��P5�x�y����=��'꛱�N+���v��%��@G��s�.�^��e1��ٖ�L��������o�&��|�[鉒�� �ι#�W����Po;Ovr%�wk��d��t�4�$_i����@��0���d'�1Ty��w��#������#|];��ؕ��	{:�?0�A�2y�l/Ĳ��[ (j׼e��'4K7�4�K�I.*����~����|U����"T"���/�5���l��&�O��i|iev鑴��|�"��n3 ;ò`��UJn#��y1N�����TN��ٟ^�1TKG�Qti�g�4��8XZϩ�r�$�-�f����"�Q�G�L|P��`P�~����W�������xk-6�爟q�(B�
����LEP�BàB������9����q����0�8d��Ɣ�<�n˒3X���O[D�^v��%tvXǕs8���D�Z�R�A���(��p�N�26�5$�>�n H ~�1���i�"yeȺUI�0��g��`�%J=�1��՝�̎&�J��g�<bW����HoF��	Sc��В�o�u켛Qf���A�5�d'���j0�>�V��2}�`�;u�N\��u����Ir3�K���0ټZ�H��jN���_E�W�X��&l�`Q+��z\��O����8�����LZd����P�3�<��ej�vX��&TZ3�C���g���*F�m�n9!*[�Ԕ�!mZ�ׄY�"jF�lnJ\��#��vd���/��3,�O�����m`�b#��w���?�z���=i~�4�I,�%.�	(ޜ�)[���Kآ�N���!���,�㬽���Z��^�{:3JWS.��0-�K$�a"4�|R��f�7|FCx� �u�h�n�Nb4���:�IX2�j�[ʻ���9���3]��]%<+��?u,���,G���g��(�(d�^����8.b�VZ��J쮣ٍ���xDe��x�h	8���e��U�A�͝�?�*6j.�
�F@=�N{h��H.E,�KXxB���j�4䅓U��O�*Q������ħ����I���\6R���)� �=���q����UА���%�3�SzK���_=M��!�E��:A~`������Dq.�r��5P���Fg�%���@��j҇�?�T����4���+���:Ϩ�G&2�J��se��.b���:y$�A�k-�������Cw�ŵ]>�� ���kE���;�Z�`�W�^M�a��[R��Ԥ��G��=���ޅl��IP�$U�: �ZA {vT���Uv���}�{_���"H�RV�Z�լB�ǲ�����&,I�2�.3����]C�x��`�gq�W�_'DE�r��z���1�Ȝmg^��|���ÒÏ@6q`�A](�����wU��Q[FiN,��)����� m8�nw��7�ܙW��5DB,��fQ?�{�A�ގ��N߰�r�W�r���>��h*y�!lGn%����Vsy�똁/�7�Χ�.��x�AC<ߣ$�|ȟ?,�� �=q�\�cY��.]�=C�כSmc
cN~%�}��7����g��)f���8����\��� [h��b��WD��kFh�����L��!��id��:� J����K�aL���Y�cy�܇�/������_3\��Hb�Ud���Wp����S:/�(�J�UZ�J���8A�L�}0E�PȦ`~�"{�Q�\����
)�
�In����[��1�c0Fz��7Z��
��M$�̣&/E(A�
�cfA�k#(a�-7������
i��/�"4�w1<G"������)�(g�x[�����F����O�K<N�&��Y:$vVѐ�U�Y��C
��Z�޴�>a ߻��
�9/�FU~�c|,>�)ۖ��ڼ�3�9��)4�`�̩�)A�h��TQw���}�C�6^��2D�Ǽu�p�Z��R�;I��p�X�U�P��cD{��L|m�s�~����9.6p�I���w3�~����L;rcQ�^��Ҹ��R��_]͖��^�8@�Ze7A|�$�J��:&���e�m� ��>S�e����W��=I��Z�Ke`��,���e���|�`EO��	RV9qRwjN�?RO�(ߐpB�
+������f��y��~FK���N���]����ٻ�4���_;���±�������6)�;��b�&�y�_G�p�j�v4|ql�K��=�qq��i�"���A���ɽ1��·K(2��C���)���
avT?���H/c�$w;H�����I����{�gPfZ���#0�[I�w�#�)���F�r<\� i] i:'q��P�s%�q�a��4{Ns�K��t����a�
��.�5��ßE�� =�G�+@�s�d�b"��t\���s�/(��2�D��y{;�Y�:���ca�j���F:����03�V���#�ۃ�i��ʩd���v�L�����i����0̨"�g�3z�WJ�����L�ظ��!Ȃ�#��"ڸ�k�kV)������na����W?�-�lD�"t��'񛫀���aq��od��@3�+k���WD�x@0���1T��,�x�5�"�d��?ikuO�4���f�3h�2O��Ň����f�.d����7���Uo��f�I�k�.M��Fʟ��	�g������!K�
�Rt�AnY����?	��Abʻg���Z~`�7�!�V��E���`�&��~e�������љ��pN�uZ�q�����Wz��l��أ}�����7��kEɲ��j�b�[��o�OH�v
ەd��g6%�z���a!i�WZ��^��ܫ���y^5�X�s=��{�;�yIxU��59�G}�%.���5���q�df�/�ѣf�$摡��������cUj ��&�'\j���.��y8z�E�B#���Bt��m���e,���0��t��D��b-W5��nB���D���_'�+�IbAt���;��1��݉�&xF�%�=i�#���]1�ř�V%T*4��J\�?E�Y �[�@�_n�@t�%�}8H,�X�2��R�%��!ڞŋ���K�8f����8ߨ��&Y�	���z#2 ���߆%�"���ļPg�N��<X\�"0Òf�P�2��uv��+�]���:L��3=��v���y=���n|p�D�6`���Nڷ	�5��l� ][�ݏ�������b���f���>�T��Y���v@D>Ϝ�Ю�E�q��>VԌ�O�,��t�LA��v���jƕF�(��Rr�R.�Dt�r��p˖^W�P���r�ɔ��?[X�d��UX�����(1��1g��4��ֱ՝��uC�1�� "�9$� ��C����~ҫ�
��?!���e�e|sfN�L���YG�K)���쐦�v|v�؜?��{�:��Q��w�'l��Eq0�������"��[@<�g�w\݅o����a���3��"3���������	'�03�/6�ۇf+3�$/���^ox��D���@�$u�|2j���������� �Rǽgh4�(3�X��w���|���c�%�����;p�ߖ%Er���{o���[BF����ʉUR�l?=���Y���q��[C�2���dgg_�ME�A�w@�]�0nxGv��[�O�Ι׃i3��UwV
����Q׊�	<N_vo���Xn���W�b´�<2��Ԑ*Ojyɹ���=9���Z?�1��3��<�\I
�Q�>m�Y�g�30�'�a��+8���J���v���ZL�d;���(�M�}/.>j�@���V�ސ64k���Nf�\�Q��>v����M1�@-�s��Mn���1C�u��CC��xas
�y��'͵}�PQx���~��t�~D�٪	h����	C�,�9F�p��L�t��Y#��5���I_pȰ��<$�;�D@d�*{���c[(�[����0j��ax�-��T��Õe�ٸ������Qt�h���� ?N�����d
�jɑ���F�}�Bڍ��=�ƃɢ�����c�a�����UO���p,Pc�8Xg���,D��o���.C�����%�v���� !���^�q�g�g��GZ|�ɸ�̀\�͇�D�ʋ����ە��~���ө��$�9�';ܱy�E;���[RA�{���G�ȗ(�qsCDEyUu#Ė���V��_�G�gC�wOD ��V��{�V8Ƨ<K�V�	�B�G�E�ۧ�C�e�� ��
�
Ǿ��}y���B�죇톷���`Ր	sO	O�X4�S��	�������RL:<1�9�^�-L����!?$B'$�c?u�W��ѯ��$:K�5Lg���82��Q2YV�\����x�2�9� ,�DY�{��o%36D���M���������}%`c�9�
�q��fNy/)�"���˜��C>�˙�$��#0P�l��=#��}�[�J(��cNMl������g�B(.~����8�"��S�>�xm�S#� eQK���N�2�1<���i��'�48l�!w@oo`��5�!l�&��&���$NY��.�vhd}�.��GQ�-�˖QS�\LՔt����ψŠ���=��b-�"+���m���b����x	d���o��X�s����B��%|�2z5�;_�=x�Cu�R����`
,�0Wp�Z�$�[I��*%h���3���ƚ���\�����p��,I���-ߤ�_��7o;䋟��w���ҠӇ`{3܈1=�*� "��*Ou}�6A!���؍��ٟ{x�����E�bu�#���_)"A[�;��6c
���+f a���vԡ:�z�V�� `%�J5��[�2�4|�����7_�{1�O}��2��L0.��O���]mM�ȏ�9W��Yն�2� &L��'yb ���5p_�,ϕ�q�X��bzv&S	T��E� �Ը����%9�i�����!�V�~�ͱ�k�����+����U[�&䊶Y�Y`��
G�>�E�&@��ʴ�����y|���l=Ȓ!q0Z�W=�a�7Ld���&�%�;<��E3���8�;=���p��$:�MZy���A�B4;����#���x��h���Ě�8�q�Ǵ��b˷	�,�����}M����	.� �&@�3��K�׊��+�j�>��B�vb��-�m�xMBmj�]��!9�K�z��N7��ߺQ����푢A/���Ĉ��Ė{�Ԟ�J�<Oh�Q�<�i�?� lK4D�+{���Uӛ4����'�G<TD�/�m\%E�/l9[���&%��gJD��DUDTٙ���qgES����NЬ�=��79I[W'KA������4�~��иOkWS�'�қ���f���<����B�0��g�h�=3ZZ�O󌽗��=DW5�N�{>E :;C�Y#��$�)��#�tD+	Hɼ�ox$R��r�����'4�#����˓|K�)�¶V���%�~3�� �R�|�;:�#���PܦK�~�Mr�z'�vw�<��R��3T��m�Hh>)PK�_�a[A	#z�k�e��g"6Rcw�+s�&���;�^.�����!"��A����S1�!�7�����`�`w�!�A6i�_��Q9+�/M���G���K�YN���x���͈���X3��,��?���Ty�U���]a���1nM|�GQ��);ڜi����+%�^�b*e��tF%��<"����5[�TeO���^���fxM��Cv�A7Qa�"�'+�^u.Er8IsX���#͠.F\lo,R���$ɵ�Y
���K�QŸ0f6J�r�����sy��"�/�3VPlO^���Ы����W��o5X\S�D���DVA��X�b?���n[@L�5L��V�}��?_	Q5�4�꾸�g�A�<g#Z"�&�PY�Dc�ڑ�s`�`Nǁ�N�ۜ��z���}��i�Xa���u#-��5,0�:��I��[��O��#$����	���	���K����I�%?���Z�n!�+u��������D`�/p�+����桑g�w��vO��Å���w�Z���(#3��x�^�e�3�R��w���Ƹ1��1J�8�^�y�t,�;���������7
Jw� m��`L�k^��7У=�l)&D�@]�S����~o@�hr�V�8_�.��q#�Z_V�3���Ӵv��L
��$�VC��c(C[R��n�pOD�_����b���������P�����0�mW�g���p�"��I�Դ�y^���7�?�v�����C������6������ǈ]��k�4�v{u���/+���Ǖ���/�!�C�)���	;������V������B���5����F-�Li�9-�8c���Zq�&�e�_�g5ߒ4�.?����WpAf�������Jh�i��$8�|U�v�9冣�+��� ʙ_�D�Ѕzz!H���c}m;ǉJ10q[.:���@v8-��њ7��0�Ɓ�S�y�T9B�r�
�54^<��Q������fx*I�2ѳD��:e�����ѕ�k ��2T��	e"�K�Z��8�+z����N�[�d0ק]�:��ؤ���k�d�lCP.�]�gL.�m�>�TJ�-hE���%�~�(.
"T�x��>�-əT?pV� c�vǝ���C;P_���� ��
��b𥒄p,d!ބ��v,��PK�ˤ��R>��Y�Wt��+��&\�"*0g�r��
�9�xn~NG�#��8�
�AY>x[�(��%}mV
jF���GƵ���+�[ϔ �ƴ�&�<�\O�[�u]���Kb�{zw� #��Q��N� KQB�-FH���{�[��ic #fsfO��Hc�e�*6�I �0{:���yL%Z�����/pǣ����\��U�۬PxqB/��� 	�R䔕i �y�:o"�Ş>#<Ҹ�|=�@�Z�A�t:IF�.*�W��QC,�.]/�[i�X/�߮���1X�{�4`��n�I��yd�mU?�}� N�֍��L��Z�����Q!�Q��x���4J��<51K�I��P�Y59�^���)K~k$4�+L�f�*k?�ڹ�z��Vk��R��-� V���M�fn7�1�C��9�6P,&��)��~�L6�\��?K�R��Fy{J�|[>d��˙�*�pv�z���ZW-2:}z���=-��Z�&�U����^�d���֘������S�A��=�16h(�ME׊>��I.���H��� Ш�h���fp��o`0t����E���
�M���\#25�/�[X/��?}�={��Ɋq��w����^}��J��E��M�T/rq�̵9���d��ܓ���7 pS�#l���}:�*�}�1���G�O�f;�Nv�ǅ�r�����^��-d��&��1;ƙ��,��&C��9�rC�4�M��+�Ӕ�,Ƀ�]8&����öiv"���L�JE���uӸr[�*�x���q��WNOi5 (�iyw�S�k�İ3�]�٢!�q<���⯂��j�KF<Z��?	{萝;��s%.x�?W�Z)���\�p7l�n%�RX�^`�	i���:b"ct�;*iN֓�I	��8N��Lǀ������T�%������a�O�t�ܝ�8V�����6G��_���.����E�\��N�v��
ԨK~e����O4�5XΚ�u�e�m����c��\Y��{8W� ї�U%��;����q��HL�QfE�1���)�<;�+IG�|v)�tt�L2%(L�x�s<��w�'+G� ��/�V�z���}T�x�(ehZ��A�9��hƜ��˅�G���h����V��Tj�]��m�Ѡʩvܳ@�-��/u�~�Η�4I�59=��A�l�:K��_�1H	���0��ɜ�q�$I,h��H�.ٍ�	��RVA��-i&աU��:�w��U\s�%o]XJ�:���e��qK��|d��A��}�\MC�,m �{�l���O���LM��x-NtQoT�R�2���:o`M��IGx��U[w5�`��TΩX"��(�W�+�A7��m1h�A:L�P� ?����-T(����(� �Ƙ��8�&���!(7o��?9GıH��v�7Ǚ!��Z9��+��3Hj3��T.�b�3ʨ�!�;y�Ȩ��ᅁ���~��=�c%�`����R�8��3.���8����B�c'��� ��Ò��>b������R
�oz���5�W�����C�����#,u�2�Fk��rk�r��c�Ԇn���ԅ1�Έ�#�ōb�a����!:��#�L	�=1���ݺ9�����}�=���Fq���@������E$�3�G(V�0�ْ,�i��*U6� ��3�&]���-}"��>0���S2��Z�����6j�o��gs�C��}�L	�}�����'��o
T�>�ٺ�̷�bXI��r�������J�w����Gy��E�����qБ�B1�,���<�3ٜ�¥_J���5��skm��Td{�@�շ/]�S��yO/�WY3ޢ��-�Hǖ(��%���d����޶~k�>���F���6L��6�i� �i+��:�THs�Q�|����;č����7u�-�(�;�ϕ.j<����,��m�9�J{غ��+��bX�^(BƥD"{ x��@�Żn���wR�25�|�*���%��?,�J�Ps�;�c xK��= ݇ 5��^sˍNɭ�.p�}�r5g�.T�G� ����eZr�3W�١*�$����n��f��0Gs1q�Z�\&l�yb�ا]��������ywy��ho�,�� �r/ց갩�'�������l�.GzTc�B�\Կ̔"`N��=ʠ�ޮ�V���+��6���stB�Ey��Epٜ�5r �a洜,V#r������%xwS�y.͋"���3��i�Q8���RL>j�֠39�A�����e4�.���՚_�SJ�T��w��Șf�쉰ڄ9Ny6��@�[�S��NG�e���&9�H�?	�#]E�7�5Ϲ�=f�I��	�K�J�iK,ϗ�4����30۴ږ�1�m?�w4do�CT8n@ӳ!��cgB��P�q]�ǜ�C����N�G�b���Ke���E����'&J�÷N
n�`�ލ�u<�������GA�QfX�б�Sx��R��܂����hl�_��n&� �q�4I敾����&����qB2�ɯk>�0�c[�1?��̓�!�D�'�YH)^������<���o��l�%�����R5z�b�]֛���� x��%�;gn/�+����kQ	�}��M���&έUS�ǎ�}�3�qZ9���
�� ����Vw��\VͲx�)f�'�	 U�=���Nv�Lc��e=��)2y?@P�)gDЌ.'s���/�>�$RɎjvu�5��ܿc��@��pe��$į��mkvb1�tT
0��2RPT��XĹ���U\���U��?�����$��蚰�}I�	�Y�%���S�L'���Hu�RΩ��?E|������D�%��f�/��[���K�|����X����X���]�!�a��qKD�c��Ý�l��x����Mt��č�3�#����a+.j�Y�V�{�F�>i��;���\.����P�$hJ����u����O9��_|�F�q�J��H�Eғ sP�(te;/ڰ~���YU�';�_\ڎ-DZ��:��{M�*EZ�6� �o��]h|٤�C/��|YjdP�9�oJ����'*�kQ*���eL�x,ST<Q��?�D���KA� �W�v��;���F?fP}�����ACv��[i�N!S�lӈ��,~�6L{��s��]�� �ӷ�@��6�P�~�c��W2����"1��ٷ˄�vH;��͂� %'.u'�ע�zk�BJ�w>�����_ߝ#k�f�@�yc�9�.�Cv�!"8`���U�W���+`��P)ߧ�N_�*K��L��(�D��%�fֶ��@gkL��d��/��f�7�&���$��HÜ^��Ӫ��S�I��m��v�L�6��	�B��[]h�ĂW��VB,f|���&ү0wf���n�����f��$��G��a���4d�˼a�%��F&�5�kv���@@����r��|v�ȓ�G�
�3,��,h�vG���J�5��ݾ�6R_G�ױ!b��Q�C@0�s��[�������6?����2������u�z�aE/n��+ڏ��8q��;ew��Z�HJ�U�0K� �����
Ldv(K\�t�ˀ�e��*v�Y��j䑫�d��`�c��
��8��;~���c
X�����_�NK��1X��!�����<�k!�� ��0�~���c��L+	�B����@3�⟵g�䡴3j��@)��@�J���ÏҟH���6���02��j���,�����
n,˔���ϸ>����sc�0"ʦic�����k�c%�R�v=x&���e���C��r�������+8P�Dc��i��m^}jW3^�ϭ|5���l�b0�
�Ȝfc�䄒F��B�*�a�d�*���։�e���\��l�Z�d��?2�������{�)���<�&�4�����iB��@*�%�<��Mq�.
��y��bY���.��������Fu��~9��-��/cCJd2H����Q���rI��	R*4�z�`t7������4�3�����þ^��;b�Rwa�&��l)h4�cR��|���ѺX�I
�p��"w�����T�D��_\5#;2��)�}n�&Q��x�(�{�5��L~��Ȟoi�]'6�d�Yq#���b'���2ݥxv8�q^�й��ɀȏ��чi1�I���4����ݘ�n���À��^�pk���]t+f��"Y�L{�g���W�4�)+��&Mz����rd�RPW�J�R�HT��N�>��y�#�Z ���;h��c߽�^$А�Y�]z,8��L(�D��GKjN�N�b�/�x��`���;��.�k�ge��=�eѿ����ef�Ǔ���(9n���=Zѝ�'=����d�`���D��I�-&N3A��'*N��j�y�fA��m]z9�\L2����W]�)`�֓�f�^�a��*�r��l���T{�ui"X�W�q�����F��=�Q�(.?�d8�~Sh����a��
HsGDS3g��ч=�:|���n/S�_qh�x!	v���!W��@�C^������lz�D2=>�΁W�}�d�B���潘AeFqw5��-��:�A1�[iH�|�3b��t�ɏ���w��-�Qi�4��u5���D����t?<�$�Yyv���։v̈E-1�Gg��_��uM�E3�Zpl_��:x��{�D�!��X{5^�_�;G-mT���[��e�1^G�� �Y5ên��	��~�(��Q�U���+-��������qZ'�;x� ؊?�v���jx[8 �T|@Z��l�Z�<.a��5�s;U���Uk�7Z��S��=(����/t�>rΪ�z�Ѩ�)�ߐ�B�^�v����̫��Y6)�
^�7���U��1�	��E�;R �o�PHs���đ�E+��3H�B��t�4�<��㖖]q�ٖ��+C������������L��L�M��O��R��Zm-�����B ����Z����6=��Kby�z� �B��(󣲣�`���G������e��g�V�.3wAߞ�9{��������.s����=�]^g \Hqx$�i�z��#E=s��o$��DR��4�z��2���Mw�	܉EF0jyւd�-�7d�t|��M�ifR�@���&U� ^ؒFMQ��Ց���c�U@���j=/Ӯ����o�r@��1�rl����8�FJ�4FC2��5,<�%�`�y���{E�y/���z6Ե��x�sR7qY���Xk��'
�9ƿ;�S��x���n��)s\r�����\�� �;}�#��B�4�jӛZ�w4���|ɻķ��L-��/HZ8�`B��H����e�iQ�T�U��=��Z�:�8V�7�]a�ץS�y����D��K�\�=g'�ŽSJ�L�T5{U�~��f*��F֟� `��K�*/�̓�	E�<8'�U�C��P�|���Y��
�ȁ�y]��{�K��?'�=��)r�%��,�N�!BB��$�m��/+b{���,N2�6�2�6;���9�4S�j�QD~d$v�Jqʏlu��ٶ����^g\8���~��z���УR��͐jf�ӳ�,�V`T�,Wo���K�����\�\B0�*0_��]6@�s�����]��g	x]�_��J@0wp�w�D�Rؘ�\c��Xdc�~�D���h|�E�~1������l�l3�Hg����C.�����T�:4�U��Js0\6������-O6H� �ӫ�_{��b0���|l^�g��H�oW���J���eg��a'�A�tv�-�?�X�	nZ�^�����	u��9�JB�=7�?�-B�jr�L�M0pE:�[���%�@��@���y�3_W!������	��Sb˂�CwZ�
s�wP�Or�Ao�n�G���q=�G���}��)��
7�)���MX8r��o(dL�O36~AAr��g��Q.&Ԅ7ОN�v�hmX �@F��ѱ�Q1�]����u�^�W���w��f�K�vs(vL�=�J-�9�o�E�6��fo������/nӐ�Ȇކ�j�G��Rvnڬ-�biH��R�ڽ�*���� �S`ow`k�Ғ+�}�s�L��,��t���Г�=�8d<F�$�zp��~?�����߳���*��̕�l.�K|"b�u�W4b��5�t��rf_���5� %�^mP �� �$5�&�.��RvҤ0�cD���2`�=�dq�,�[�c2-
��'t��4,�8� Nq��c�[_��X�,� *�!AI��<�eo �0#�Hve���'¬�9\��s�6�����0[��=��CB�;W�m9'N��AUm=x"����H�nm����ړ���M��
Q���9u��h�S�Z�?�5�onY�_3�˝B9{��6�̭Z������7�E ����ф��=����g�AB������[a�3�F����1<�\��A��8V�0WEn����k�|7A1a�	o/
.�^�0�Y]`$)�P.��l�Gu���b*z��?�O�	�`\Ŵ�T�����z�B)&�hh�}��z&�e�e���;t���Gh���"[N殫����P�'�M���ߧ=�N��9��<ul�+#S��y˷� �*������9[˸!�y!]�5ra��MA1�V������W��Ŏ�����>����V%Q�m�ů9`��Oq#&��S�IdC��LBe«����]�5T9Ȳ����s?��wE�������?- 
�CB~��Ch���Q��i�R%_�V� ��l�V�f �h���ѽ��z�\�3�C쭇���I{����%�m
��A� �*�#&��7�� Kc��\�+����q��� �mc��J�;U~[z�좓�X*�eT���t$����!�/�ښV���p�4Р)�K���T5�Y���=eo����y���)�^w��,�j�%�,q2����%���V�|]R�nkr�p\Dem ���PI#�����g.��^������_���iG�t�����Y ���ģ_�1nJ�	y�{~g��4����<^{�	 �-�$�:K7������OXά(�(�R�x��+��/%>+��XvK����Х�N>#�,0����[G�d�L��c��@p���MR4�	���)�>��s;�ju�uu�r+��!�$z����lB�K|�R�2;���?GS�q�Xh��"��c{$ހ�H�UI)��A��,J��ӪU�\q����Pu�ߝ��Ǟ.@�Bҵ��ҀHG��!0$��&��`��u#�/��l�P���6�� e
���':^��$��K�:=p~&�F�.G_�+�pB�3�;�u���n���A�׷?,���4(<�S�yM��(�JYa�y2󦞋�8��Vxm >�/-:]��_D����퍿e�[wpю6���W�����Z��h,'���U��FF�u/� \��D�# �E#�RJk6���<6�s�1 '-�0�L�_&+ 9p�,�x��^u~p?ƭ�M��S�_z���ͮFx�'T܏���B�TU�<!w	p4̳�@|��a�N=c`����T ��:c?�^��,�(�9 �@ך,��-�|/Zx��N���G�:��=��~፥"Q����.��\	���<w̈�ؼz�?3��3��11��vgx�{�]un�x;�_U�}��J�֯�����(k�p|Gc�>	��;
WӋmB�Ӵ4=O�2��o�m���y�W�V��Qԥ2'Y������'O�5,Ԕ���jlIb��O����?k�X)���
��.�vL�?	�uJ$�����W�Њ�f��7�E�I_����������ٞ^2t16wA{������}����4 ��&��ni����TP��.�8���)o
��$�3�1 *T��A�z��H1�MH� �_�����S\��U��I�t�3楆��]��¤uPp|�GY�~ZI҂�P��.ͻC_�@������ZT�����1FY^^s���Hy;�����S,;K���3��*��M;W&��ݜz �T*Ţ��c萉�Q�g�Ԙ݋>nŕ���Ý���"������e��ϊ�AK���� ����İ�������\I�����ټ�b���s��Y���\7n����s�Q��N����b���鍉�O(�Z�#8���&�f��x�U�&F�WݕYJ�u�I#�UX�V������ļ.�P�rC@����);a ��=�K���nM	H��^����܏�b�D'�r��}����%�%1'��A����$k�S����R}�������%ZL��ߖ�|dU޲BSS�Enњ���
��8vxa�C)�h�F���ؤ���u��n���8�d�ӟ��j��46~7���������
D���)y��N'�A�A��/9*?��W�#�˸�L)5�x)8!w!�mOV��ģ/2��#�33i�����4����2H���",��x�HVq
�8?µ�Ř���f�8�AU���\���v5O���s�4�hG����9K8 {d�|��Χ�5�	����&�<�|���m���g |o#$K�)c�p��gFF�H�#qMOj���Q��� �H�Xz��u�"��D�Y�v����y�؍�g�Q�MȊ�����\�r�Ѝz�����<��֡xۣ)��;�O�v�Y��Kh)��ȫm�vx�0������F2[aRZ�l���꺜����}/��x���Y�@v���\�Y%�3 Fn`�N�[����H^a眐z"�^���DyK�85�C X�*{�q��Q�z�g���$�?]��Kd~���r����=[pFz�n��]`������=����K�p��y�H����ٿ;������Y7�B������j��\q4+�v.Z|�3
����?��69�K;)K�G��}�B	:��)j�;G�@�|1,��F���u3ꉝ��>���)�{B�:��ܹX��0�)��d`ԑ����P-�"�?Bcz=�s�f>~h����%�����B��cڅ�P��W�%��φ�X�!�N!�<��<�N�TD�!Gm�P���L�] �����k�F���7�s��u�hc+��Af��%/1ݗ���@**���_П��Z��Pڏ",��	 �<p )�ތ�YL9N�>�������Z>-���������w`n����2�sm�-6/k;��C&�5�d�/�{mݐ��M=�ҧ+0�`c��Z~�#�~�Q�����&��o�z��RҮs����]EK����kGx"��x��k��'�e��=#�G��� ���2x���Q��αf�^K�L;t�K���+q�Pc��2�K�#��1�CL��t9~��W���n$����c�<�I?>�. h�^'%�|�/�"LܣH& _I�����U�La�ɧ�����y�ÉlUĞ��(�������kdpn)T�7�uZ��¡|������w9����\G��ZOx�h��6Gr���,��t�J숧�����V/����3d� �����ܕ���T�{'��,8��8s��@�Hx03d8���tM�ҚB�E�R��J��w��q���))J�9e���E��Z�f���<���ʵcpU���7@w�������E��aQ2���#	�0�㩡�2)�)w���忙I�pX�~륞�b9�s}gD}X}0���x���s�>Y9W�K�������kf�io�^n���n�r�/#�4<񿅌�w��\M��Ԙ�		�M8	�̂{����h����nǥ���xyԗ�.�����lP%B��tf�J��촢�؞W�NB�Pzjp(;�N����A���M�������%Hʕʬ�F3а�M>��B1ȵ���������e'^�M;H� ������Qo#i��U�GƄ���tәjq�p��`/��^��(x[n ���ͩ��0��}��k��jI}�%W�oSy`����2���9�4�Fg;�^���Z@�
an{�k�=��g����A���.�Y��H�o�%`L���Ţ�x�������U�W�2�p���u��K{��}��j�ta�����48z���������W��u,�]�7F��D�x�$�jG�A3�����A����9���mtI���>�ϣ�l��=ȭq�Q���O�&�_�O\��w�;0���b�r��/`�ɸ�f���45�wLe#�%��:��f����7e��g�1]���o��	��R2W���b�h����C�,�:��oC��j'�<�w�?7�Ck��`���^�s�:���6}�˫�y,��mz��:����$!�\I)�b]`C,�H�5y�V����D�Ǽ��x@h�D~�R��KR����ĸ����5C0��o&vp�!h�[�bk�VD��l㭣$���;S1^�6l"��Eyh:�jro�����!v�T[���x�+>�4�e�P.wP�$z����ނ���Ƽ�R�ӱ�p��@[i�� vC�K� /�>�ޞHj]��P�(y�~s�B��GkCg1�l}"O&�S�7��Q���߯�-��
�S�~�gX?�c�T�ne'{�,)�\�O>%�t�t<I�m���W��C`�?^��k��Lb*;����׏����\�#����h�c�9���\��-����6�3����'�/t�.�� _t�Y;�o;xL����#*���|.(~_�U05���$2�M�r���D;�Hln5���d�/{��Bӌ�GT͛ 7���XG��� z	�����A�OJfv�$�Ir.�`���[�R`���r��wmfu��=NU�$��$�*��}ve��b]T�����∳��u�/5ȋ�� �q��ɩ����\"BBЎ���R.+�!����k�@*�)�Y�<�_�9�2	?���U ��6��|5�p?l�7O+�<�� �E{���Ȑ.�ظ�^j���@-h�ܤ��r	��D�TȘ�.A�UgBi��GE^?���k��|�!:�ʀ��X}p���l+�ӿ�|�%�kU��/s�����	`��Gq����fNY��Fs����J��Oݾ�Y<L�����4����d�a�C"ￆ W�ġ
>*�X��/������H�98�7ˀ0���H1���{���=ŻFuW���u ��I�j ����ӏ]�y;���_@g��98ö�^�2���R�� ����ì�v�GޭQH�*{l��i��d�"�}�+x�	�@�Ri�:��n؉O�s��m^���?�P����޵�7�!�bfT+��69�u�Б֓�~�\&(Z'k}`�x��D���w��5��3��$:M�w�T�t�)���p��R����,f���h\�wZu�2�U"��7mV�D�|�	B�si��m�[�o�s�=���CK"� I�HRRxN9���~B�(����o�G��_k�A{Y�v�$
Ja�HG�?���G# ����u A����50]}�p4y���Hж<��\b�"<B�|���)^�����h�@�.`K�]��U,�rQ���vI��."�&��N���$�RC�X�!@����ah�*��e���ۭ� ���oM���JH�0SE�I�y-_{�O_ �)�+�����٠�)E[^P ��g	�g�e�D�����f<6����p���ֵ5�E� ��dY��B�h.�@�";A���A���7�������+9��(D��\��Թ< jA�[��Р�D�"a� ��44Ϋ`:Q�羱��0{w�|e������mB�����p��w��n-N�U���Kbگ���U&L5��s�;��ڮ���� Q�G<����Z3�X�\�bt�8�Q�.��A4��up�L���~
��m)���}Ш�ш^���P��D>/�B�g�8�����?3�F�`�+e��0u�آ����h�0�iz��Y�L(���Զ����T�.]�o�
���!�גX�����0�Pmk$�����v�j}����tr(>�E�����$k'I�a-�|R���ae{�&�4NZ���Ld}���g㬞xB�K�|v�9��&]��puwO�%��10���G1.�/���\Xv-�a�w�{�����*x�A��������+��;��1yAs�bC]�CBh�Y6 b3�p�S�M��������IZ<��}%��� 	y,����~��o��RU�R���qܴ�Zd��k.�*Y�T����Q�9���g5�P�n��{א�̑�.W�^�����wm�69j�G"	�$��1�L\jf�Gbs#Z�ц�:Ǝ�(	t��G�ZYl����nV��d�#��ǔ�����RqZz���p�������]��W��`]eL�e8��5�D�����H�w2���Q� mSq�'�G7MZ.�)�6#� [ܓ\s�Y�5���&Ҟ&l��?�/W���Dm��_���U�Im7Iܠ�[圜�N�k���\�g� P/b����<�K{}g9P�2�s�$���,b2Zך��])�݁�R.u��Զ�Cj�U6����K]�s���t�3�{�Y����f�6*8a(ũ8�gzZcSɦz=
Pq"����E>�l��!ش�0�(��gӆ�"J��w@/���]�Kb��>���v�F'���(��_�>�G<�r�꥖5�}�J�(�h2�@#��"�uax�`p���Ӽ~��4�r��}�P�"�3:��t��@.�g5A���Iא�_���nZb�-,�.��\o���O��~#�����O�I>n����{ r�zU�z���yeӮ�&-��E}���'~W��#�_Qa�Q�c�-Y�m2���Y�j~�R�;�T�n핏���N�{^���Q�Z�9^-`�i��ᙔv^/h��՛"��U�3*W)ջ�򸛡=9~�~��I���:$��34���IT�۹M,P����dz���hx��qEM_���بw��F�@��A]kԠwy�ӛ]���OF��q������$yڬ}�����!I����ō�2U��Ǵ��o�<�D��*�b��b󱏥-v����3��,Z��P�sPF
���e]"T�u'��䦓�=r�����eק�R ��#��@�~�N0��+�w�4�[�eL4����
]z�~����P�_��Q#��T
��N�o��SH��2�X��ᇎ�4��+Q9�����p$J���_Z)�yj@O!�Ne����\{vh*�aÂB�Gƶf��*�W�1ŏ��|4r�� !�#0�-g��mS�,�����
i����z��t?�6��2	醃9L^�H�k�a�n�=��L>������]ܨ��Eg�[׫��C��x[��E��ԮL�
�~��;&�be
���k����y+��X&�l�T�ԅ8-�rڠ#9�;���L�����9�,�4/�;�~�?VH>;����w��`�3���Gjm)\��DV�5bڗծV;�z��������V�CҺY�W�ߨk�nL�K34��x���1� Cl3*;�:�����U��~4C�d���2v`��6�r$�H~�y��}ow�'5�5�ɞ���0��;����f��d|�"a�����οp6o�C.#Ǟ0r�U&�3���J$
�?x��w\���hE�W-`�x�ǀ���,5��Kl?9�y���-�QM�����ݪ��ɦ��y�;ޠ�uD���7�Zh�@:�3�z�^V��w�M����*���}�`�E�&�D�P���p���m̐aQ����>,�x��->���o�Q
�: `�̡8ɴ"�Wf�7f��1�����լ��)#��i1��C5Ls�u7���"`�_��u�^�N8��
��0��H2eZ݂|P��i$'���k�*�v^~GC~���#�uLL$u���!*��_-�ۭe��a觇��`���@-���l���$�@@��K�P �6�4��;�X���;Q�TՠiȎ�m[W �qQ���
3��]	����5q�1=��xF��xd�ֱCw�R�J��3�H	��dNB=�O �'�9~�.��p�o(-;�\�C�̮�b�~�ܠ��|�L��#�pϔ�,�I|����,�]Uh�Si`����1C�En�я�<��ٮ?:=a[�m0�ַ��M�rMd����EW�f��g4�j�ED��iI���x�uwAx�2&>����OiwZ�~��i�ȥ�ʨ7,� �F�ifp���vX�D�쵋�[>\[���L�i�U��.4�2?�Gg�H�`\����������-��4�Q�;bZc�^?+�0S)��Z��~V�ڋ�.-s��3�m����8Y�J�At�g����� �O�mh�G�^��$�������&0���v�gf��uf��bv�(��K�vo�����IWV��Pk}-���2�ӹ/teNL�.�R(�<��R��_�j(�mSt[�D�A�+Ts�J���BJ��樂eA�̟��L�M��ϳ���㯓Tʊ�3UG
�꽱d½�wG��g����{+0`n�$A��j]J���:@C�f�t�֩.c���r�Jm�kt�"�A���Kָ��F�奻8O��'�n����$O:d�Z�Ѻ0�� p|�Yl6FK�*n�NCo���Z2H�YT�#9Er�b�W�:����$���Gs��q[^9��>��͝�6DP3�),R���xE�;��f�0m��·��a�ѡ���S��ЍH</��S`x �C1�塽�F�/*�v>���e���s�Q�kz���6By��] � �ˮ��O����h����t�ÀiG%+�A֮��?F�@�漌I����ñyn�-��� �Q`K��g�Q{�*��	r���Q��~R�b�����PJ�fx�L���id�u;�Vڇ�򍤟�f���J��8 k�dJWZ�4�f�4v��j">өJ4FK]�7�S��)���H�_m=����$u�y�g��f�6�I��¼O�>��=Ʒ}�>�xxw��:_��(�$ɬ#�q+ܘ�b�³��<�����U� ;�Q�*�gA���\�I�M\(X��w
�t֥pb�H`䫎Q�Ȥ��������j�"��V� �}�����o�B�'�b��a�3��-z� 2�y�鐁�輔-����w��X}�����(�2z��j�l�1s\}���j.��.Q୑��5�s����P�1���	�С�CQ��ʎ�=D�*���ڊ���[��몒��M��HI̧r^��q1�he�S��,H�'+�q���P�>GUځ�{�aZq{'��˳��-YO ���o��.�;7�U)#RC�Ó��pZy}����ϻ�,p���"q�C,���4��O��u�����3J_F7e�].������/D�sm<��,N���9����q��;��ZH|��<�ytҾ��ʣګ�~�9�d��mI��j�8C��ϞZް}���L��	��>���-�=8=��:���b��#)C�#~zx��u�UD���/��N��X��/�Q��k�M��7��y�?pd5�׏Y�	 ���N����B�\lLO�N�w2���`w��T,&���@Hۓ���=`���A����1�-*Zk�}*��C��a-q�m�>�`ޕ���ؕJ�w۟��P����Ő��#ԃ�)M�ym�RaJ*^k	�����Y��0����/��-�� +��lE�)F��|{�Ao�E���*�ԙ*|^���,ct��(��40��;�_����|�Vے{K0D4�<��p��me�����Z�-U�����E�r���<� e�� v�5|׸�c�r��H�xd�X���<�*4�h$��1l	#G1�JU=OTX��11#��#BOX�)u�[-m��(�g��l8�t�S�\qx@{Lg�bt�$���=�L�ԮE-��$j��	o��o���}����ݺ��	F8�����e zkJr`R-��h�PZ� 8��S �p���`t»��˜��	��=d_�ܣ4t����&�aڧJO׷O�ᐫ	�*��1��K�����	a�d��N��fA�����Z0��������餻���hXSsU�>���/���@)�'�W>!V<�u��eݠUi�j���ݭxX$����nO0��s{��<�cս8���$p�exL�l�1�u���{Y���1��
�$Rz0)�H˫L~�J]�H��V�Ba4v!���	멒��ֱ�c�*� �!������Q���[�'��Q2�v��En,�z�xI�a�E�HO=�/o��������`X�І%��f8?�d��z�R��>� $��9)�(��q����O9�}r�s�Y��ԛ���
��.,�B�>����ᑍ�Ѧ�KZD��v;��,���f���o2J8�������(ϑ��QHw�r@�7�v+��ʵ�c����N�5g���r��*�]1�>�J�_}.���9r��3��VFؕ����=��(%��'�����dE�1+�"*�����Ѯ�T����]���c�I@�,ռ�їm�u��=<��!j,��(���	��Q���+�. {���DYn�tH^��n���� H��K;F�	�QJ��^�+�9@Ş�o4#�]8`W��sd�x�^ ���@���.����g�S�Ow��N�A^�1p��=.����l	��s{�z(��nΒ�0> xs�.������'g����ǚ�|3_e`���-�'dT�E~b����<�tu���/���e"0CU%a*/[%��J���9�^�(Y��̴�X�Z��}^ͫڨ��4D�:��%�?߆,�Ċ���_"�HR�gM����;�{�0�,�!A{�҄�$Z)�+z%��g�A�<��j���aT�7}�LQ���㈹�ߔ��z�q�Y,���Jdon�(?���汤��@�l����_}��)V�m!�z�Im��A�0_����x ����$��>E�4�"�[ev��W�#�x�P'�oّut�A=�\0{��@�/-��T�1���Ƥ����U�*��\ij�p���Q�	@2���)�y<��Be�b\P�4���Mn���
��	H���|rD4ʆ�jyU7K�d�w]�U����	˒��B���� �<�U��%�j.@[pN�&�AC� �����/nn�YU2���=����h/�D�5W"��kʱ��+��?�H�,�o!���@h�R��AhkR���m����-����mD�KЁz�.L��XMO�	W��;"����YǨ/iE���Otkqo�"�T�[��1�]�	��)cځ�/�6����?(~�T��� ec��B�'AfY7�� ��!!\��[�p��D#)i=~a�?_�H�>�@i���&�;i�v�ίGP0���:����]x@���y����Ug�ͪ��Ii7P+ÍH�Z��k��-S:ke����WOR;���M%k�odlG�Y�FS��v���(��
k1%� Uڸ�A�S.�SrjNc�_��O�;lq^Źgc������-js���PN�N����xL4.JJ�����2�0���|�1X�>�l�w�\��W_V��6HH�z�1 Ls�xG�ֲ��T�W�8�&���=lT��_��N�ǰr�\�$��vqN��> \�����cUBb���ϥ���Ԧf�BU��u j% K�ɍ��HF2�`&L���g�5J�̫�[�\�sC�� ���84��|��τm\�O0�S�yY��龎o�؛B��0��L$�$p��X�h�$Z����|��*pAB��z�z"��1�ݩ���P�u>����H*�ౌ�w�3#[ I�K��G�^�����SY.�(�ԗ;�B�53��-�Rd��c9����<ׅ�T�&
�QF�*������#��u�0�C>���QD�;37 ��ۖo"�������r�27
��q0i����X�$65��'�D��a��x�̐��iy�E}�F0;�a���bPC�ַ+t��	�&�wP%��U��m�G�E��ꇊ�qR-�h� &+�x?x_x�ȥY�O���H��	�녊:�$��|Ԅ�����m��r�܌�`�z�
�[�[TBܙ���@��3l��G����j�����eB6���x��m�eGr�e �l۰��5���A.m�ե�F9����` O������"�Ӑ/�1�./��t��O#�^�~�M�m���SW<��i��-?{�W6�+��?w���q��
�˓J��>�2�N�ts�0^+n�tç	���ȯ��{��5pgc�Wk8׷ �O)k���x�S���|,M��:��W��EȐ�S������w;�����l�rM�!��bP�+{����@�����v��t8
�_�4kr���-W�!�au�&�R��I�~M�rtp������>E�X���;,ֵ��\0�)�t?��T��NQX\�ڧA�H�c\4�������p��nH5j����7?�TKUz7��5�:�2f--/��O�� �\b9y��[�T��IB�=-`���f�)1Q�+�F���Q0�p��F�/fl&���F�G�ga0Q��\g)#����;21�閶��	{�e����������mp����"��(�����Zy���q�>�7�>�}��BZ��"q�	S��iclZi�t.�o$� ��ov:7u��y����/��)_>޽IKµ�I4G[���j��}M>�C�^��<DJ�g[�R���}���s����O��̹u�����#��U�+�ڜ��Ө!�Z��Q0%�/�c$`Z���O���1p&x�%~2�(U�47 e�щ2�mul�(�ϲt��V�J���[�~V��s��X\f+5����p��4�r7.?7�J ҉.>E;|��RP�u�n�ń3_�<��2Z��f#i�AV�Ƙ��AX�`�q��Y;w;`�vދ��Z1�����Oћn��+U�8�j��j��?�<��5�#�����*��"�`W���vr:��fP��mS*��FQX�$G���_��w-4y6Y?�PW$��ـ�a����?�T���v�=41+[폰"x!���[�y����C�JXuO^4��ɚ����v��Ⱦ�~cSL-кku�<dh#�����r����I���  e[�n�"Y+���ă�
����@I�A'E���6�;w"4=��@K	6 X)�Y%6rk�0.�
�10#�h�=�I$i-�&/�.���/���~_Z��Uo�� �`�U�#���5�v[{�7�6�v����&�ɦ������b�t9�.Q��Y�WI����!�W� �Ab3��p��`N7�%}=��	*�^9�;�D�� ������j/,'m/��ߜ�Lw�V��XJ]�I��e�ɊQ-XS(hFƈ"^��gF�hP��so� ���#P+�Gi���ˣJ@Zp?��-Y�B�I�͵�D�' bl(��mמ�k}n'w_ǯ�t�?�Q>�}�V�h�t�V"��Yw��sZ���'Ո� 2r<hD��F�*�hZ1�M�=�2�=�F�c|�~`��f�[�ʮݹ��N�2Q*�O^�2�%�P٨L���h�j�_J�@�FH+��?"m
zvax���=�?	J�P*H㞔ق����I
37���h�w�tLv�a�VN.1��;�b����}w����U*���u�l�S�����\��[�~�/Mt��!�|S�
�������N7��}�����u�_��]��5���V��æ��;�y]I����kVM�6���ʭ۔_;:���e!�`A�2�K��͎)�Vn�Y`���]�=r�mnv�o�N	��q��?��#;h��6}\�uƐz��z����[�3.{�<woC3΄H{���z�Ť��F7�򸈜*��	uڮ�5��#����DH~4?,���q:�*"�%�_�L�3-nGM���|�+`�\E֍	���2���G��ut�t�7A1�J'��v�e�L��� �x�Q�|ь+
� qM�NT��}0���,�}�~"����xR&�t�E�	�v�i�,�H�~+]��K�3c_>�Rɾ�j@�R���B�0n�� }* Eq�X�?�
Hv}PI�ҊCbC�����9o�v��j߇�Y�/rM���ױc��F8��5 �Y�	�>^��)p	[�GI�Gd�M�s.��z�P�dht��wIz7-�ɠ?_�|}�ts|\�����[C�*�AD���� ���|�I"A#�}ʜ����S���
�P:Y7 ��W����t��<�KN�t+ǂ!/�'Y=���)��p�&�w�k��F� �]��������P��o� �[��3@'5V�E�����[9]�s�f�cP=�4���ޚ�K�I�ݻ)�N���7��wK��W�zE��a��J�]ȵ��Y?����L����U��"�u�,%0��-W/;��[~��Vm2����,ð��y6������T�$��>��r���kM7n���q'{�w�i�W8.�w��-~易�,�L��?���X���F϶Q۴��
u�t�ޓD��d��xBǴa�Cp��ϱK}���e�eg����'�t^t͘�7i�v^�6���k����@��ۃ���PY�J3椕�]���~$�{��	
:�`1���y������`��j��"�XG��[7�@�������
��v��5�C'�k�`j���M�٢��<K����]8mՕc6XhE���S&�`x�,t�@O��'v$�6��#)��}��t���U�e���{Eئ����.]�W�堎4�3	@]��ȯ�����3�"��{|�zw#Φ���2�[^��y��O�;S�1�.��zfJ�[�����(�y�{�d���X��y�"��B=�_�eY)�H�l=is&n<+p���a��j�}�n�� �g��r�ǦG��w
F�*�l�yX���E6<� �7n�ȫ����w^� -cc�##�O�T��[ʃ��
�X�b��F�cՔ�U���UN1����,_e���5��4�gr�l3�6<Ű���mޯ�̬̍�F�U�C3�g�܁�K7���n}�o�!$�=層�Y� �J�.��	A�R���|�k���;�Eee�LN�5}u�פ�����'�F�N|�%u���a����τQ�IϺ!����v8E��z�v'@2]u���w��@Ù_���%�㞥��U�!yTP9is���@��2�KŶ�n�FA��t��Dݮ1�cj~����g�ǿ�d��t����y!��m"��rN�e"@�;�/�#}��S�X97�	����5��"`aC ���t``��P��@�:JA�N7��>J�1����RA�Cj����R�w/_~&	�C)�p��IC�\~���e��M���Z�z+�[J�O���"��m^�ĵG&MP��S�=w��O	�R�3�p}�Y������~'�k_�!��v���K��0����&�WL�5��D�n��Ya.�����q$�2�eI6�O��Q7�!{�`�ݶo&�;qP0MB/�ڜMN��N�<��s��Y!K�4�{~rM���dXS�bt���ۄ�8�1]�UF;{��Z'��(Jl
],��,4���	�}��F:�i{������r$���xU�^Vb���+��x�1��l�~a/���Wl����*��{�����:���;�?)�r�6�e:N��ꏔ@c*��blY*L���m�2��5x\�I��݈�0�M���X*�6U�<a��ᦍ耐 v#�&�!��X�o �Ӱ.��7A�l��Ǫ9�hO���dȸ�^�;C�z��eO^�-Z�l�%���|�^���k�4|�s|IĆ�Z6i��ohĒ���9�k#�(�oo˪���"���I��Vڹ�}C��}�M��qle�ζ_�Z�@�G�6����H�Z�.U8Q�[��D�v��<L>~R�#a��a��Yn��p�/8Ғ^��>~ݕ�%!z/�]�6g���s��dAV�������V�H�#,N��Ŕ���y���k�狉��B�u��դ�>k|S�.�[C-fnG=
iq\�D1��yKI%�(<	��Q�k6S�і	{,�D6���љ b�ɝA3�F(\ooz� ��dL'���b�Uz���GOˊDD�o��~[�z����T"��)%d�֧��wC9����j6?�����V��we8��P�*lc�:�5	ZTu�;����7i�ͦ��I,?��T��C�G�v�Hн8O��5 qT>�M�MJ�#R�dQ�e�P�+�^�&t\�^'�q�/K�'��k��#���9�S���@�FDo忂�(��ŕ�=:/F�l���4�E�s=91�ݝtG��-�'�d���8A�Ku���
�c���N��B�eA0﬽��ǁP����W���^WF,��e��t;�!�%�7Gb^��A5L������TM����ݘ�^�Sj��S���疱�{�N�]��I:h��$5�y9���H����C?u�;�ք��$�Ó� �p�9���"X)�����Č�x�M���gQt�7�<qh��,�r9��@�NP���{�����x�����x>.¨jEi/~�y�������o(b)p�h�:��.b̧c�(\ң�YOQ��nl�nO�_�b�m��妲<��ոN};�����=h�j��� ���D��m��:���pDn1�@���Al*�Q�e�2z%ԭg�� G��3�`	29�(�2�N�<2��K8͌]$ל
;X[ݚ͂AI�!b�8������f��BI���[u����R|�ZfU��E=��>�n��r�u��g
�*c:V��i9-����ǯMF?��8�}f��3���p)Z"⣟��s��,6AD�I�/1ܥ��;��1�&��UM$d8[��������wP]=�aK�т��[�ln�[�ӛ���U/K(���� �i�E-%YL���������4k����aǐ�b�l�K��
�Q�^�PÎ���O4b�CJQQ�qPt{X��pxr \��j������������1�߁Y4x
*�!�]?a�A*�H-�z�f�< ��.v�r��p��E�����> |>���ECh��{�Y��f�1Z�C#tB�2:�����ZP���|�=L� �_9��yF�TٵFwfР�
���7nX
�/����e�Z�,��XB��<\g��IBs��8��-��Ҵ�n�E��;��0	��E�"�D/밗|i�O�M�J9�ez������S��IT�MU�*I�9	�2t�J�0�f¼B�L��Cf�[�2hv�n�yԒl0M_�xZM1;z��7|���L�i����Z�=��i�w��]��Ռ��w��VBL��c��c4��D�9]<�u�L���-� ��Lml��e�_�*��B�,�����������i�[?��bsGlJ�=ϔּ@��i}�������Z�̾�1��ų=�fˍ#��їY��
:r�����mIZ�3�s�xM4o�_�7㭄R �ॅ�(� �Yt����ZF����O�{�b�m��]����8?1����.�6vrff���-WO��T��Y�0�+�����5���u6�c:�<��B��� _�D� �`��kG6 �"^�_����2����Y�0�W�>4����q��`���[�v#F��]2k��0�&��MU���=�y��Mu�~��1w�j�!:���e�E��(Զ~-�C�J��h�PUWpb.ܶ�k���=�>՛�%�����QM1tB�ۮ�p|�:B(�5�nf��n�q�S��`3���-��u�Ow�?�0;��&�q��Z<,\��Ĥ�r���˴��N�.�T+?`� v]sݺ��y�h �����\�s�$%�s��@"�,e|�D�+�Wfs�j���ť93�W5����/�k&�X��K�x��а�᳻O��x$>��)!+�KeF�5T���"�.8����s: +�~!gN��:�ԋ��m��$�a��N��J;�<=H~-N�&�]+�����?.�T�l~�MTt������M��b�E����S�q�d{�����'�^��L���~������2��xVg��Q�c����x#���1��4�W��8\b'��<V6��U!v�Nht��@M�+��粟��z�E��>��ՙqBò�Kp���*#
�}��x�{�VU|�KVSkE�ɧ�A����&��Qw���-�Ft+�Pw\�^m��&��"%��_ufI�AE.*� �8)�ѺFV�k��7h.�Z�.�q�`���ufif{�g1_�7�u���)/0����Z�-$A�2yyNe�'S�S!Ż9�Uy�qZ��˅�5��qߗ���a͂n	oZ�~�xj>Pk�����Z����q	l)V�m�ր�_ ��m\"CK^FX�'��F�r�	�혊}�Ɗf�أ㓓��l�E h��m6_��w�?���!���Z@�����^d9��i�큹��^�98D`(x��ġ��M��QC����sm�Z�U���L��/��4/g��T3G�گy.?�%�u�y�_ݒܵ>r�*�wֶE!��xt��a@���F���[������&|g,�����u�}:ء��@̺^�A#OA��!r5��g�O�3^G��R�tX�EC@����3�UF�M�F5Y��R�$W�������Ka���'[�Ta9q.�/lA�O���%�л��H5�^�!����b�O�ȩ�S<���	��Lh�҂����_��i�V�o��S T5<$fʾ���3��p*�į5S4#����ӋCP�ti_0��a��{P0�>�'������c� �|�d�x����miG�M�֜&9��6��N��5���q_]�x��3��>[T9�2:M��B�X�v�'>fĵ�[�s!]���	�R�$�b�1��j�|긒<�m%��ɲ{�ޫ !Q�X����q��M �k�b�$��RUa����v���|�Y_���cj:6���4/V̭���G�ٹ�>��%��>�`W>�U�V�Ġ�"K[@���q�R"T�"r��r�vy�YL�Մ����3�y���{?�n&���?ƃ��&�\���t4�r��� �s���n�4bj�-@�*���ד�+Yz�thc���j[~@L�
ڙ}	_��"偨�l���oV�kc�֣�AW�H�R�0,���ئ�P)�M�.���f���2$
z�+�0En��F%:�Ik�G-&� �E�� �ƣ����i�B=���GU��a���R�IQȜ۲��uV:���3"����fx{����k�W�+E{��7��|�]~����*=���	~&�޽w�q$rM2o�SqQ.��>��k@Ű�Ol%��u졂����E�m�X��N�]�ٌt4#!�����K]��*�-��`<_kZ�+\֪:�^��	
dc�vTf#�|?^�׳�ټ�L�|�>��;����4aƴ�PG�@����;����V9�}�Jj��v�~7s9>`�u0/w"ʬ�N>�L�v���m����ƿ��'��{�сu=�{���~��n"�E3�Ǵ��\Ӎ�d�v���~KGt'��<�>��"�|!�(�q�~��$��6��qi� >$a�f��wT`B��KɎQu82U���Nr�gձV�Um\�2�D�K_�>��K�hÇF)�������wW�s瘨�[^u�ԙq��4����E��E0�p���{���6H�	�6�B��e-�ѓ�A�X��P�*zx����仙!\�������u�Z�fX����|��<~H�cc~�UV���X�<��is����aw�d	�3f9��rq�sg��z�>��&�)���BzsSCɋ(�d�M�ɝ/��E)�M٤��|�(�=!>xg�(�:ܫ�3.� �� 
��y���S��E�JrS���7l�m�rп����6�Ү/i�ҥH0�J= Fi4;�jK	��n~��c�J\qq�E��H�����!� eX�&Z��7g��3�2!� �؃"ST�0�I`R�7�Lo�3�E$�hդ�F�`���y��cVAo�	V�X������� �i�qksw��6nIB�p��\3P����Eh��c��R���b�H,��VT���|׈�)w7V�X)1>�OP�DY5���� lT9�/KZ�ئ�ud�.fR3g�L���^��=,Pѹ�T�O.lF���i�N�֐�gòɇS|�����DR51@�G�B��
�=z2T=�
�tr�G
Z�@�%]X̐��H���amv+�:x���YF�K�(r,�-9Ћ��:˃����0I�� �?�m�TTm�$?���P���c���dD��6n$�}[î�31~Tk3
��o��aҏ���$�B�����Xs���P��Y\�ۚgط�P~�0@�� �iY��+�(�e��t>�c5��M"S�׆�2dE@qK
��r>:K�Ȯ}(Ӂ�A����qA*�/����c]OgZS����8��Z)��f��`��2�;�+u�#������*^���g����_귮�u 2�6`n��l&���zh����VX�d$s�)�I�o>���q"6�!���9�9�q����l�Ԏ�D\C솯��[��W���ˍ�rIT�<��}<�ڝ��x�v�$.=�1?)_�'� ��='������l�7g�J8��
/i�̧F����ob
����p�2ň��gS~ݶf�ܙ1�RƊjvᦆ��G��_�h5	L<�f>���'L&�ۥ�B�j!�z_��L�-I%��k�G�<�u�6�e��ӱqO6���R���o)�X��h�W���F��1�h�=Fx!���c�@��Xd	��Q�M	0���Q��w-���G���҄�`Pd�sSAXM5�C��\�R�w�Z2�Y��6$�����1|l�?�\�+2��s��ΤʋN��t���C�ot�����&]6j���(�l��,}��Z�AB���acc���n\j�c��v�)o���Xr���œ%t�2��T��à�l�_|.V�y�V��i�S�Ђ�/��gjyh#sz��;�x����ƙ��WH�⠧Wy�Qg&��k�U�0��4��U���r��ʈ��Z��h�a]����hI��Rߝ���T<����-��+�y�Y���0��j��Y{�H�Wk��E��L�W!᤿hH�I�|�?�wM\�SC=��� 9�S�ʕ���٩U���'*;N��[|#f@�Va�&.!r�!��zv]B3�𴆧%��h����~��9�����j^���~������[.8���fU�� ��Ƒnz3T}��]�_B�עf�;��x��9"��ʶ��6��%�x��8^��E�L���k��`.ͿD��`�ub�(i�5@(:�˃�J���->9{(b%��p$°K��FJ�dh���.����A7
�`+�Ъ(ٱ�/@�~$�w@ƫlT��c�G35�KV��Z�:Z�;�&����]�?����{�?��⩇s�1��V�����t:'��u��塄��R�k�)5��Pm\�Xmf�-��Mv�P����k�G���+t�����
��l�ݹ3Ԟ���4IW"3��Y�"s8��ʖ,�C�.����%�ƨê�O����@���Qj��k?�3<6�Lj�v8�j�t9^��>�H�r����Av*�a@<�IQ!j'}�`��DM%�k��ц�Ǽ~w���4��#+��n����Ք���K�c�!&��o�X���u�h��r���Qb�=w�=�Vl�x��o�����AXy+_�fw�e7BED1�"qc^��z�����~��0<p.D��,Ԣ���jW�S*�⨡���#}R$ͭ@RE�cU)U�����f�o��v�I�-(U�$���7��cA�W��*$�5�%��iNNxR���+K��gD�d���Bcc���`S���r���Ԩ�OF�R�ho.��y�C�)i걛t?�v�?T�%�p'd̸`��>�H�MU�!:7 ��ʪ�R]��4p�#j��.]�9�����]��|\�d7�z�
C6�}<҇Uu��/�rMn���L��46AC�#o�1�Ρ��߀*`�ǂ{#���;eKz�Q��%<H��u�����ÀNvY�ѽ���fo�#ju��"	�������x�����]�?�_���-��!cB񃠈+!�B�<�J<�J�o���yݶ��wx./@����!�3@����DO��R.�����:x�dm-R�)顒V�q����-P�^�ZQW��|�P�yD�s��b0yBċcI�RDT��26	ш�_8={���li�}�Ͷ���{_��A��l5�3�|�|,VCsm��olXH+�^(M���,A!c}q䆠j�T�]��
�C�9:u�HfG�	/����ky����7�X��҉o��T��yC�����ֵ\i����k�h?��tdC�!A�mƒ]��S;��v�w�{ҡf���R<\e^f�j���������,����*�;\�'Ӛ�H���c�1M�O�4k�����|�>Ԟ�4֊�)a���{n�W�ԭ��RZ!���u��*����,��&��"�O�c�G����eGw��4�OH��眷��[�� *�dPB^7���B|�&/�t�I�?<��d��U��|v�v�&J�"qV���[���s���T͇5��)�3���O����Jh`��^����TR��]��5S��ش�{�~��=� �#�H*����K�~��=��AT@��*�&r<� ��x���3���cz�`����t��C���*AIf*ݍD���Q�
p��MնM�C��VOwP�]D�V�t�������4P8�͸R�P
/i��R�7yp g�R�]-����b֍-���U��e�fgm��gK�MIgBO60�B;]7�CY���j3Dڕ� ���!�s-�U�������M+j@<na��B�m�e��Q��b0���أ��<��V��[��:� �6?41�գlS�L�<��s:?�����/��� )�~�xȧ-�~�T�}A��O��fo0_�2���0t?�A`f̱!|��m����3�z|��HP6�wI���u�d��3���@}�NIŊ�I�Sf�\2ӑ����onP����Lp�d�a���<=���[~;N���x��Kƛn�$�5��͇� h�Q0C{�}
�k���b�]1� )*o���(Uxz�\��r��ō�ah��J0g�;ʊC�3��w�X�t?��At,��K׎c��1�fN�Ej�D㪗�~�9ID��X�1tq�yý��Dz^.��	���r��rJ��$��F,��f�}0<�,r'e��П[GQ�9�F�����G6��y[�;Ƣ@I��9`9fom�*5交`<EW[3�7)J5�يZ�/�vbp�������OÒ�$���F.��OPJ-p���4@���+vJS�j��<�=QK6{�;tcgw%؝�#�7wVk�!Z�w�4G��ޛU�ST^�ִ�&���|~���SR�^|����^���8�LZ$eT��L�g+��Y�Y�~Us+6�퉺j=��籏>��Qt}�w���[6*t�S9���?�z��&�^��I+��r�u�/d�ۍ}�J���B�q���\�/�� �&�u�������<g�Bm Q��� {U���v��Z�ߛd�*��O�r�,�}��Xq�=��a�m%:m�:�*�t�U�V�U�iW�sx����&�ce˥��[GȎ�J+���-�:�r��U�#��n"&��ވ�R�1�)��[��䧄Gv�'�ޫ�p��ҋ��l��c "V��2�tWy��J/I� �%#)��VdT�b�ǭ.����`�g���k�j��l(�G8C�����b�*��Dv��n���$�ִ�r��̗գ�"-��e @I��3�(ׄ~SW2]"4D��@M����_��k���<�І$?A��dʟ�^�4^����7�c`H����G��~�"�gf�e/����3@�N9�7v|k��g��:p@�&l,���j��Y�ܑ^������(7/�jHC"��:=�PDʽ��@��ECm�U�TMa��Ǫ��~���R���]};
�÷�ed�����Y��a��3rbN8`���j�y���e���@x;�LcckGu�J-;���E���!Ğ�{���TA餸��OUy;`���y�xܽϧ�n��rN�q�@x����5��凑���cѣ�^����{�e���Ym���Z�q7��i�.��h6�Kj��
�a���8?{���:�꓁[�'�*r9F'�ަ�L'=�z QK�u�N��`��h@�9��ؾ�Z��I�kr�nd���(�bc�Ì�7��K��+ƚ&Fn��@�?] � G��{�Y�kT�fO�g^L?�u}ǈ<��abu���a�[���gk�GE����žh+1��mC_-����u�h�̇����Ʌ��)���;W��t�x�O\��i Z��������\xL���� ��@J��a ![�D�F��/s�s���6O S���R�7W՗>��s��j�R�K);t��/��4i�������M�ƚ��Mӷ�$�k�u)ǯP�^�nYi�Ó���ae��}���R�rb c�X9M>�;��F��!��S4�T	ʡYл�W���w)�����rO�y#����LM8����|���p�щ�ݔ��D���X-+!ʂ�d2�3�ŒS�!Fb�8����N?O�Y徙 :H����U�
�$��mC�����&��O�{�<�`Ŕ��]�^������B��`\�|<7K��v'<k��c/�R!�?e]�@]�J������E��=2��< ��@�+���R�����܇�����&�߄Ε��&F��Nx�F��sâ>�kM���r�O�ۖ�\jx�cz�;�x9����U��܆0F���g�����
=B̶	"�P�᪁�tǈj{�(7�$<��yЬ��AO���CT���R>��.֥ ��]���k/���T��z_�3�����[��=�~�ޭ�UFD^텟`�]��`�<tФo����B��߹���R:�ĨȽ�2[�Gw����o7uj��:B��-��+�n�l)�{,�M*<�h�#���H�"bS�,�?��(�eX�*_��'8c��r& �(��H��z�y�%���J䰁����(p3�)������ �m�E��Ql����J�flv �Ī���
5+ f��̦~Z�6�3w	�t�`I�&�z�����J�-�������8��mW�/�%��?oi��+�'��}�yYK�a{���o���6(�ܸ�5�=ڝwo�p��|�Z�'S��R��/z�
�i}��J)YY��Cz�?��.��&����L��Ih��dl�{��� �i�#������8c����?l�Ը[ng�F�b�����\��#��Z���4�0��u�	��Y�,}�����r	������,���×��70	ʌb:�����4�����Q ��wsX�
�&@�T��)�T�I��_�b�G���+��.=HuI2b|�
F���۔Q���!n�&�>0.�F@X6T���G�v�,8���^��d��%�⥸t�t��n���x�_��Y�ש����ڡ�Fa����h������Jw�c�X$|K�G��ZV��Ǣ�͙Xl=��P�S;��F�f�V2�mU� ��=�Hm�.���v�h���N�N�j]ka=�y��p�"�`|�-�^/�{� E�v�$}��մ!�$�Á(���C#��5�������6,c���1{-3�zg�z0�0�`�up�ΗN��*HBF%m�)�`�!�<���G]�������P�Lr_�\���^�6"���V�ԙN��B��徎��'�,������(���]ㅋ7����EP�xl&w�B	J��hҘ�o���Qz�(r���@c�=�����j%\�%"|����d�l��Ax	���L�H0��cKݮ$HZw���%��%O<�oG��3(���H3�3���Goժ��J���xMM!�o���<yX����-���y60�odO�h�s�TLs- ��X}�l������
�N�z[ɋ�"�k��h�K7i���E>E!�9�8
h�nX(@�>J��Z�IB"����x�nvk�d��SELY4#̗7+i{3Ϧ�If!C����z�
`@��|��x��A��7�ɹ�Ffi���%WX��n:�y=޻��(z�d��U&ٵ胎���\�X�'�(n�<VxJ�x�%��_%�zS_=�F��$ދ�s�,�Ak�
X%��21Kz�,(}]ٌ8��k����X��0�ܛݞ��"Te3���,rD����q�DT�j�'uG/r�ۦ4?^<��a���$aCU��ޅD����=c��z�v·��U
�:Kse�3���l.R��T,�o%O�_��{�fc�W�W%�H(x.v���Ms�~.�,���6����}a>��?��Ƶ~�3W�w�c��F>�	yƊd�I)�H��~XDq�ˤ����;0@��)"�z]#�qv��������K�s��o��]X��Q�����I��m��meR�J�߉�q�*�o\��A<�.Y0H^����'�D��M䃆B��Ɩ�:�x����4mN���Ǌ� ��Nq^t��Z�tz��9b��B��_��f��5Mد��}�$����8�M ��б���Hp���a���vA�f�X���@X�O�����n�dΚd��?��Hek��������4�����G�/�t���+�	JJpxS�=�^������� ��2c���.�n�����}�~N��HL���j�$M��)X6+��	�D�{i���������GuG�������_��[��@����NuM�USNIb����J�,�2���B��{��ǂYa$@��=!d��Ԝﰨ��z��FY:� ��:��`M��@��/� \n�y�]ْܯ$?7�?M�ռ-�u�wU����`�7o5ZCy�t0�8�����<�lO=�EB
��p�����`�!N��g�U%���L5ب"�����|��>��ֆB*=��m�������#Ie޹_s� �8�Ù�7�M~�=x��N޻��Bw�SLe��F��.����0v<�+�W���s�\s���N�Z�{��x�������Ԝ�_�3��b8[m�	vK�A�k� �/�3�]���~ �\�\�噠���k���
V��n��5�+.��8	��Lw�~�񬏕f�hx�y49"N;�I����<�j�e�����8}[�c�;�4�����m�Д
=�3Y�M��w�w��NL�\��	(a!R���[�Ջ��y�d�t�j�e�hb�ݨC�Q:����8A3p�	���&�6{�A\@�y��s����p�V�ˁ��J�~�k<Ax?���E�5"Rd�sY����C�����Np�������ኦ� l�'H��*N����m9�ś|����I4c�G$������y���
��lH2s
�Z��u�.u��c��F���`�Y4��T��T;2P��<~N� .7%�Fz������N���O�Wƴ�y�H:V�c|�$�q>���P�����md�s'm�7<����550��e^����	�[%��<�s����#7���ȍ;I��6-i��L7h>W@m��;O^�d��E_6�a:��Hpۂ�Nw ��qJ�k�����n@�7VcI����w=� #�zG�R�q�`��Ŗs�(�xe���y�?��v�^o1/rW�[��$���ۻV$�GZq���u���Ǜ'U��b�qN��9�;79������b�+((s]`�J����+���v���J�:oT�F�;�`M�q+r��S����ݍ�з�~A�>��r�s�b%�?�	�)x{���k2�=���x��(�.u����B>������B�`���R�~��	};��
g� \����&���|�$��pk��(��t�1X���8c�Z�0��6��Dv��5KFs?	��:���']kWv��	5��L}��!�l���g��W[��<O,���b�ŉ(s���Z����P���Vm-O��E"�2�-�x"��A>��qW>8�F������%��BB��?M8Q�ot}ϙA��ivF8��ȼ{�?{�]���h� �JQ!��W!�:tKM;"�"���.��h28����f����O0�g�!H.�ۃ�}%y���[Y�ւ�8���������4V<���x���,��}�4��la���~ �`�E�t��;�6(��eL��XF=���6_)�:�ǜ� �Y����+=� N��z�1��?��sE�e>:��`@���TLcĩ�0�MHÖ����S�d,�m�H^7�!�����߹L��R�6�l����hI����^u	�O��B�ȷ�"����>��+9�ISsp�^�)��a�]
�Ya?R�X3�8�eډ�S �6n䁽} Qw�}�jކ4���������ƴ�!~�1����(�_٘�AS]�p�)f��F�R�Y���V�e�p5Uz��z�[���A�u�Ly�t|�Y��ھ�2��K�l[6�l��rH���l?���F����$
�
$ao������H�z�/=˝Iz�ІԞV��0	� :#�I�9����%�w��I( ����?���;ٗ����Y�G2���չp�ѱ.do��%b�&�����E���*|�6�j����<��0F�U[����6H�r�;U8�S01�D��⁗��T~�>Igk������q�Vb���tN�(�9])�_�C<�V?�D�l�k��I��H7��I���6�΍��e�dj��;%q'�r-0K3���A�����k7<���q2��Q��#��<N�d�tJ���f<��֠j���ߜ�n�,<���S��^ߑ
�Q�Ɓ�k�_|q.Q�Z�)�~g �Ռ�1
��_�������.��]~+�p�%����P�M/P؂�n���T0ҽ)�[D7�����& ��
R~��ϡ�k��g=M�d	~����������cnn��{]�&���v'���t<}�5 ��a�1�7���֏����<~�����Q��[�����٩Q�:��L�C3+G��T:��P/+~�a��Z>�sN+<ps��},2}Q�֕l����+�}���/�!ɻp�YI�Jȕ'()���4��p�Ó4�?�fR��Kg�BXK�^Z�ْ*�-alS�$v�����bc�l�/T��5�:�A�������ۈ�eϟg#lc��{�%7_��x�GK����7�vq�6e!į�hL�햰6O���w�I@��+k���x�ɒ�s'��=����|r����+�X���� 6ZΙ&M�1Q�>��R�F��!n�W{�	׉��g��!H]�_fK�Ň��h~���lUw�@�5@�Q~���gh@������D���:Xi^G�ڀH$���,�fex�.I�_�,99�|�o#���su{�sKhY )5��5)�.�8��c����:7� ���-_o7���W}e8��P��li>>LG��R��[[�s�3D'�Vq�ӫ^M�����f���~�SQH:�;͈C��݇Oz��;��:�Yٜ����y�4�``�L�q�z0�1�G:fk��S`���b4�S�w^�'a6�7��OS���9W���>7�.@޹���� 0�UT��[]��c��%H�K�U�&�������ʐk�ڇ��M�����8]�Ў�ң>�H�&t�!Z�mG֒�\eM`nOLVqY"�hړR-�#_K$���&q���0M^wf&�IrbS�$+�C�9��VeF�pG.P
��,�M�"B2ʭƨ�E����$,��4��u۾8�Yc���z6H�����l�:te=��7e�S� 
G�['�
�[�mA�������[:�����k^����,q�d9"ڪ��g!v�WL�����"��8u����"�}�&z��~|o�7"ڀ�)����=���V�[�D�.�پ�y���ON��Z�?�|5��UO����H�'3A�hД�R$m5�G0�j9V�\��F�8�Tz昴.d�����0U���M�ꤳ�գs�b��:�Q�X��E|l%Zo����L�k�9]�f�.���
 ;���Vug����'*���/rBӣ����:)�Ε����m����[o�����,����`?��{$�M�׏���@O�UbR�b�2��5�0��)��}�nDE���L��D	�����H1��0�%�ƽz�#��x�(%�������lA�5cR+B�j�q�ؚ�w��,L�I�_��, �H࠭���5���Vm�ќ*�}=n7ѵ�*2.���'z�V�m#@����)�W� ,<�Vs��S	�!qD�-G���"�����a!���uʞ/GEds�}��kW{�=9�D��'���nd�[b�7"r%RGR#��!p��}�>%G@2.xC"�P�#��O���&C��e=��&h��A��A�����
��G��vШ�3-�S~&B�׷����X��-��+�')ky�Xߕ�G�����W�WSP�W@�G/bq.���$�QL�֡�L���wNb��A��i+��0A���������o{��Q`��_s��j����ݏlD�����<��Q�����&� q�'�r\Rq�r��E��\��7�\�ˈfwы{QW�{Y�@� �%u� v�vEQ���afQ!�7���p�,���׈"OP�e<�V/m�
�8ClTk e$�.9*|�C���DD��}Z%���qX��Uu�m�ס`���֎�k�w�q���D�W��!@�90w�v�O��(e�I��/ed�2�� ����Ce��%��d�i���=h��m��k�>��<��5�l���=���2������מc��
��zu#isU���*,ktLr���8�e��6͕5�@Z�Ts5�evB�$�{`5Y�S�:����9Z��c6E�U>�S5��gX*��	��˧U	�h�]���.��L�� 2`�
D���?�Аp��m /��EÁ�ݼ1�Ѧmn!)1+�>N��4�:����0Z��?PZ��Sأ����l~A?h/
�61�j���!/����O��;�Ո�#u�ܹB7}1����� U��ri!D$å��zkʨ�ky	:��FKa.��@�Oc,	k��jɊm���}'�)���go�#�����^� �F�i�q��ۄ�mS���&O�X��'�}��oNM�g~��$��"*t���>�v����T{S*-A�/eͺg8`',���~"�6}q��=yu��SK虿��tc6�)�ѻxM9�+3��"Je�%{���I��ɴ��ר�c�3\y��G��������� �ȸ!�gH�ET�
bؕae��D��Ju=I��}�%E�N[�g�Q;}�D��M`0�gL,X�M_�尭g��5}��b���Zߕ|�ȓ�ZP����	��HF{�$z3Z4
�^i�����jIg��>s\K�X�Oȸ��Oj����Ym����l���!�|�_����\�V4T=�1��C�(p��7\���/�q`/$����0�`���#�����ϔ�^2ӓT0��q+Z���e<ޑ���(W�Gҍ$�Γ��hT�6"c��gwac7{���J��G&G���n]�ߙ
�3�I���!��-7��2�o:��{/�ّג(��Oaݫq��T�m2�n���7iR�Cx����k�0����-+ywSߜ~�&�d�Ę��	�؝F�O��r(�7*W#�Mn&m��408r�����TL'a�aAt�Ҭ�'��V�O���ɑ��U���|E����,�A�^(l�qn�*g�6�xKj.�T}�k�����t!��Gvw�_��M'�}Ҷ���al�$j?�#z~I�U�����݅���6H�G0B/���d�vΠ�s�9�:���"���U��y̓4�D��7t!#�r�`ac����_��iF0czZ�Ӥɫ5a�i� ����`�Ք��^ň/��jTb|ak�,N�w4hG����>'�����7�(��{�ғ}2�#�.k����a^�)�w���z>���;��
�\od�x�^h��������\~h?��AT��Nn��>W3u�(F4���϶�l %��{�N��u���K%I�o	.	L���b5zB^��i?bdp�.�9��#�E/'B�o{&i��ۂ�:П������FI��f�ުK��G�_��=��S��H���g�H��Q�m� JA��X�{[����� �����6KUU��A����_[�(�X��c^���D����#�;������Խ�+�W1� p����bi ��ѧ������nj�G��i�p�G����|�A��h���j-D����G��	z:k�qɃ�~�U���y��3z=�pP��B���
3��w���vMZ�B����7����`t8�ї�q�U�T����\W�db�������?�@  �PP������Ȧ0���t��>G�
���S}�/��HW�B���.I���mY��9DI$��I	��n���l)O��>
�<�f��]G�Q�f~WRk����-{�׀���8,ke��/"������/���Ah;���ew֖d}<gjS��Ut�h���cG�A������*�r�a��㬄W��QIȖ��9������;�8Y���vr��@���]�fK��Vaܜ�5��Ǻ2����ge�����+;�hC]��A#��ŀ�j`��1�G_��	��� G�y�����L�_���(��U���#���J��&�~�� �`�(c���� ig�	����F�L��g'0�-��p����5�=%f��[�j� U�@ �[싋  ��w�KOפ<�����G����tG����P_�N�y�{�����M�0��1o�:�V���N���,� �C�� X��U39�g���Y���&̗�a6C�E��*��!vN޻0,��J"���bE��0���:�w�T.�7ӷ�m��f���҈cJ���<�1\E�Ҭ��S��!�u`D�0���X���c�鋈bƂ�X'�M�%BM�E+��rݓ���o�7�S���%�,����%�����
�v����@��3��>�,�ZFQ�jI�m�S�l���2p�K��p>��E�ޟg��)���
gTV2$����f�m�E��_#H�RoH�g�XF>�B��+�Ex����}'ų���G��5a� �����^^�� q�b�S$al�{ivy�FUF`I�ә*��&�x�%8���;�j#�H�^��[1{0��w���ޞ�x�%�_`���R�ZB=�	���'5K9	9���-J�Y�V&��tihs��{=��OڰMgi��N��'�R��!})h'ɫ�P�k��hv8�k�i٬���]r 녺C`����@�,��R��|h�+��C���<�}�Ǿ���FT�ϲ��O#;4��E�eH�o`Ox��z���A�@���f׬LJG05_��=�f�u+�!Q#[T���z
��w��j��>6���&���C� �&�;�����z��N���t�tk���p�ս��$"��u��	��x#ٳjۜ��Nù�����`e!�Xz�3I2�����l��a�I�������e��+=VN��7�j`�
.	��8�`��9nu��S�$�/����奴&usrj�<]J 0�o���׎�ԏ��Gs/�90��ȂY�iZν�~,�|��hF�O���ۉM��e��#�XJx"�rٟ�cM�ẁ���5Bs���Zv�G-�+��K��y���
u�_��rW:�}�?ŋ��_��@��$v7Ø�� I�Nv�&g����b7P'�q�c�ē?^�#`�k�TN/|(	����t'dMl�[=�&n�
Qf]K��U�����B6_���)ʖ��#k�@~�q�Y�uM��JW&��O�Ջ�B^aug���7'&)]����(I�Zi3�i�������R;@�]#sk3�5����N�]��yW�Ǹ�=>�ܚO�^7˷!�l�c!�fh���X4����\��E�w�?�&����Y<kG)��Q>� �2�jhq|u Z,
.�d#���W��}r��K���u3�yxO�uy�3u]��hR���:��]��@_����WQ�>��6x+����7^E`���H��jRPU_���?/_�C��g>�	�}W�7�q�[j���]_j������C�9v$.<�8ĳ���I�9w��Ƣ絣e*A�F2J�i������[�պ�+�$�kv����ָ�>S����P�ص����,��o��x��m��;�;%&B崁���wϝ��׻���4vG<�R�]�kk��"��~u����%O�/ubֳB>2DsF!q�������}�ta�eβ�Zx�U-�:�D�z?ҟ�*��I�����)���TH�t'��N&�؎�@6©� ��;>;�>�����X�}�����5 D˪�4&^F_Y;{S��;�{*�s�	q3��!\!l�7L����	ya��ЕSSW"�^����kڱn�S�o��}��c�h��=H�g���=ZOP��k�%�"*��D�Y��]%�PMQ��֬`�;�A �7�Z^k�\�Ġ�@��{�uNI���3
$B%�q��d⟶���H��j�Xڐh/�*����g�Mќ�#$G�5;Q�k�à# �"�~Jf��l=㪌~�������!�oWK���?f`S����H�G���.v|*6���+G�$kE�W��8��
�����T�9t�W��� ��Y��]�0W�Mk�V��{�[��ub)�ia��� �N����!w�4"��c��?�U
=���Ѐ.[VJ�0��ʏ[�+�/\�1�_Ē����i��؂�qg��0# ��YT9F2�6�(���X�.���=M0?��ؚ<'��f���8�=��B�w/�E=��X�U��|=W��?��iR�CM�[h�wUZ! D��e'5�ۢ����Q
n�1V��<-���������<�;�tu�Lj�tw#����= ���F��S�ۨ�rC��A�qAi�����Y��	b�Hw˽����C2�YOł����]����W.>���`�p���o��aQJL���j;譟��}Q��&F�3.�pI��!�n᪐	4�5�;%7ViRl~'C.���Lg�N�h���4���?洮�՜��/1��ff�$��l޷k;a8V�ֶ��V�����f����_V��")�x(���2
��T�&�&(J�|��\�	�����Y(��%s�l�`(s�g�@7�hNN����Ů6]�����o��jdr[�N�2w����hmދ]ɏ��Y0���Ab?���~|�8����S��,������1,�5f�|�g�5���H�X���J"G#/:�蠨��K�3g?�/I\|�D!~�I0�j��58΁����祢��e2��ˢN� Icx�q�ə��1<������)�XV�wk����0��K��h����/D������W��6��) sD������`����U��q�@��_c'��y{�)��bz���Į���E�u�t��ȈI��A�s)F	i�+3	�Rz�ƕ��ܭٟ��ݍ�.Q�MF�������-���U���x���C�O�D���0w��$��
�!�cM�%��s��M��[�����/�tP^��V�H�����s��R��L�M��# �0Z�N�'-7v�b$�[�A�8�D��3�!.HA+���{b;	�J�8=!/CڈD�U�:)F0A�)�+�NkE[���۰��D�h[�]vL�)��'Js����C�oj�{w�,!5�F�(�����録�L	�A_��MA��KO��A#������0����`���eP��|���М9f�*#E��G���r�Z�JP1�d��٤��yG���M�ò����Ie��&k��g������U�]d�HŹ�ܥ`�O(�R��kZ�Y��E��}m�tV������q�!�:��v-C؂��4�/��d��&�f_��K�ܹ�]�KN���?�_���Je(t��I`�;�.��?��΢`�q�`d^?�]m@��!�&9Q�o�؂BV��'�w���vG8����IG׳�EOxM3Z!;�4��G����zr\l:-��Ĉ*�?�[9�s������J�%�C�B��7��$* ��g1���F������[;�IW��N'pUd�e��<�*�����"��zR
Ä$ݷ�y�\�	"fPi�C�8�8���l�o%a@�@�[�����Բ�:O؊T�DŸ"�'�2��](����د���/�)�&_|�_�Ai����\�a��ڽ���"6(�	w�)��^�~$���n������y4(P�	�H
��������$�-H�ɬ�2򯳿
NI(�z�CU�v:�s�'	���Q�!,Zo��mM|��w9�sj�׏ ��M7����8������ n��I��S�sԿ8|�wt��z� h��@���zJ�O��(&�����G����}�i5�l-��+��u���9�!��mX���_�v��/�u�������*�}���pPY�-�:��u"���,�e��8=W��Ci#��v�NTD�O���B���d��E�`���![��`H�K��i�vykV�&�T;Ϫ�Lsn�4��it�Q�o�y�{�����d����*������y5K#�4�$\�`��?/�~�3���i���"�=���>���W����N\�����Gh�Y���~����^kCV����U�F���J��������o6co��b�~��$�D��G�c��^:��@̺�����m䱸��P�\����l��(�8\��@̣N:�_�%}k�0�z	�~�HM!eux��+��B���7�]�W.��z�a>�.�K�U��!j��䕫b���f����{��iB�mp�q,��w<y���Lt�Y��\#l~ճI=w`o�y�];o��|�LJ���ۮ���Z�]�J�g�T���[�f�@�)���f;p��a��xڇ7?�Y05�V2Dgf|NV=݈�4�^���P�㜊�c�;�+ݪ���y(�ك�}��㶅�:�OWaPѰl��|�c#s��I��Q��j��/�O��� #.tT��>�u��bz���-�|��'�{�6?V~���~�O��e<��zJ�n7�˸��ߧ��[F"�^������ r�8BF�!<#�m�^L�����]}������&��h��جe\��YB��
'j<����}�l̯(o����#ܦ(���
��z�M�T�It�����co��6d!|�����;�z��qql[%xB'j`��.dN� b�a�S2�'^D���Jz�
 7X`��P��A�wı��f��#���o20q�o�C�#�EC+t�^w�,�L�O�t#��S<O�1��S`�8v��+(�i��dd��~�r7�l<6dꙢ��5���ܖ��_F��eJ��k  �Ÿ[�����gt�W�=>�f��5$ڛ,���w;Lxr��	�f_������=#g��c V��){��a}"D���h��H����_�-�\�$3"�q��~ʶ�\�1�` Uz��C)��c�t�"��v�"��)�>ۢ��O��b���%���K��J"N61��������[�0G��&��NM�;�a�.R�x�G�;7�'y\Os�z0�Y}�.�Mfi�䕵�Q�;�<���"�t����N�/S!���~�"(�[�x�D�������������e78�����Ju���g�h=�'�� 
*.������Z�)��16l���	�/�w�(9�!S��%��1�����s,ү����$b��n?B��=:�=k�"����	1�K����ѵ�+�e�h���s�q�J��M�'��-(N�gVB���I��I��E���L[���iܦ�vXO�%�F�`割��D��i*�^#<���2�T��2����.O�-�Ҧy��/��eЍx|���Њ�5B�f��d\�@N˴="t��C��K-�14�4�����]������{R�f�{a��<�� 5h�쀜3^#e��������󏠆j
��;��i��>Ro�\�%`�>����ҵ�����_�Z����d8�5Z���ͫ�#�R���+mt,��3q<��w$ʦ9+�R(/�lo�|ӕ�Oi��A����H��䡗��p�7� x�鐌8e^�O�����۽pt�s-����Oi���_���Wa�@���K��D�סi�1�;�>T[��v�k�����xA���l�k��~��sk�Tz�r~u�{.Q+��Z�w���yb��V��XX'�ps��l�Ԣ��G�9�� ����>�%�R
��
.���I��������ڼ�@ҿ2s7�T�<�=�P?�K�_��4Sw�mo` V?� �C�W�l>-'x;����������c7�O8�_�)i�M������q�=Vc�� �)c�u�3�a���GTXyd��{�_�d�P�2�f�<��?��- �����\	1{,/�f�E2����| F��������a�G>Rn.e&�Z�S�~Њr��L��oI�τ&�Q]�to=��f�r�B;D��� {����A�=���Q�=�ޠ�k��'rn�|T������HdS��7��-*��EBwsx)Fu	%�i���E={l� }��S�`Pl��
��c1�b���vA&�+m�r ��(�H�TS�Z��Ni"pè�IP�+�{z�z*68�W����De��v�%U�fh�L�����q���}���l�w;9�����$��b�(�mF����_�X�6���8օ�ϗ���ek���A��PqzIҏa
�E��?�K�^��2��!��T��cQf0f�
��d�tM�U@�H"��_*I��gH��]�������cb.G??eG9���k_��j{/����nȇR!l	��l�̗nz�Ք��B�T�D�g��o-����=賑��A��g	��=���$���R�}�����(����r(\�ڠP�t���{5T1�F����ycW H�(���V�_ϝ��+m����!xAذ�-̠���N�0�~\��t!C��v-]�5{�I0�k�|=fMx�����Uo��N�B���b�3z^���Y�)%��fF[d�c�#�ϲ/�Q���-�v�2@��iΥ����t��`D��+�� ��	<��FB��D�\a��K8�e�4c6�=�ξ�}8�Ȩ�*���zN���L��*���G̡z�L�FL�9X� �,RY������o>E�-��?h�r��w� *k�>F��UQ���❎�4���RGި���Z�.;c.f�8��jIњ^IM��=G�0��4J\3��!��#�c*Z��F����| ���s�����`���X� P�/]�+u|��+��)�V�J��vW����_�$ �o�$�B4Q��M�!t�@����q�=�6^����E$Ac����¡�h����k��V�)8$��u���5y2y�	����`���Y��ؖLV�RȬW�5�n�p���!KT��|��'�����D������߭UT�}cn�<kn]��"=a�Ej�~*�m\ƕe��dG8���<�%�-Si�~��}�n&_���x�΃Eio�����]f�Y�R'����e��P�2$�=�BOMSґޛF;χ�W�|u�T0�`gw����_f�>38����{�3��9��'6D�̘�����,���8����jmH!��p+j���d��l�a8��ٴ�|bH�v�}�����M��7�
��f[�*u����	S��CN��Z?�"蹓��r~��쑣�i�WO7L����wL����\?n��ߠ.h߲.�R��w���Ec*�-j�Yj��R}�tQ�J���b:���	8#yL&)5@&m꺜�4�s����Zw�d�h���'ٟ�_\-�l�G��#����w���-`0�og���M��dXT %kH�i�����}�r��s>������r�U)I������[�oֽ�hi�U�}��*��ZW�JW�RdB,,��>p�v����E�`pDj_\��o� �=�CA�!l���C��}�Mw�%p\�fU�����G��"����0�'1Q4�Z�L�ڤ��dѼ�S⃝W������L^�Dy��:$�3c$�Y�iAr��E�Pp� n4�0gc�7��M�rX�Fx��I�j�/W�df���j��!* �/�����Q^��F����57��O��Q�R��B�̕�.I�t���� o��u:y�����?����2g�7����;n�wa耮v��[L(�WD@p ��/2a�y>�<_&[T�C��y"��}�$+�hKo�������#������;��>�E���Y%�]w��!J�خ��$~���^6�lM��O�V����{_D�آD�xbA�?��E]�nF�a)�淙�g�Am�v�!��b�wɽ%��D3}�o��Y:ߜւJ�>?!�;�ڼ�H�5Y�@P'g���d�u3ج0�N�4p[����-�:�S�%04Z#�`zjIm��e��}�O� ��Y�<�";���x���GY�=�&Ej<f���E��*	�������>��DL�D��
D���$a]VƦ>�4i1�Ub�9���&ބn��é���:4+S��ب��~^����`��b	��C<��T1�����O�t�e�ۖ]�@���"䨾+.w|��F�=�ק ֩���w�k+���G���]��\d$Z��u�2�������@˃N"vp�7� I��1U'&�ֻ�ã�P�W,��xT����b%\�'���i$�����J����G����3�|�`��
UQ�t<�#�'���{���<w A���O �Fca/ILk�z���U�v!Ā�ݱP�DKfɚ�CIzN��M�ܪ6���'�&���j]��u�8�wJRu��w*g,3+,(��1M�g����?W�w^��m�.�ޱ��ڲsh�W���YqKv9�Wh�񊎀�������z���V���˰"<�h�}@�҃ �8��2x�_6��e�ͯ2) ����F�p������Nh�dQ#9���ID��T[L�l���:�|I�h���H�U�%��g���
��B2���X�#�h�L�lv�f<�L�8��H�.m��	�.4�S�`^0�5w���Zƹ
 ��s��c�#A4�Hc�&-�+r#nwg"�#���ۓ]��)R(�̻����Z-(��v�&��|w
�W ��R�7��ٍ즧!G�Kb����n�#�mpբ1f��v1�?�{S�R�]V��k㛓ϡ�t)�N�+�e h�'�e	WJ�� �=Q0Y!;�M4q����O��8�Y�,z�0��Q�5F��҂w�ڌwgX�h��b���E�#���h:����3ő}ٵ+S��l��l$�wv��>�d(���',��J:��m�9y�!�)�A�̲����J�S:�O=ӉK��S��W{LhO"�-���`Ӆ�zs_K��+']��wu���_2z{o�hp
n+� �ȝ�N
��p`Q  �H�;��鴂?Yp��"iyE�]7���;0yJ�I���䶛oƀ�Fa+]q_E�"��h��X;�N���,�<=*�/���a5㗉���z��� F��"�H_>�K�Xot7Ж��
�
�2������x���'A��,�)�m��AX ��٨ƭ�������|�^������Fy�B6�c��\�U����'��f��h�R}/�??�=m����<�����c�u��t 8��+#d�ۘl�d=`\JS�c�/�/��SK��4a�j/�|�B�ouy�7z����dM��?��e�"���MV-N����Ԑܧ�1p��5�`�b ��t&z���<��6h�	�˪�u����@4a  ��	����r������!�,��4�lL�'쉽��}i�y��,k�c���i潠|���5d��E}���\ˌw��F�ǋx8�dy� };pf.\P�T?,t9К�!�0#�r<�u_(��Pل=T��L����d�%1�}f�^;�0*�2'x���mp�B���f��Z=�`g�L�z�K�n�	������l��O]wѻ�����Q3ٌ'���gh�ȡ\��k�0g��}� �j���(��}���*,K/ڤ�x��v�������q"������7�d�hU�/ �j��=��g��xZ�;腵C�dX�����q��U~a�:㱆���3z�о�e_���Kְ��X%�J-~�ln�` ��v�.+h�^%zl�Wb�<�3���0Q�1W ̨r�|d>hTm���%��@�Çw�R��O,s"��>�5pKE��%�Y<������Z~�7�y��#�zʅ���s�Oal�QYE��F�:#� �>q�;�U�]~�N7d�M�z �R{[;��Bkr6�7L;�w�5����3WP�s��B�7|�i,
��{�H����1)/������a�c�{�ް�mKҵ$��u��כ	�s'0n�-ٍ�����U-��I��Ԡ:hPD��*��? ��d���A��H~n~�#�{;6H�iAMB�O�3��3�rka���:q�"6j�&��������mW;ɤ��ƈ���^9��d'�Z�0��Y�$$�D[�	�^���RB��R�'���3m_��P�3��ҟ&�t �r�{=��p��-����:u��"�A��܆�{���{�RlYd����Zg��(�z�s���Ӿ��ܰTjs�Ó�rK��.�)'��R���
k���6�|F
/�Dp�5�N܉���-p,)�ۺ�>�dp}���(ܟ��r�너^$X� �6%�v��x;���Ii��~��9 ?[��OmjF�G�-V�\�A�P_�Fh�� y�|�U�˺*�RK��+Z�k��f%~$ �;��h�x,��o����/�;M��7Q��>�Vʵ[THK�F��(�*���hHe("�H� P���$@�P�M}>× R�>������;���1A�7v�k���['xɟ����*���y��a��y�����I��$	W�{�ߵ��]�۶�_�&���������-��z�42���9H�lORޣ>�8�R��)<��+�iA�G2,8v��Q�n01֚��eue�IC��&�5h�wC�g���\\���[�h4.m���<�m�Zn;v�;g�\=}����Hm޶	��_[y	�H�X�[HD(�ܕ_[f�.E@������ݤ�X䀐O4�N,	��~2Gq����2I�9@[��y�Eu����� �TvXy��'���I�L���)K�9� ߬��[u��Z�Z��3�Q���M���_	�L�at.��w�@�z��0��kHeL^��?���R�x�����W����<�q��R���X�6}���FM0e��	�^F�k�M���s���WmF����ܱ
�_F=�j�e�@���Q���k� ,�o��":�s�v��Q�$s]�\D�~����r6��\
oۥ�������
{+9�r^
�R���iNc���P�H��'��Y���J���jǟK"~h�|��b>9�n�]�o�oqpA3��6}����k�d���=�Ft/�X�{uC�*x�b�S�V���5*H�Tuz�?h����H��*��VAr��f�Ȼ[��/\��s��[�QB},�M �hC��VI��>Z�7H��$m��>b�lx���TQ�G��6�GIXCFzi����#�cHO�:��ffvx��4r�CQ�����!�p���� $��z�6������ژ�W��[b�WFA� N5�W'6==KB��E�ȫU)_ۍ�%u�:#э���lf��[y��xy��2��?�)B��4iYm
�D���� ��IH.�&mJp����R�a����55�
.�5P�QO��TO��s��Bo�aw����(0���Y$���ҡj�Q�(Y��s,�!C��!�]JU�b�d�i9T��ʓe����d�mJT�>ב�����۰���`=pH�*��t���_����t,L�D��;�;W/� �Rs�nr���t�����͢P|C(n-�� �f�����KHj��T�%E��H�����b�����F���͜�$Lbg9��0�D�tx��4@�C�>�O��X�?�!��K���E��].���0�xUΒ{ǘ]���HT���n��|
�*P����#��}/O3��=�����jV~�\�#=�l.���6[	]Dv�M�����I��&�	�V�s<������dG�m7X��/m���x6Cm1&F`r�{D2�|�� >f2�q������)�2�^��>�+�꼌ԅ�pm;.�\]Lzk6�R
%F�@��m��y�[�-�;s��@/?�֐՘��J�H���j���"0G0��&!�ҾL�)`��?�O]ŭe��YU�pq=��c�s�)��E4��c]p$�#*y;Ad�ض������瀴sF�����o�sm�@Z
hhz�O;�L	�ok���n?$~@|�#�.;�vY+xN�9�̺_�ĩ�R-�EL����4�j�)�I��ij�
TG�
���PF�D��̛��-p%�A�p���xR���.}��Xg�b0��z��Re��C"B@/�����H� ��ϕ�{��%��F��$<��i�*����۩A)����I�@���1��y�֐I/)�^:~0.ec5y��CC���{Ŋ��
�e�|���CN���k��m�%1����O>���ݛ2Y���n{�'C��Ì��FP��&Zļ���	�茩@[��2M8��)N�i{M��db4�Okϩ�����LǗ\J��N�v��us+1�;!b��7�y!d3a-��M����5��OI�X97
����^/[
%��Zl˳�X,�2W�ӍM,�z�ղ��xn�T�Ծ�[$*��i�5,v
��V���W-f�JGHh�IF�}NwmX��f\d���>9�����CNn�n'�9
4k�l�R�h�6�9La@�J%�_�X_��|RgQYf��Xa�c?z���u��
WǏ�YM�;$��b��������#s�j�4n��듋��;���-���r����KƓ���!��?p��[hM�8�����6|�������T_�),�Am�Z�|7boƤm	�%��e=_x>�F-�'!8k%��Y'��F��w_(��p�A��PξpXK�K"�#g�C�f��d*��t��.'N���ʎGP9�6h�%}��W����=��c����ꪳ�j dT��/e2 �v��K# \%�cH{sڛR͵1�I����	fQ?�ؾz�R)�4���O�x�̒���������#i�����h��L�ނ����,U�P*v�#��W]őK$LA���:�K��sَ9��`ʺ������_?r�����J�	v�u'�
�Cxbt�`fV��U1&���V����gO�q*.:��zP�:��s���V��϶����g�gl�!�]C�vs�u���ڸM+��z���@ѳ���R��ԍ<�`>2Ye;]洉���3t�� diJ��$j�2fC�w�}q��-ES50Q�{��b����&'>ͽ��J3<��wJ#���)1f��Y�J����Yx	NPP��t����y�؜� [���E�����(m�����v��A�Ԍiܤ�mF�<7G�r�i�H���i�e�Ҡ�A������wj�:�s�p�Xg�����WU�X��l�|���㰲z-KZ97��_۶ u�A�/�1�p�!sI��/���+�B���M�%.О;GC�<�4����#�_�
����:�Gg��ݽ�"��"��~�+u3���bdCY6";P#P��� #�%��$;'w��~ڋa7�c��i�V�Yǉ��}=ۈ	���Y��z�	�Ŋj�V�S������!;WkR����8�(A��JT*)���TP�ѥ��:��Bj�n��%<���d+q�x�[����)de���]q��[C/��k*����aF�6]�3DR�i�f�T/Sa��bE� 7��|�����H%9K�>o@n⫽EF�aP$���Ё%H$���P9�V|���{N��"�<o�>�?�t���@��+�-��wheǠX$�-M=h����%
X= ���TM/�H��1+�S̵ø��7�D�W���8��z��H��y�	f:������������a�+��e�˩���kX��fvR�z=������.��(��pu���=j�rx0�>|�[[6E�k;7��a9��<����w@r�d�w�����o�#���4S)�l4g)q�΍x�4`hPiҳ�b	��]�6��-ٖe��e"�-vS���'����|g
�::َvpB���k��F����ԯ�+���|Y�����uK�@�1�颥�af�B��k���xbUQi���9�'ޫ��Ʈ֞ڽ
YL����[����}a�ˇ6�(�,z5q��;���W`n�T����/��߬�ZQ2AWS��7Ӵ+�����\��1�K�!���Q�ї�lvV?C�s�VA�|�_�a��e�8
۬�zS��l�{ŏg�U���Y���v��0Jd��e�G4L��"��_�s����'�8R���u��Ԇ�E�s�͔TBK��h�Mp��?4�N��|��ȑ*]#�����+�>�Rj���(v�=23��h_sE�0��[}���x�Z����w�P���W;~U�H8JYۘ�%юH w����d�� f�l���HJ;#uͲ�X0w�V�`)F����r�.����f��J�5R{��1c{4^GP�+���)KM�p��rɣ�֪!�4��g��+�c���7�T����Xu6��,�����㻓�e��4i���^�}�N�?<��hj#���:��JiM�=ʟ����n���Qcŉ�azA�[�8ﭓ-V3׊�F��%��L��=Zi�xX����|��G/�A���Ki����-m�&g�6�Eu!W���#�Ga����` V�}�Gn��:o��ϗa� S� bF)tq$�y�x0㒀l>/;k�����-� $�c�;_b�D�����o��:Ӆ
q�Βrv@�����嘆R>�^a��4��OΖ	�d��}|Eg�h��KPKp_��U�j��,5����v���.W��vCn�P1��]̱�}��=�Ga�Nb�7G��"�.c�i���=��ѿsJ��"<*�h��ͮ�q�(��/�s��b_V네����K����+��+��M^���5QM)�C��<�?�y ht��\�)]��bF�3D�X *OQ�P٩Ǽ���lƚ��0'�b�2*C�	�<u��u7;�. Ggg��f3AO��1'���L>��b��vc&!�ߗiRu�N�z'y�`���ϔ:��V���F�9�=6����&���ߡ`����.'�� ��I2���6�(��;���4\��WCq�Ȏ��r�6����3��#��G-q�KS�D����H_�P��[��˱�p�Z��gH���Zj�ei�ǃR� i���}��~��	H�opL�.bE��Y("�٥��֫����\q�aJ@N�]��)Sȯ �~�猆nS������q��\��RYƫ���/� �w*-E#a��Y���*f�<��Y�6k�q���#��Z�X�ڙp�u�RT�L�/qpj<7|�t������g���_���!�D@�p�L�54޷?�Km�s����T?DmLj���� ��x<J'T����-�Knغ��XF	���?@�W�Ž���Vs�"k_�Z�6��B�v��.��z�d��"=~H��LA�%�y���W7���"�3�BC�r�H�~
������n\
A�.��L��4y����A"���F��"zԼ�)?&b�D6�XV���t���Uǔ�y��o�)���!�KC����<�����`�,.�gm1�̫S�24J��:��}?���� ��������+�2?Y9�hG���:݋��H�'���!���N2DH�\���W-���J��͗�mm?Z�t�v�B����#7�g�a�!<Fh���[��@��[��L�xfT��W�/{�AO��<�J�x.$��#�F6���-U+E��;7��a�s���s{�E�����9؟� H 8���̼������n�'�xhzKa�"T���P��m�$x���O3�(��Nc&�%[�z�	]��r-�w(�q��>ōק���i0 ��m���*ch�`R�N��S2��W��$Z�Wl�Gx�"��M�%�RV�?�49�JB����	rޕ����3'(1�;YBh�/tF6��㑣�XI�����1���as��ݝ��,a���Y��;,��-��'��+:�;�ş�h�%����a�����sagk���<���b���`?���#�R����_�19�-�/�`�	��Y>��LIr�Y㌣�k3��5�;��K�io�\�>�F�>��n&y�y#=�Zp�j~�J}U])^��9���4T��m�C���J�-����=ԫ�{��4�y�ai�O���'��-p���@�u�eA�f���ޘ^�ʃ>AKM�@�c�3��# �������}�?�S��+T*�������3m����=)���:�#��'�,��$}�E(�ME*���:����c&׽
`��ޭ(S����}���Kk�B�=m���.����0-��*�$�:�=�9_����k>���s�����l���Q��v�%=�>��C���m�S�6}#�� ��W@;�`_�Ά�{F֯�=�����3�?;���w3�e�W��.E�����@GX�=��+mLK�����j��F����i�ʳ��L<��?�����3����.b�p���QPP��x2Aqg�D��4�M�(ne��4N8ٹ�6M�Js#X!c���f�:��s"d��v��י|�Quk��"�B
c�__����AA  IS�������^8�cq��{[����p�
�rxU�j�l��5��s�����K
A���k����i83)vs������ݭ<-���4dГ7����&{�#��Q/̭�?�Ý O>u�-�̐A�e�x�3�a��/����NTں�,M������KiL�`ځ�~u����8ì����ʍU����Bȝx��wBm�?�}q!R����.?Β�F�"�We?��9��w%!��k���G>Mߟ&�y�-���,�����]d��f���~�̌�%� ̰�5h�w��!��JX�$Ӳ���{m�(�l��#���(3�1���� �_�Dg�fDwPK�&�XV��Ś�"2��B�t�0��`���vk_� a=%��zע������N
Wd^�a�^$�,��l�*��J	�Dv(���"���hC��,�M�8y�O�\|�u�����;�3#q2E�r�bٯS=��x�P�+M<���XAS���5��@�^~����4i>��k��K���L{�W)$�n�<7?C�"���d�"�r��5�X��C�I�Ř�a���wl&�q�>�8z<�7��i�W��c��I��T-l�N�����~�s/7�b���M�l���eh��Xl��=��-�	S޹�q��,��!&�i�2�V���-�d�4���Q9�<��=�p��"9�mDы@@�(�|��.P�w����2��  ��$&=w��.o^�����	�[�&I�]V���b�%�/�Ϙ�;Z-:Jp�RH$�mR����F�.A����w�ygލ�����7Q9�3li/�ֲ~>����vKk;��M�Q��˧�������+�}��/��R����rE�x.�+�^�Ub���4l�K�a�@^�mVpʭ[�|	ga��J��1��G�Ȍd����JZ�2U�3���g��gϚ(����I�5�u��l� v�_���L���=�v��i��1t�x�lǜ�P���sn�W�s+ہ�%�v�>dz��(��|�B%�D��ڭ"��n'�Y�r �Q ��g��=l�ۨ��WS�9�ڵ��pn0]m�%�扲;i����/��<��d�8n����9.m���y��!����������[�� ���K0�H�$�gq�7<L��;|8e���� p����f[��@*:,'��4B�D�����\��L%�Wqڅ:^ �� "��7!��$SV�	˗�|�����K�4[�
.�S��W�o�N�>!�&�I��en�{��b#��� c�緑����������NS6���b�� Z�;�W�I��n˓V�c�N��<��gƭ%���8Il�L�R
�	q纙-���H��Il�{��6�����o(�p#WQ�Ԑ�$�G��<��=<S�=�Յ���)��*.e�nU[`��pe������@���}/ƃ��!�����kq07ц��^Mg��@U�E�}�Ѫ��U]7�,ۋ�'�oz���@aQ�,�a�ў���j���t�ݴ����
�(N��S�(-��4F�}�C���z���d�O�ߵ�%�7���J�Y�Fwm6{���~*c���������*�g�Kا��RgVm��s�w�b��ک8~n���-Z;�@��.�����ˆ�WJ0'K^f�!׼{��+��4	{��q/�l� ?��^�S��U#���0�C���/��I���bg��\�w<�x���(���pM���ʚ�Z�`�N����Y2f8J6�T�<��o[���������#S�s���E����#��;X��Xi%a!�Vf�A����~��_������u�e�u(��3��l|g�U�]p��/:�+T@��7qEс2���O;9*6��Ĩ
Ea] ըH�iܭ���Nr����S'p�f�Cf���V����)>�A����c���9J�c����E�g%E<iZoҐ�X6��a�R3���g�>��lTr�3|c���q�as-�M�Ꭴ���:�Vƕ����[��#=��Mm_���;i�)m�Vm`�Vd�ڰ��,��j��H�y�l����j���+6WrB[ȧ��}h� ���8B#L���3��섓K�Z��=��� 3�����o�S��z�W2�������c����]��R��S;ֵ�<�4L&�]u��b�9}R�8C;��Y��b��������oXXk��i�2����Rw�����;}��"͢��N��< }SD
�
O���oD:��(H9N��ǣ�}2&�s���|�YEx3��岵.�c�w��Ʌ�� C iqw2r�:�]���Jh@�]��Ic-�%ejpY:���G��C!]���2��/������>�a�bC ?�^���#�D�PY��7�f?)�Sbb�E���,qW
�>��,�������t�Ry���;��\ XA���7|H�d[kZA8~x�����\�d>�[ˁX��u��5�Q�8�i�T�Ғe9��L�>����	��K W�w�$�T6�5����)����dU+���Ζ�����]�M TTs8���<ڊC�!�y\#�Mj���ҋ�q��v��1A��D5����OEJ���_�F��Y J;_���o��.�tF�G-Wg:��7�]?�+#�ux���g��3��z-X���zU��z��b�S�f������K,i
-�6o��r�@�xr�߱�#��d���	�;^ΦlncJx��,���'|z�OE��o��$��d৤�|6�$B�N������DY����O�-�
��J���w��a�w1w��qR��
��R
�W8�5�,K�8���R��s�2�(.��f:U��_�:�˦bU $��~�'r�9ƒ��)Vk*V����$�����o(14��U_�l�l���h��
itj�K�1
���)
�o�ʬ�R�ԍ�+�aSa�Y��A4�����C���U7��H9���y���,Я��N{������	�؆_s�T����\K����8�m����^8���T�N��\m�����\��ce_А%�����$�'\��Ě�*�+W�A'f�w��,�@כ��Q�=�+�[�G^nV�v��P��7 ��⛿7�jH�|���d�
N��@Y$Y8�d�9a�x�
N����K��ł��G�l�=�Kp SJA�c,�Z�}��/1fʪ�w0^����|QU&sܔ�1s�Qdc�����e������B&u�����*�}b`U@AzþxƝO��a�-�·��)C1��y136'"}����%�_����
C��~ө��%����9�r�x�T��M�Y�PU]p�ym��ۉov�j�4Z�~�i���b�/���-����ރ���x�L�����P�o�d�z}Ɛ��ي�6Ԅ��3!|�I�vG��u�����_�T�GG��������╝�foA� ���^�)��)NY9��)�|��+����	o�H{���\���ȤJ�s_�+��	��wwe�I�d��xd����iO���B��i�7RB��Nq�TC�ח�m������Le�c��(���A��[� ��yz��8�o��m:��-&�.Fm��0yU�Xc�j�,HF������ʫ-TSrg��S~�ӧ��$Q��"�5�+D5U�c�Bk������ʠ�Dc���0�#�N e�;}1�>�0-�>p���?��2��;Ղ�����;��YBp+��q��K;���jX_�*:pԷ�{}��:�Wh���U�j�j�<�����j#7P�1p`7>�#��Dڣ�6�	`�_W�{Y�@���@��R�0X%��sl>a�Hu�?O�#���ڜw��l��fj�����d�fhn�^^: �%5I��^�HtN��4���g�u�-)I��!�GH�!�q�Դ+Y��/�F�[Ӳ�T+ZQ��b8�a62�{Yx�--u�Fm�vsѝ�։�.Wg�MA1L�=
�q<�0���`�JQ(�g����wx�§=f���H^'��{���O�A�M���
<ӝrx���Ћm��# $�$ ڧ���p�VR�0�՚�������7������T��Uqy2z������6`_�N֦;zuH}�aw&$�3�O�MaTe�e���Cw4j�HG.	�E�L8�^Q�̊���,H���Z��Ȩu���G.aa��,�E[��[�I�A)5�i�%�z�I��?Ƅk�p���W�"S��aJܕ�E��_MNH�����u�^3A����%�\"���;ݔ������8�S�D�n�?��'���J�-EH��Z*�<'�@xG*%Ҝ�5="��)}Fp��On��)1]�}�e���n�X�y^�a�j�a�Ǟ="�u[��P�b[��|=��(���pVh_X�M6o��*�������t!��6�+��|�	վ.��b�'��ݻ%M=m�y�x�'k4�+`D���pk�a��^InAf�3
4�Y�U��6��<"�5�ϐ�J{����F��B����S����#DbC%�'��߁�2��V���E��9+_�"i.dҰZ��x��
�+}7�x��%#Ę0=�[`?��ؕ;/�����ܦ*�'�[8FdW�����\��cW�ʜ}	����!}f+Yt�<b�gLȜ!Ջ	��J��6���.��5Y��=d����8#�G��=V4,�g
["oc���
ȟ��ef�8�J�L����)f�����Y�.��IG��]�O�#7�%�Ac��Z�晑�5��R�=�ڻf�v��tdP��1����������MKa(�@�����󆪫��e���E6r���!�vB,f��k��w�GNA�Ix��9��PB��湖��/���!����T��ꑶo�:�ϋŷ\�/��C`��#�9�ա>]l�X�y�\x�<��*�~͹��X�LʍD��gP��ҵ��>�'Q
���6�0�[�@]�I�Q�"�8ێ ��i�{�E����p<���8�~��Bf��h\79b�P���u)�i���\�^0 �D�wn���u[�v%<��o��U@I|PXr�]���_�:���N����6�K�8��� ��l����S�z�6����+@2� �/F�UV2�۾�	@���r� MoD��D5�R�G0�_M�f��ʷV�܋aK�LP����~j���SuƢ���y��8X��s���8Owܙ����"��rPtr���;��N7�AM�^a���	�Qf�w<��Av��4���x�Ct�#���GP�'�::�� �i�Eھ�MObu�����&�=M��y��$I�xWM35�tV!~X���?�27���"U�%vy�h�� %�cZ���X{)=7꽽)��Qx�y��#�I�<�iF�2D�6��Oi;�����D��9��j�p�5�����F���N��7]L�,ʈ��u�Y�6�u����V讓���(ylP0:L}�[�.�P�\��������~�����B�!!{؞[< -W�����ō[������5 �Er��F�XQM��w��<�0@������1(}IU�(��������
��.���SH؟�W �&ԣ������U>��v���Dr"��oI�k��V}�@@
�DU�`���lD�ږt�*����(�hgP��w\�U0Q��=4cSC��^8hT�>���eRƬ�|���t�,���b?������tl\(s��/��z�����P��8��6G��'/�>��������Hi���bO�r(Hm���������ۉID[�0��N�̒�fW�C8�L����I�n3S�)�ʗc;k�g:]���w�h���y9��_�g)��`ݒ�7�!\�b�ݪ�F�FD�Þxt�Sf�p��#b!:f=e��y��kN$��>4j�ozf�-�M#ğ�c�oN@*|�Ar�����+kɧ��9ַ�!��C[�Z��ۤ��75���k<��5�@��6�SzR�{S���yͅI���&({$Y��W��qX��}0���ٟ�rR�ȼ��8vt���[���w
i�_�K6����F���B�B.��� K?*�~_;�����Ϙ��6T/Q�ؚC }�/����ι!7��u+��(�w�i]c>{�-!��؋�4����'��O��#��Pٍ`��4Tc|",Vn[�6�0D䄫�Y�J���1�i��yɈS*�_xďs̏h1:��5��A���lT�\|�=
1V P�Uwu�0�ޮ���C	@�W�㋷�}��Pn��O�p?]�b�+��ڊ1�#�k���tqI K�ˍBdރ��a�{+��զ����+�����u�d��ufi�	�i,� �*��5�R�����r�!����Ɨ��.K���bO����b��7�o�3/m=��t�WMkj��ߤ�.|���7=�t�ػ��љ�[(�Dk��L�f�d=V���U��1�֩ $ŚMi�'<Ϣ�^s�)�S\��R��	��Uڈ�s?�q�%�~F�jQ��kHN�%��u�@����q�0�|��n�fVǦ���l�7D�+�M{"f��K����}j'��RD�g�;n���rл65S�f��^Xel][��(��_<ܿ��Tw�[�H5f#��"��j�{�:5�ml�Ǻ�_������Q��A0�z�ՑPN�mT��<���T+A��s��`����,+`d�d�+uVmꝮ���~�~3�@x]�z��7ƞ�?Mn�V�¡O{}u羱� [�i�*�
�z��APx�I\¨�,��$ъ�5� ��#
{�&S���sa?Y������S{��:Sa9.D�U�!a��U�E�9\O�1�y�P��>�f-��*MY7��#�I�E�P���Z�0"{\����L=In«\
���?�(ꔒSC05*���E�JKZ&�󀨆���63�u2�
eW�����!O*��6����'ή�xxU�N����#�y��~<[i��rR+��U,��F�p�I�_�7{�\=q�U(���p��Z��L!,!⮋c�qukE��r\ΤT�<]��b2&6˹��!hsh\mʸ{y��2j�Vu������C�Нֺ�0���p���\�̯��2@dJ��������4�¼�5"��W$��*k�f�(g�X��d]i�$��Cg�7Nz?� ���
�F(��b4 �?5N� gA�YRU~�I��O�I�B��ˈ����Ŧ��B�$�	��8��t�c
j��ωZ��7�S⺭G���Ƿ�2� �"{��ʰ�9UG�C�SD�+|��^�돍��I��#�[e��u&`�G���P)�8d���z�v,�ɑUA脑$X:���1Wr�� Q�o����j.�����9[=�7��`�ʺA7#s�o�J_`�����|oɍ���B�#f,!����l8 ��}�KQKG��Z:�i��.�~�8�������`W�.J����N������~�n�A~��2�kj�(5z���i��I�V�p�<�b��#<3�X-ˋa�o	�\
\��WB�a���Y���X����
*��5~j�տ^���܊�6h?q�)�R�#9��P[,{RF&�����Y������}�a�X�l�}E�oB�ڀj ����a�ƫg�푽&��в:R�L��7`w�/�-�tM�3�/���#����Ҽx���	Tg�J�\mSO�Saxx�I/6��y	���?������9�R� ��-X��Tt-�$CD��`�=m���}�Ze�S��T�l�-h3�5�Syk��In+=hYBgI�t��u�P%[p:Œ�Jm��HaLͻ�O��3h|;��/�*�����x���8(�:gx�7�L�$nP��pL'B�A�R��&w<4���f�ɑ�,���Q2elbL�[ҝ6x^؉7��J+4�]��dboT���q#��$��pɚM{��4��2k�Y�%P/a.c�Vܼ/9�0�+_"E���d�����B�T���iO!�1�m*�Gj�n�"�������x��Dю�W�*��,�߉
ѲoV1t� �P�s�hzu��b�O�
�����p�������	�
:׌�>�K�Iz�$�0��� ���QQۂam�,�	��,�&:�	��4��O��[���Q�[9an,AG�
�
����a�~G�kL�����׃%!?uȄs~�I��
x܎��22m�^���mZH�rz�i"��2.h��P���.G��]����I�an�������ޖiO����3��厭!�w��K�!0%���YJe�[�	\c� |�wZ�F���!���m�|�k����#TV]�S�����X/`�R���ƞ��6�{����dll	��y:Mƙ	����$��L9�� �y����ڏJ�)~_�i��/d0�'�QQ�zu��I,K�ʐ�� �� �ȫC,�#(b�.��IJJN�C4�(i2�D�6����>�0�����{KI4}@�k�4���]P4�(��`<\��K�ސ��d,�F�%�Ճ�81�r��A�Ug������/���t����vØ�@�uy�%# '�3��=���~�(����F�)(�� ����&O4��/���ϳ}��s��YT���K��\;��o�th���3gVR�ݴ�����S�N�˼�K�*��R�ߐ�VB�*���&q���)N�ZW^ׁ�j���S
p��C!��0�Np�F�&@Rti�z�s5=Z��<pP@��5�j�X��"�����س����R��h��ԍ�"V�;�M;(�_�2��b�@�KY	�$ae��m�a�Ė�,�@���V���s���ô��� z���e���X#y�}X����lŀ߬���&�g�g ���n&6sz��-{���|Mn;���q��]��%�8Z�u���=��4>���9
��u���_��5�&��4�R�1i�b�Kx�$bC	����Zm���ߖ��Y>i���^��t)2]��`u��w;n(��w��9�Ak��Jc,��+e9k��~;ͬ*.!X��w%n� L���XְY���d�Qc�\լyfA-A;O�薍��۠�V$Yò|W^ ������ �f��/��S�l~H�Pr���NU��&�<���}�F���o��b	�wݺ�Vzt�Ơ�C�)�k�o����"4��$[�B}��G<&S��r��m^	(g�/x��4P�����\rМr0*6��\H	�r�R��@'�,��h��u^��єL��V1��=-��4�h�O�Z)�<^=B,�^�&%S��������$�ʖ�gv���=C���y�[�`�8, (;�����d�
��P�p�X>X0����	I1e�#9	��Y�|YRh�ڥ4P�H�y�c����;Z���R�j�fٔ2�wr#OR�S��<Uۧ�*�3zU�&��i�b��5�n `�$Ӷ�r��vdg�3U��D2_�`��f�T'�������� �t;��J����qNڧp�O���X*��PJ=ߴ?\YUb�'�����vqѓ�dG 1�a���_n�PQ)Kp|�� Ƽ�g�3�N�('䨃��;����Ō ����c����S|�����=,���}�@��EP���o���H+>"|W̭�H��E�J:�O��oQ�*M�u���tBދ����P�?��~h۴ �rqŒ�M�%���0����}n�_����̹�*����,ۂ4T�Ũ�z�|�dM���N�Py�PX��,ܭR̗�b n�O?I�C�
��M���(�ӏ�L��oh�:Ֆ3x"j��0'Q�bg������)h�e~�N2&�E1"�V���\��y+Y��c�B�/����͟~~&�?:���uw�YL*HM�.���t���܁V}b��I���b��#�$}�\���S�qwGVQ�3:L����hת+�* ��О*ߤ�s�q�4��k˜��zVuRݚv��4���c��N;�>��ja͚�9nȓ���B�D��k	�49q�9�z�j���Nj��k�_�
���������l���̻��e�An&e�����j��`�\�o�e�)J'f����)��sWs;���gu)��b���T����B�0i�j[�-�!CGX]'��I�� /7ݜ�c2����o�X��И�gNI�^�����E1��}�-��8$e-
�� e#E3W$�Q�*o@��w0�}%[j�P��?�W��Bb�A�it�*K���,Ir��L��"���X`��ހ��\۱�au�W1��ݻp��F�3���s�ƺ����y����?�݃-�F\���~�V�i�}�����.p���B��RԔ�G�t��E�p����R-�'�P���G�8HHl��'��w08��9*?vOq��}�:��V�+��B���f,����=l%%��;[��:�u�Q<�cDժ\�6��]å�M0��[}���O����i���#,��;��i��1U��o"2�ao���Y�n%q�z`�����Ȳ۔k��{�M��>ʪ���{�9�?��Ӱt,%w�H��d��?/^7y����kt�[	ZNu���E����U�I�{�O"A
��`E�s��'xJT��g�џHű��m[AS��;X�	T����ik�� �����c�W';� �S\Do�A��=��Qi���'���V[{Dߎ��^Tn���X�j�tv���#��	��:��Q~(\e�4��Sā�m�, ����&�C���$�ц�x�MR�^����>�B�W�QM;�.Ͱݬ�j�7_&����T,�X����*,*ՊV}���Gn�������O�y�U�B5�ko��)��7+�x��$)�G���_V)�Fc��ᚸ4TJ� (ċﰪ���[��0���q
s5�&[������H��0^;���l�_��f�C�?�6�L���5Os���� ��ء�x2��3J��R� ��u�fG̉ݪP4yQ�OF�����ukP.��G̶��]WU�!�+���k0�w��Bd>& 1C�E��d����u��%DX�� �L(|? �����y�����J������V+t�I�f%�ϫ����Kn�l�?U:�U��A3S�y�;��AK����a�CSpE��ʊ�&�O:���a����/�6���J�j�B9ݕ"vM	��Oҵ�0jp=��g%?���8��E���f�{���y��5����|�E��r��&I��~��uw��P�_�CtH),��o7b?���r�;�L��T��/D��;�f�c��Z���^R�wݖK��#�i��V��̰�����D���{h^Z"��$�͚%>���K������e�S�f���㻓�[��,������\ۼXVE��/��+ʬJ�U�.�?+�����x5n[��}�2��iR�R���}}�{9���Z��j@�Ao��m[����,��H�gw�,� "�[����t~�﫥�p���RDb`+���K�X|8+f��lQ��Rб�Cf~0h_�ք+��y#�-�G�#?܆��f���Uw�|�8�Ո>�'�L>���D)NzC��q�
���=�8T=������~ltr����Է<�~��1�X�Z���`��f�OϽl��� �+u@:��D���YG���&�兦������9�c-8�{�"@+�R��̈}+
�l��F���t?���PI0�k�p*�&��y�s`S �V!̬z �^U�k<�e��.�V2!*���A���<����f$̀��d�&ߵ{{�J���i��� �>���^|�WD�T$;�ə�L���
����Bn������x�F�7��x��z[C|�����`�P����1��"Y]� ��]t� �VdY���/:��+u��; Ѭ)����#���#�������e ��Sh���Z�:�#�M�g�T�ɫǾ`&sk8(#y�>�58�	��	�M�i����e�_�%�BZ���⟚��N���4�I��pj�C�}3���?6~���M�FD\`a�H�nӽIj�:�(�0��t!c�! ��
C%l��[f�v�6���ʮ[��$,F��mk%?d��/���l���D��^�)��h�*�銤@;4��!2&�b{/%�O�JȲi!���q��̗�����eڱ_��,��t�����+C�R���ڻ\�4�9��@D���?��B�Po��	��vK�
�,��� ���H��ћv�<�%��H*���>H�=|��L��ƨ�^1w��5 fM��72�,�����>�τ��=��C �}'�U�k�O�b�/�/���z��i �Y��v�0�������)�g�s��<F���>J՚�_4�z@��!��\��>�	���N�
��7�B��~�1�����'O>�OUTX9Gfazm��}Z��rGw���j��H��tp՘��0G3���LZ<J|�l]�\�/��qw#G$Թn��e�j[��Z=��/�'��ۚB�4�qOՍGT��JP' J��`B��tO8��p.��*L֎�`�_t����� M�4���B�Ia����z�`��-%1�8��Aa�j�3��W1RTZ� Jz��K�\_M�{����7�n[��R�VKdR#nO�Q�bg��Ls�T�����:�qds*�z=��VAϩ���xz�#��kt ������Z_(��s}� ?�7�%Z��hU����X�G��������~Voaō>��F���]�.$����5��(kA��z�;��}��'o���.�%|���M���5k��
]X�b.-�\��#���{@���-�^ᦶ�sh����`S��ؚQF�<��*�Xqi��h5�[�����7���߲ZM ��S��d�T<h���w�����$�6�w횂�s�$O�AC��m~'VN��uR��0�?�ǭ��{����Υ6:O�o��dQ`��5�㥙�2�5jd%`m5O*�IJ�]���5���+�a�uy7-���M�/,u����'��_�47'O�ll
4]T�,�V��7u�ݦYtמ�tJ�*��Ie��<����Ӓ�l���P�1�������lzMN�zY�\�;@�� �)��x
���n�شRDA��<u���k�=�P�7z�x��s'���_P�@]h!p���N��*�vG��]T�;o/�C��?�S�)#X���@�C4:��� l ����l 4�%�.&�Μ< o��n��H裧%lP ��2Y��:-ehF�d��}��c��o����3<����[�t��'���W���a���%F�%WDw�z�CO�����In�˝�!8��t������1�;m��I`�N�qb�V_�R���&��WvWU9PD���tS��sȮ圓MS��2�u�wS{�S4��0��O���d�&�6����l�IV���gU�՘�=v�b�O(m�bM�R�1`WWS�.._uD���<m��jnCg�u>1E(�a���zhj��X@a���́����.P��~2���7cL���pS,�Y��5\>2�?�m�,����ۑ/�b=�z ��>GmC3*�'FU�2�mb���o.ɖԺ��4��-�������ʉ�z0*��HS��=�� ܽ��/IreH�Q��2�\��0l��F�V�u�Ik.�I�o
�k\��>��� *e��o��"�u�%!"��e�!O�?�_BL�� *�DA����@]�+/�jH��D���	K�=|Ǎ��o@*h�w;���=�\��/=U �$.��Q?>���H���2�����.��І֐(i'����eM�Ik់�o���Z﮸:��V����нi]D��n��ܳ�jK����^���5;�#���Ϝ_��~�zS/����?!S��cR�rs�'�d@����l���ĭ�%��xD���W������ K�l���Gw��:T�Q�Nj��8}��>�p�0ْt;ݓ�$�"3�|ޓڑp����{�5r�cȊ
�l��pN���h�=`0s�������Z�Ij�Y����o�Ŝ���Q�qp�wÈv��YL��m���h�gh�T0%1�"~Ks�����ցbtҷ����mE�]�w��p�_��R O�*I�6�A&��gt�#���.5Ĉ��!�鸌2<�2�CaIP>70WZ��L�gG���=g���ym,�\
��\�<�%�I���`�AR�_kk�y^��C����8��#"���
�P����}f-x:|c��
�/�!(9�F�TL�jsd�߱�b�7�5�N��6J3N찦�K @.:�j�P��ީ? B��e����1z�(��
"�)�������c���+f�CWXbW��$jr�j�y*q�L8��fMg\��tܞ�yu��Yb����mX��
�.W�p�*��91����WfR�LR���d���TY��mU��* S��q���E��T�(A��V
��/O�Xj����5�T
�[z�w8FֵqOt#����p)I���Q�uf-I��<�5Oڹ)^=���*Z�H�	y�5��ə����'�Nn�.��>E0Ra2Sh�vN( ��Q�����/*MmB�l":�0��k�-T����~��㓴z� fft�k�FZ�
�Q������5ц��H��\���X
h��K
)�w�t��S�����+F`^�m��1 �k���e�L)�6f����"h��nT��l��/�ޠU�z:��d��T��Y�YUG�g����l��s�x).ms�Z�N`辢�- �uWt�q�-���5]�{jD��b�:p�K/�[�!$`��{���٪/6�e���Ʒt(j�(���-�x��b�Wݏ�)/g�w����疽[�A'm�iA�U���88�7�7Z�i���'����9�5�K.]�N��`s���r�ύ�4�Tb�0�v3$����M�ݙQTI�T�������۩,mùCD��1N��XTa]xt�'��1�Mӄ^���&~Gi��X���PYt.y^�x�t+��Au �]:��ںJ��vŐ�^!3m�]m�u�ZU[��?Z���=�0;�;e�j�?k'J��Z���n
�M� 5��Z�;��c���">�aPx`��nU�U�|���'���e�U���D�-�n��J�
�a���1��rr�H�t�����	a��z��� �N�!��M�yGU�9�þ�e��$g�vU���U�P �j��ѻ{�{��V9����sP�> $0�Z��+-�'ox�\��5��7°��%�)#l���{-	+���R�i�J�|����7�}��o ��o�P⥁c
Ъ"�uN��^��Q5�z�y'� �{U����ǣg^&~'Z�M�c�-DqA=�1�g�_�H�W�`)�S�n�#���J\ʚ9V�gЯ1
�/W�x�[C1��`�H��#���m�R���0�A#$$�<co�^l��v�wQ����M1e�{U��+���9���'S��d�J#`��A�4�R	Ɣ!��?�JՅ�7�+�^�M�k<��_4�أ򝯠л��:�EL�y~b���.����P���S����n��,���p��.e,&˻�����U�lK�c���VO�g�߫�;b����zAf�0��Ϡ����u4��τ+!h�8[OJ���F*b��?!���縧Z̄�h;o&~f�_"�= ��(����^���ݾ�������`�썊]���1���
�Pߺ��)�P���\�}����(Z)���{}
�"aV�8�¶���]��U�oW,�Q�Ȗ��fdeG֣�%!c�'z��H+JHt��O%;��95n�\hՃ�|m���dg��y�h����.��%ER{j�vǀ���S�y�Z��]�WCp2i�bA�	�%i\腝��5���z�hHI����x�kH�A{�IA 11��J�ػ�/` s����Wl$�O�Q�0��fOj8SsQpM�����c������@����?Q2]<�;s;��k��opI�xٲ�m�~��A�>O�D�xU���*!��nr�A^�^1"7)Y�}ӟu�l�o��ai����qo*	6\�p/��[��4F�bI�\|�ۛQ��A���s�U�V��i@�#�2i�e� ,��e���_�����]c�)�$O�,��(Tr�G�7L�#6�, �*�0�~3z��`���^�t��f�k4�����J�j�?��B8"��Q��
f����n(�E��G�P�.�7������{��-j"{�	]��!��E~��dW�&�~l�zЌ���݄��w�w����A��c�Ǯ!'��,+���c�����F�sp�Y#G�Y=o�Mw���+�yz;}2�3��抩g>�� `� (�|�Z������%�l0i8��>�̆OYl�ʃ5�̚��A����=���U-� �z/��eTJ1�E��@©�����p�����
�L���Y��M��� #?��_������0j$l��I{��vB5�z#j$4�G���0@�Y{e'aX*�-�V�p�U����f{��Z|���5Z36��؏?�,�t_��B�GT��Q
*�i��4����]_7<�ds��lL=%��x�vb�����3#��mA]J!��[ꘓ��뻟"xg��x:7G�w?E���O|��z�"�p����4g�>�EvA_MA��7�`��I��{� ��!"mU��y�����bKhH��6�3�D���y��8q̎�DJi��ٌ^�k���*'/�3t�B뛝�����J���)=89t��r�s�#^g�7��Uo�~۾�D����F-ѐCޝW��X=�M�vS�nY�h���JK�,L_��!Pm9���q;V;{,�ѝ�����/����l�*tB�|���fy.�sQvι�����T�Z���]2Ĭ|Ͼ�A�X5:i�E
xv
v�V������B�</��g"=��ա�X�7܉�s��a�A��o:����z���}k�t3�K$, �yau	r���9mh�*���V]� _~@5��OO[���Y�RuKo>
�k^n�����(��M��(P�'����쵙߮bcN�T6l<VyUJ�p��3��ew�޾^EŜ�����s���].)����Ox�
2 �2R(�N[~B�`A���h"��Bi<&i(��x��/�|�9?�3�5�/!|A�5�-�F�OD�:{��r����8zlDm��o�]���AN�S�`�3{n��1O��� �x��-��p���Pw�9
:6T{�}ҳb<�m\a�pa��Ǆ������|A�m�(�Q��n���;ś�-��T��3@q���a���,m)|��A����\d��G���- ����\��Ff�߈�\ұ�M��.g�,#�á�c�(�'������u�AK�hS�_�J�����2q a��;P7��y�z���C�'ak߭��);hGAC9QRp�NYd��=��i�����b���</���Z�(Ү�� (�1N�'��Ik&}��d&YPio��jjL����."����	��-V6��!��8�t{�dr��c��m1ZM+�+@<4?c�����&�2�����"��8d�G�$�5��-�{��N� ��f]�rk�� ֱ��am�S� ��/�M�M,�2��t's�p�9IfƣǴ�+�L �C3�����q!�iz���;�l*
���3��A*��x��_��m� 3�H!#O}KE�2�M�]'E�q�Tqq���7d�~Y=�w~@2����Ҝ��� W��4��9�*���ן��{��S���q��Pñ�S����nv�����(Nu���,7(y���A�� PEű��#�_�,�M��?5��oC5p]D~������S3tA\�C]�<f�_W;0�K61rW�[_a}+h ��q#ӣs'��Y�6^X�@��t��g�J�ޗU�<���|��̥�V�JI�_ -�Ne��vq&�s9t�� �/��k��@Cǌ1{�LM��/�=�k���b�c]�Հ\�.۱h�v��B�PH���*X�.���0�0���jB��K3��,�1�{EY@��Th�坖�DE��k*6�uub��4��L㠝uZJ2�B�z�K�<�$�Q�$W�����lb�C���3�1*RZ���٣^�����e�J���>�t�}M�ثM���-�j�iP�B���z ���������;i���D����b�ɞ\�,u#��7���p~��Μ�
����֮����kʁ;B�-`V��H�f��&$~�+Kw�5+3��u*��X���
�i�֭���@�\8
"҈���!A�R��"bͩ�3#�U�W�;
R"ט����i���W' Z0A?v���=�<�eK%���'\*uO������#��F��
ˉ]�NfT6%��"�.���Ÿ�ԭ0|�/_وi �3 ����6pnkvQ��\H=�n:�nܗ��q<�d�m��»�cz��nJ4�0:![X8�k]>E�D�U��-1��b�ڇ������~K�Hƀ�=F$�S9��U���Ð�"�`�e�������aR��	&��VĜ����&ӊ7<����H�3�)I������g(
���asq�+�D:�{Lс�-�z-��/<J�`���(U�y�f���i6
�� ]�4͇��>�A1%p`2%K0J�FQ>ڧ�G�H�8�5��t��>y�U?:7u���7U��9թL�8ZAn�c�d3����}w��+u���*���T�7�E���8}|�&X��f��M�,�F��F���G6���fn��V����<�#30l����M�	�X�#!)�+nZ�� ƶ@X���Q`����[�HI'����:��ڈlf��F�|1�'���GL'�U/���N#8V~��?kD*�r�l��S�;_�]���uf��D�h+�?ޡ����"*ʬq�_��+���O��z#�o�@�����BfK`����ȴF��U�q� �pCl�G���Z��aq��v���r%B�"��>����Bx���]Z��҇�뱚�/��h�(i4]�q��>�v������IO.J�P.�f�b�U�j�`����l�ݝ�G�/���LY=t�<�e�@�@R7��+��ҭ���C8e����� �$?"�<�������	?X^V��O����"�H�$Yٍ}9���iRr�l�yݓFr�Xvw)x&�MYfvot=c��j`:�(-�Ɯ ���U_��-pI�����x~�X���}��V��o���TE�S��0*���0�+�k&��Z���I|1Ƣ��F�3�E�*���]9���Hs���.@<6AL�ap���P���b��[��y�����$���H��?��D"�N��%!��؅���K��D��c����Ωv2c�ZY|�N�U��,��P���3�i�%䰱Md+N�p$m6���rkCp��3J%�V�!_�|N�g�Y$d:e��"����{P@��:�+���}��.�ĉP�9P{���欫3��>`.�a	�58��>W��M�)=#��9�1�QJ{^l"T�:��p!-�*g6$>c.�ɳK�FMfJRY>������i�* ����*��� D�뀐!2���/�pr����<A� �vr����ղ�����\�a���'A��i�Š�0���RV��kT�d���0�,}�i7��x�� ��]�Lz*��28����{x�Z�(�ۑYMkJ��0�H��{�[�����E��f�L+�.���-���n���%������(�ܾ&z���Q��JT�8X~]�ԁ)�[vw5Z	��ZPW��("�j.��.��C�o�Z"�`���Pt��_2�Izl���B7+��&�g��'�>B`� Ǟ��?�HY����m$֋%�sD����Bc��&4��w]ЈK���:6Ө�Z�pz��=����uڐƬԴ�zv�bʸ�aR$ii����?M�ɳ����G����۷?����A����1��x��?ʾ��4���Q����TH�"Q�D�f�&���A�g�}�}���O�˳��É���Sr�ڊԶK�.�t���iE��֕W����>~�����uՊX̥B��tt����"���~lS��9(ryC��~�����pO׋M8�&Œ'��T����n_���"4K�6�q���v�ܾ5���H�R����jq�Cg�g�f� }���2�AW᠘;��L;T�����=j`�����W��䑩��	x|��r�3t�yn���A�dv�X~��b(+4��a����>Ud�ko���K�� �Zw--Xf����t��&���H�L9NӒ\l�yKl��hA2M~?��������p��E0 �$bq[�H���OGUn�-{�5lj��Ev���]�*#F`gq�:ҍ[
�;W��<L&���j*#�6�̞!s�W�
"��_n��V�����B��Y�����+�F��'�4���fc3#�����ћHU��y�c�ˮih�<6�FX�	z�@$_�����OuY��!!������f���%y�r��s ]9��Н��8�v̄:Lv��#���n[��2ntT)C BZz�j.~x!1=z��4��[3�"7�i?�Y��o��g�J�B��vA��^
��I['�$m���8@~�wY	_�ʧ\Sx�`�8������_a��C{��H��:ka���|̄����\��s)(Q⦙0�$T��:��ڬϸO��a�B�Z8G���J�=({\,�!�Q�9��Gᢾ���w���0�7��=浼B��瘎��`m/�!��O��=\癈v@̈́�
�}�t���(�c!� =p�MB�%�ɴ������,˸H��&��*�^t�Z�K�Q0��N��|#�֔�¹�A��Q�oQ��SPz�+�ޱ�,4�����E_�1v�7
���G�o��ED�Zr#և�XN�,9Y3�a��L���&��u�y����,��ҍgB�vݧ_�t2���3�h5�j�Jf~V��� j�ORyg=��[�&z������lX8�x*���Ep�J8�n�-3�8%��ެ�▅�Z���\G@��1PX�P��*�8�t��z_���/蠾�w�S���W��8k(nO`f���i��j��a}�-��k�|�D��pu�<�=qd�K�e��c�%"�}˓���������-�	t�X���*#*4O�N#��f��F���r��"YҞU����ymГ�2t<��Ӗc�CQ+
��)�k�l5�Րmɩ��OT�?����͜����4��D�7�)�L1Ҿf�ۛ�(�������En*;�T�sT|[u��E!ԲBU+x��`�&)^\� �:��!��Ȏn�!�J�)@�D��E��>��4+��ɐ�m#<��J gX-HK[������������(����Q�DG�ˢ��o�����ϑ�R���}X#�$>����bJ�azǅ���x"�@y`9�Lӷ�c����j�������/ھX,X�S��Svۚ2��n�TVFX4��~�F��޺�NAP��q�frE��0���/��x�����O���Z�i ���Y@�X�\�eW;�ŋT��c�j�=��<2���@۵�y�<R̝�7��w�`1��:o��'K�8�l�]��e>ơXL;�ض���)9�����!1ɻx6ɫ;�"���bޏ�E3���!Yn�n�/ѽ�M�H��= Mq�1�)�Kj8V���\~!�U���b&}����+��#k�ɤт�2w�b#����P�è������[cy^�V("�IQ3�q��1`yU2�����+Mnh��?�y+UL��a'�a�)�»;��P>͒wx���6ur,��"��A&PU�vψ�<�2�FTc��Ż�+�ߐ�&����vTNxṢ�Yƻ���2�6����7P�I�h�0��s���h�?�-���n�VQ�@l7	̃�^.Ka2u�����U�m#�0����8�E��d�����I�z��dn�t��n354�RtO��A�ݞ�&Y�h�m�mu���=Fc��[Z�aUu���Vb��~��a�%���Oo�,ɽ�S�L�D�`�o{ �(��zpz˲x�P�n�[�_��:!tXQp*-��e�v�>����$H>Άx>Gϓzb���5�1*��W`�;Уů���պ��4%��NtY��B��x�!2j�[��N<O}	G��_#�0�j-����3�O޿�n�~k�5��W�4�ve�3�f�a�ҋ��h�P�yfM=<����gM>�J�����`i�XOw�qtކ,!�t�*g[RhΞiO�1u��6nK��#�a�9Y���V5x���3yj��`~��N�/�jMkjXh�lř9��r��,f�&;�m�G3䙛��%�m�@'㋻�r�F�*n#1�����%�602δB0 t2B��OѸ��z�)ތ=ˈ?���~��]�:v������8�,fF�Cx��gz_�6�4�s�,��Hz�!���(��~˺[y"�@�k�gD^ղMrU�����c�k֕2��������D
w��x���H�8�\��Q!�*��A}�Q��Xŕ9��'}=x�NB�, s��q�9�� ����x��½kV�w4$�>�>
��Q6�(���^�+z�������aƸ�M���qgGw�M�@�Wg&F�qt&����.�����2�-l���X��0-����Va�\¹#y�#��<Gu��ٲ��5���ȝb<��i�	g�f���l���e�����ܭ�P$��]�C�?W�s��"��,uy󷫶0NS��-Ax�`Y�[�m�ֽ�m�W�������l$T�|4z�vs^����k�AD�.��C��:��mX��joS����@nR�'�/8
	h�T�㍜�r���[j��[�lh�i�֟�2�5���Z���젓!ٜ�6�Kn}|-�'������rwz�F7����W_�h�x��VA�_./�,��_�������e�:i%%$�>-u���-/�F�V�����Xeˍ�g�(Q��,:ث�9�Řsw�\k����1�d4,Ó,��)�adjZ:�3t�v͋Z�2���ᚧrJ��ZXry_����R�CA/���1��e�q-dP�ؑ����t&�C�HY,-�g6B�)-�%"�tٵl4�5"d�h(W���O��L})Z�-_�P���S��Vk?���R��hsLh�D�B@t��4��	q
r����c"��ĥ�s��8/>2a
}x }�
�I�5B��0��	.����Ȟ f�e�M�D�?
~��@�f���w��x<^b�����?D��*�5�a8a�$)T�_&Y$�s���iUB�G/XAg+,Z�i��槯����=���Ly��QȀ�!v�@aC�O�_�����B�9��N���y�u�z����e�"�Od�*��c�3HM��ǲC"m~ ���T	��s��bdH����d�JK�lb��λ�W��'@�x�����aQ�a|�wP��n�����d�X>?�=a1�s��x�(��*��YC��/*"��#�	��n��RG��=]��o�*����6��s�&*�Q���%zNwʯ4Z|@��GU\�G��q<`#�z��ѡ����,?H�R��{��b�͏�&�nk�5 ����o�j��ʑ��ܓPF+�/��>�_`��J�9�7�)q�����H�Z34�!�l@��z�d��3"�������,bYv�9���S���R���Kh����&�D�ˢ+G	,�#�'T���79�s�<�6�($�aF�"(��P*��"q0?�����	(��Wgn�St�������K ����L{?i7Lp�B��1U�4(��]��ɩ�;z�����c9�O��;���b7W���/wl�iNT;b�
���C�OAš��Xw������g���FL���r���X�k�����������7���g!��e�<�J�6���&���m����wiD���ֳ�/E4*�������?o$�����17�9o��X� 6߼Bɾ��� �|�b�<E���� �U9X��Y(J�'g�$� _�;�G}�g2�<ru�����`� �(�V\��?5��,n�1S]g?�A��8��"���{|��-Uy��1ȩ��?b�>�HLK�{�x��M���ӓ+��f��MҊ��C�Z�w�O[�M����3[M���W���t��TM5/͔�3eiEP���ట�T�c0�Q��;BoE7wl��_ϐ�l�<I�_ˣ��y^ǳ�g���@b�K�*�^1��R\�L�-{��V�y�-R,�m��������GB�)�(%s�p�D�t�f�ڰo=1e��A�~�:�ޮ�d����{l	��ѻ@ ʘ��xa�;[�?��K��c�j�#^���A
{���>A^�,�{��b���%C'����0j��z9x�"�1��y���ųJ����k[ -i�-��� �Lvo���T����G7��'���D"�C&lߔ(T�=�_t}���y?��iOb�gh�5@@1.<��l�I����^�*�t����I���{�w�Z�o?�����
wԥ��뤲2�_��C`=��]�\K(T�pk��x���Nw2{7�us�oo�t�,0��N��49�P,9�j?��,�|�t����+���r%E��+l���i��%<�*�>;���sg��{l�g��l�xr�tv�m��|�\l� �XT�ۘC7#䪓>��O�9��.�� ��*�����H��^i$Z���	,p�����i��cyY�y=�۸��b�3ug��N<bs�1����^�"j9t.5�u�˓jMjܱm��M5��`�d/��n�N3�q�:.�Vl���Stuv9Fj|��i4���<kCs9_I�����s��k�T��NR��6w��*U�<�z��-k9��De�6#�AX�[9'����%};�aQ�c��������#GW�Hk��Y��DD�˷��`C�!�8�Iw��lB�DR+^��۷u�j����VҌ��lCE	��zʞ��џ�f�
�B���gH�\��0T�����+�\D][����b �@*>�S�Y����-qoBa���m%q�/-�Y��n)o5��
�z�UxF/����gI�2Eׁ��DdQ�+l�Ip��Z��
�q��4J�Ȁ��TeMS$�i;&0D�����BQ	;o�|\'��� �a�{ϭOY@�&��䀀I�H��� �SD&�]����uu~>�����4������.cY�Wq��[� �~Z��3����ZRc�A�))��{�
�f��
*��ԠчR��Tz6�jm��y8��,�8������7�@��GI��S�gۻ�L}���l�U}��1v��
����X�M�#;���_�vs��}�v$�H��T�)��i#@5����cH(�@��n��#�o�9�$*U��IG�����/��H��'�;9��Q��Z�l��ay0�i���:	�ع��!S�ľ��|��+�Kv��ȫ����i%�v����n8�������՞�O�ļ&� ����=��U2S��X�!8��ɭFAZLu�*@xt�������Xw�a0>��?��� oEc-�]{�Q��W �"11P8�S�4HGk���P>��\z��T���tqp�5N�	��ᖅ�{σ%�$f�υm�]S�f�w45ms�˄QZE$�`�B���r�h���ы]ب+�G�l4yiP=��d��@�C�*ѣg-V� #Z����1�ºQ1�]���@��`��_��Kb?7��0ql�)Қ%F�bZAa-���,\"�H� 7w���P6��wz��Ԣ�e��7���Y74����ҨZ�ZX���-��q�6 oh�����52 �]��T-�,�,:%$ � Z�p���a���e�Wʁh��Aф���>t���>di��@�Y�[�e�����'�T-(-{��;4���:O�_���?�}�m2H�R�#�~�ιb�ۓSҶoNiH7�p�|�+k^^y{��㪞�
�ˠH���ʚ۠O�}��3h�?���w� D�m�f���(��V_>��'1:��3\JMH�}���K@�2ԛm���Z�՝WU=W�^e7R�]ؽ�c�	i�k�v�B�?�5�i��r�!��.9w������g�]�VXrF l<�a�I<V��h�-����;�ؼ6FN�`�E�(���̭��얎4�p	�a��$�e����8S�-���o�K�,�����",�p�FPT֛_��U�&x���A)~vЖ�u&���)Š>�`6���.��C�	t.Ĥ�D�����q�`UZP�ux�`�B}�o�ҩ�g��K�2�J��ă�m˓���J�d="�j
�5(��'}y/rq؛�q�3.�:F��ro�%%��ae���l���v�P(��@�$v�]�믿N}�����qR!��p������r�2 ͈�?���h;���` �++5W����j;#�*a��<_����X�O$	_7��?�c�ӱ�Q<����ӓ��L�Kj���Z0	��^�i���.-��D撿����&J�GU�Hf�H;��v��P���M0��!k�A��(%hڸ�g�u��λp�4�n7+m���n�VElF�@!6�lA=�Ok�;��XݪX��<6�EJu�����P<-�����}�x�-�^Ry�����%z{PD*R&��վaf%̮�u�(>�B\�F7��X�>��1�O�ȧ9Ow0����d��*��0Y�!�����n���=��mH���%��o@�7@x�|��!I��(4���Ƙ���k���i�.�xo@�m��ͨ�����&ŪH��S�o�r�צhۄ��Z�S�nȿ�"�^��.gUi����s���Tbw�̔��9�<^c��	��%O�xй�d�U�P{/އj��	�u�m>tU^�Ͼ��{�H��i�ݷW���������|��q�ڢ�
q�/$�-��<ն�,YǔD�6ݠ�)����Ȝ�s�n�Bzn-�"�D|�b˰��Z�:u�_�v�����Z,������c-W%������zw��v"�C��フ��ȽD��s�;Ɲ?-5��R�?��> zͳ-A��x��)"4���S�yV�;�|�:��m�!���ޜ#&��-�7��)�gк�QO#|Ԇ�W������3_X����3d�lb���%�`���l�����.|oHN@�9K��=�#�y��I���X�'�k�oJ�^�9��X��e��[������f-�"f��:�C����6����gi���G4ɀ�*�F�_�ZO �,۠� ��eF�nҰ !��HIKH��y�bk_���ʎZ	Lfn��8	0wz:K&��J2��`��CM0Vq�5~eE��MS�>����i D���mcY���\�Wv��ܝ�"5�`��/����s���r�5��-O֨���B:���:,��/R��@-G��Nw|��W �+�4�R�9�V�G����>�������2q�]�� %�?Q[���e+�4�ʸ�rV}T+��T3�>1�Kӗ	|���"Q�����xu5O�@O�"�!Wu��脱Ŝ9`,��=� �D�����7hfS���0��?"����#�ۀ&<7ٔ{Yы�Pc�Q�&:u��v(H��_X��j��I���C�tf�R�=I�_Z5A��hذ ����׍�}�?[eW����y�F�Y�AfZ�
}g�/�)D;5��{��ő�z�ϻF�`Ma�����\���k�ը��w( ���{k���f���.�=F���l�)}��%9��X�8�
#(M�,�[��3#��!o=�?,4����Z�m��9��G��2�&�?=�0��E:[A��ٔCW(J1I�)D�N����L�~�����Ls�?]I���;ڑi`�|PX��~l�����y���Y�� �M~����.��&e?�������)ރ:�TQ�IbD
U �j�\�����\��0������D�咇P�>��hZG��5����.��D.t�/�����W��g�_Öo7�zu�)i�|m���P7,�TJ�c�~�M͉�J#�%~̍�T<���+b�*�X)��2��� $-�2�c}��](���!��>�V ���1YZSV��_�Zi���bě�@�7�"�d��:c��>����\�!����3����P�����IA;��q�K8�־����A�������8�h��� �%.���>N;i2���]��"y@��RaRB�{��/C��(U���_�yq�za�Z���2��R�F��k����<��Z��a؃���N��0��I%�v=Ð1��[��_z���X�&��#�F%��7��'1��=���3$������kw׍;`��71���q�1�SQ=��*�0,a�3ӏ� �͘o�����^�nY�_E��>��m�a�v��:����ʌ˘����7`_�<��X���\�r(�+�ڱ	�(��[�!$z�.������k�����P��V�"��4���Y"��M֜���m��K�desⅈ}��6����Gcػ>͂��"�b.�E
�3iTC����y9�,M�6�N�P2x3�f�0*��:���ŰTu�Krjw�E3ߠ��ĸ���`dL�uq���~0@\���ėE���d���1&��Ɗ�c4�����ܕ�E������DD\�cِ�mQ���b�̷���F��=����h��0/���S��3|��;�I22w�"Żǀ�ժ����wo.~�P��*�S�)k�l����L �����}��^be%�]�+g�܊̄�n�O��<�5�#� >��NyEun�1��MQB1��p(�l֖���MR���7��E�ɤv�䅇��\D��p��Dn���m׫�ꆾ�X�!��/M7�$$=�j��1 ���c[YLC��Pg�$�낟�7lX��_��j-�@�,���Ą���:|9��R��ve�����|RWT�X:�Z�/B=��;j
����N���O��T��!�]�}r!Y����n�j �[-��Zr�"���]�s��if�,DW�c������sk����.�ͻxˑq��*���eI���2l"�W���8|E�g�W�Z�0�d����YئǤ(wYvLץ����ZL. 0W��s�aQL���)�>�`2[ �q�e����o�t(&m�)���(��,s�����4_���uvGYdp����꒶�%�c��ΏPb���Ŀ_'�|�X�/�?�=���V�~+���%?�JD�p;&��g� :Q+�78zfs��ϭ!8X��]�c�J����I���$(�*��H�G��!��3h�ɉ:���bWW��zO���k��@ҹ�c���ԃ��MT5R9��ò���4���o�,1�P�5��4���uQvG%�'�|n>�T�r�
��4͠���
a�_�[`6��>����O!�����"S�!~��)J�
I��%r�
x��pz���g�CW��[(]��`���cؚ�
�r4u�I�Yu�x�'GQ�e\5�N��L징)�JB��	?	8/��p=g6��ο����ws`�u��C4v��W"��0�"7���Q(Q��0��Y�Xl�v/J�-PܟlT�/�t�o�!���^w#Ĳ�=O�v.�*EK����sRL5�.� h����.7^5��s����	�=�h^K�1���n�C��(Ԋ�,����9"�<+#���	�[2�����w��m���ء���V���*y����Nj�V��ޤ1�X"B���I�ds��T1M�J��wm����U��ˊ�
�>g�M >�������N�ۃkk����tS�B$���d��?>ҍ<����F	�i�Hm���y�n�Hۍ��ˎ�#�ޚ��X�����nk�, N����V1���*�DH �	0��ӱ@F .�#� g����1�(���`T�G|HC�'>Ǉ���� ft/�g���|U��&G �8����E���r��T;k�%DJ@5J�K�<T]�������3*�������"�Q�H�R��h����+Hf=l⏧�7�ANVX'9�I��ń���{m������� Q�fl�'T�N�؜:�qh=X�3���{Њn�U�B�:1�A�e��
�}sCJ�\[|j�%��w�@��_Wc�`��,ŮC����'�Sŋw@����2�N��,��SB���da�X������#n�A?�5�u+@�e��`d��S�0p�i�R�/q;�c!���ZU��j������%~Ÿ��椒'9Y��o��-@F��G�z�*��B�_	;��Or���NHY^t*�v�6�w[	�^z�cZ�l�'�ƕ"�^��XC`��K>���_�ɼ�$`^8d3�R&��4AԒ�[��B��˲� "<U��pq���ØW�a�t�ܡ ��O~s����a���p�֌�5'G��mZEeN�b'���jƅ�#bY�aE�y�Z��N)d���������"5	��|2p<��/���Y7~]�Yw�	 *M��o2����P������y@��2�1T�#�B"Kn�N��;�i 3�SoF�]QG��c���X��S��D<��i	���G�#'5�;ղtG� /��N�F{T,X	�%�E�C;AU;������"T�m�بʋa Vt��L)c�j����`�Y��-�����/��A���:X��%�π�r��B�^�7*(��>�x Sq����(1�@Y_��=P�%2���R����YODuM6�T�^Ml�j�B�-��h���F[xD ��^-dY��f���������VZ.��anJ�<5�u+�����Cǉ ����P�Bl�KJ�72��+
rb�	l�Ӂ��D�De�"	]����M@Q���:^N� �¥��Zg��cCe_�Wn�kĚ,Mg��$$x�<��@�L���O��vz�N�����G�i����n7����PxT������n)��� �x.VE+-��x�[�����=���2JL�I�mɝZ�$.?���e��V�`m�*�W��J4���A�z�+OP�Й�>yPFH�C���-"T���2�@mx�C��"K���$�˿_>Y�Y��ϡ��<ĽW���Q��L�����Ɏ��7`��f����,����U0�-���ĺ�9�"q0�jJ�������_��Q���nxa�ih���R�*�羧6!�T�
|�U뒪���jfݡٔ=lC&N��1{�}uM���;�Ju���o�75ØS��:bG�`iȽ��F�4�^F�u#Cz*l@�����IrD����)���&M��R1ni����h�E��+	�LN�|hb=�o�T\�l�w��3
��C�UMH4]�lƍ�uh�o��ƩW3�����/IH�,�Fx:�m�TP�-'�
֖G�cSP�����w�C������<X�`���a�P�j���㠴K��^ϸ����/=8���\R���	�6�S�	]؞�E���� �F�֠o�P��t/�\�L�?�%��l���#n���ˤ�jE!d��gL]	�̧|녵�1FѠ#R�ӛ#��l�״=�^̓��d"pۍ��� U�JPu��C��dR���XI�l��g,_�N����$���+�bpk#�5�-%\�5��ĳ�|a8�Ұ�	RdK�s�|_O�$fߠK���P��m"���$��AG1�80OF��>�ȯjy�Q�u�/��(욪j$m��M��J?[!�+gap�*�7Yd�un�m_�m'���M�icvR:n�*͌50��瑷��9�ŗZ����Ą�YD��0�[Lo���{�9X����0:���o�my�Qa*
�=����z�Ɉ��F��]�a\�����.�h�@9�]�d"������Gي�mZ�Q�V�m`C�Kk�X7/B�H�6�gG�73�9�������(Z3�s):�c�0OLi�6! ���JS"{��l9�*�5u���њr+[�vӓ��W3��Y����.SҎ!�cA�Epc��L,�/ �����!VXR2��J*�V�jI_�uT�aNN�V']W4j_��f���_�9I�(�|P���Hi���6�R�/��٬MHQ�ks��G�zߌ�@�����:T�}�i��,����ǟ���J��J��E�ر��_-C5 "��
��㬣(dTNع·ə;��E8f�BwBf9���P^�k�Z�x��]��~��8���V8׻�sS?nv�@�Z�^��OkF�Ob$��̄�)è+�U9��,�6R��s�[�V�1: [@��^�Q�IP����U�Q��Q�O^�b
�JD����X��Iq5�6c"�����Ff��[��P���70E�Z|��aDP����Z@�C���>E�
�l�yX��Ο3�B-g��GH��L���/z�H��,T�%�y1�t�� �	�Nz�7hD�8�9�Oh�_$���5�����#r�^��FS];�f��%�9��ߙ̪_��GF���X��e�a�9��,�:3M���+*�8e�u� ��ż��Č"��tV�I������˥��_	_�]n6���~P^�� EA���v��D�H�c������:��ƍg~Yz�|e^z+�q�����yi���q�{��hsytC<����N(��8:�L��ۙ�'�-���z3J�`:�S��_!�kV9ϥ\�W�$�\T��$WƼ�$aUƆT�g��������0�$?���v�$xF�n�8k��-V�bwa8hpV�����b�2��>���8���6<A���EvDg:eb([1�Q��x+�����l�*&m�m}�:��cC����(˫�՗p��<!Y������Ii���P�Y�:��S��"w9}6���f5�u���ȕ��v�}:B�X�D����do�/�����CB+p^�bn�Y��W�;� i-wȃ��с���Q00���?���7�V�PXނ��N��A�bk21(���0�ѻ��^#��<X��R�ȟ�D��o�:�*\Q������*x9##̒Ɠf4�ú��ҫbf_Wo/�\WӲ���jl;�x��]s1zWw�^���,��Z T}hk|�\�N��3��
r������q�5Y#���3��&r]kmGvZ���)T?,n��@l���'E
��=
bk0����M���
�/�{�)���������Mp����뱉�8n���T�����u�C&�ƣ��;υ	]�w��:����F�y�a����*�b�!�tvx@}������VT��~x���\�FZ���IK���[dTG�碍]{X�yp��R����$�Z+!TM&`'��0����e������{g3�ǥ�� 4��FΚ�p{>f�_�L(h<ɶ�g˶<�v:�g��g�R���o�< �#ƪ��<+�����D�͞�9s��{��f�9^wNJ�V��|���'Z��l
W��W��S����\NKN�����L�w'�݌�	�I��V�[t�s�\.�i2�A뽠/IOy�c��p;�I6 &G
�[qf|%�	r_lB���)�H�}mBu]a5��o�_ڴd��*kߗ'�jB5������ٛ���'#�/Ŋ��{Tnk�
S��kE�2maK��F�r�RR�Ճd���+{��6-�zD��BGGe��(��0R���D���:�A�D��4u�
V���_=I�Ou�����=D�
�ڄx�<Sa
bXa�����F���V�zd���K�q[H��v` x�7J���Χ�uv#\�Gh5�ۚ
EM:hC��Pg�s������� K��Oxu��/f�F�w;xˠu���lK����gc֣\@�|1xI�$ Y��/�=���B��u�X��AI2"�������e��Ve���g|���1,�K�ȩ����0�s¶,ٽ���-���@��)G��޵`w"��	Ӗ��O���&��R���l��s:� �����C�eʇ��#e;��ϭ��ND�����ؚT�X�=�zӌ���L�+ܘ�Y}k��oJz��`�L��s�
7��%\?�@������ar��;N���5
�k�5���#/{�keB����ZR��J�-?[N����M1�|{~1e���5w�^2�u}6����g5D�h�����,�>c>>� �V� 	n�&�|L�z��w�ˋ�/�\,K��ˌ,���϶i�`,}�V#�&1�� 'F�y�� ���}�W�����9 ��o�J��g&aȿ#������)�[�����i ��,�B����2q��_J��h�3�x�W��X�]��G�h9�@���:`�Po@����\V�LE��g:��o4�N~>�������I²�*0c��u����gӲ�E�C���W,Nj+
�3^¼����j�:����ع��HC�b�����P�ۅ�&��0�뜮�B�ɦ���Or0s�'qH�߮���ĸ�y�-�@\�t�r�)�c1�^�9���$Y�S	�g��g����FT!�*����>U�L�v�(b�Z�+�v87�^<`V���&?��B;Q��?�z��w�@��c>ׁ�<mwG��o�s{l�{�|PA���a�d�剑��Ykң���+�� ��Z�{N�_.��ؙ�sS�{jN[
�I�N���Sl�����8�)�e�I/����4�}W�<�\�O����;Ӱ���f��L�%SKm�E9h��a�u=��u��"�ǜ�{=p ��=T�hȴ�i�2�&�Ly�Ro���z�E�V�����D>��E^���׊�JJ�-�#�]/�R՜��9�<A#�����38/��_7J���bՐn�f��A�z!K�5KQ��俐SB4�T5���V�{�x������|��Kj_҃��e ��g�~�(B�&��ֿ}����g 54a�"��2kGWא�ҿ�p��NqSW�w*��][Y�%�	r���U�{�urm[t��t&�X5U�n?nqL5;v��^��e�nl�)T=���l�=@�u�gw��T	��T�L�y�e>�0���)$m�!��������
"%�>S>�&>���_+-KLq��ƝAӼ9���I<���:���h6;���X���;���D��iZ�l�����:ȗ���d!��,�O�{���_N��F����Ix�1��c�Rݠp1�qc�/z�:�,*,�i�9�X��-��m(JCW���7���̢���C�[��ǣ^����$��?�Η|  ���H�G`ݵl�f��*^yK��Б��m�7ͬ4�Tl��CZ�G���Wa�_���*XGE�bT9r���.s��Ą�������ڛ�u��opE,��nS3�|��a:�늖xs'�[���ܑ��;�1�aM��Ɓ,�w˲#��f&&��fs�g��͘�h�d\.�k �tz(-�q�8������M�,Ʃ�I1j3
R�LIl���Ty����Q���b�_���%��/R�����Ew)-"�&uE�x�f�����'�Јמ0d�s�oW�R��S�?(azX�����@����_~���5����N�r~���j����VHI��+��KP�K��$C�����i��䏉yxWp�_�	�/@g�9]�y��:6���� �vS��&�$'��ֺ}��I �S�n�_*��/C�O+��{��+�4�ټ���rbo@�; #ԑՒ}��_��j�N�j�y���]Q�l:]/�<Y:x6�����	�N� b��۾>��7&�W���.�|�7z��/�V�- ʶp7��1Ea:7C�;~�o�ym�t�`�ilz �Xҥ����įqҍ��ƍ=�W[(|��Y�B���U��-��  �懬�
�8�|�JdJ���bE�Ts���DM�T�������;�嫂�ݯ�Y�Pq{�\Ba��)�`�:����^�R�rO�ʟL=�d�t񹓀"��l�ǭ�w��%��#�3�����sYM|YC�2�#���=�����a��_���U�B�����p|���e^k.r�hg�N��*�ղ6-V�u��+y�n����x4�����KXZ�/S��w+Y!q����XR���Q�`��w��0��dn��\QX�8s�j��נ���E��R�j#P�B!p"��}ѷh����<��#�Bj y���6��Y4Hd�5;��ر ��l�ϲ ";toz�9�t7|�`�	�Rԋ�Wf�QK�G_�� �1�;\��a��07����e���� �8wc��Ƥw3yN�� �Ri{��Z�Գ�]ym���r�昉�J��G�v��Bغ�]��%[*� 9@.�4[�vŦ�H��R#�=}_:	����-�Q�=�T���^�x��)�CK�5T $�Fėʗ��u�0��k�̴�3#��XKXnQO�q�0tۘ�>D���ƹ��=l�C�P�x�=,��/^#.�_x"�
$�%ô��A�tV�YZ)C
ܾ3�$�O�/_?�=+���j�F���`t�)����׾J�u-vf�.��*�po�e���YMDu��e����dXDO��� �>%o� ��9�%�)l�~@��W�$zq���C�
��RZ�e�ƅ.ȭ|��Δ����&�F�� ��|8
,�O�~Y9g:|%��3Y��'\����\�\Uw��"�t����]����9��$�:au��.������A%J��[��r��!��Hڂ���S~���cF����`��ȥ�c�1�K�W�a
���6)i��<#�[��^���N�9�Rͻ���G��9��z/��pv�r�bh)Լ('vG��ܨ��������I	�X�k=�(��e�W�f�f�j0	O��g�̜EQr$B��69H)�l�O}?�r�X.��PU��P<;�w���G�1nq�\}��0K1�=�\z��xה=�}�Vkwt3�0��ZD�tݯs�yL�#�S���޿�)�R��!CM��9y~���[��q�h�sS�]�������R{#e�2���6v��LyRz���ɜ"yW�+/�拸Y�!�`�tVj��i�BVU�s��@̎���b��[��Y�X����jq����-�2X�RjՃݳo��ڂ,��brO��m�+-��(_|�'q������|g�9�Vd�����+~�v��<a���䱄�W?�����@�x����9wb���#c&�����+a�Ӿ������N�k��xi>o|�~EN.��Y5L�>ܦ��PLwQ�6kbY7��銍��mF����f:
�R�_���z�@�t��s@}=��G�_tKKB�"�Ei�Z��1uYď�8C�{HN��H�C{����̱]�͔<����B<x�2)a�0
V��ȟ�2���_�Ha�5a�aI��9$�^4��aჴ܋^ϲ����b��;�h<Lz�ٹ,}�.�!A3})	8��.&�n��C��q�l��O�;9�Ln�IV M�3�`��x��G�����Q�*4c��,ꙏ�G<K|��!�?8htx�ii�$&��MX���wd����We���׉�J:��3$����F7JP���g_'���sQ�N �I�@�M<��<F�+��dp��9�J�� �Dz�+`��#QN}� *a�<( ���cM��U�%6Ҕm_F����_8��gE�]��٭���<�����Q����* A�Ǩ0puj=ƺE4�v�%���4_�xR�?
��'��U0�0�`<��B��^���F�z��Ʊ�f�ܭ�R�Spd�7=�� ��4��à3��fG���4`?�A��LΤ�W��������bj��7*��O�0~�(|Bƾ�֐�I	��}
x��P���#(;��?a�%�XӍ0���y�H�q��{�C�!�S�3��-��淪��t�iKk�H�-Ƀ�-7X�l������;񣬲	�x�꼵��(���%�lhmU��J�hGD|�kFOLG�f��O��q}Cn�LΆkx����<�pw �5�ᨏ��S�)�*��=�������5d����ґ�B����=�E�Ggn�U�[�(X���%w.�]+{�;(��d�k���=m��=eQxLo>�����%��5�^k Ki��	�ǅ�D)ؐ����hF����;�qd�tc���)�����P
�º[�呮0��״qf}��u�Sc�՟�R"��4�5(���b�5A�󅸋��U>�JoL��%�VK�Y�1���!Δ��k箵��N�nHB����6�/�y� >&��Y�H���'@#���7ģ�"�s5��kf��}��Q��,� O���/��]qA����H i��Ќ�/*�Uu0���B��3ps���ՂJ�o�H����Jy�ĈJt#N\���^ۑX�>=9A�wk7.yqE$�{�ʎķ`P����V��<v�G�QsI��+�T�B�,��L�r��A$`��@�����
V�Ȥ�	#��*y��ʡf��&9?&9mD_�A2�;��Sc�����.�$�{/���qP�m�D�N�+H���?$�@\e*'�%b�#3"/�'��n)�]{b�g���[炬�UOt�������o�al�8�D��TR[aB�K�Gs���;Y�;��o�<ҥhĔ~#�<�w"������ 7��n���Bx��xY�\fI�ռ��9�5��S�/ �H6�>�,]�F����PWWϥ�M@.�V���C:��FP�8;@���(���G8���ݽ�����݆߷��邼�C��?T���/��-[�1����I��M��Q�a���a�!==�'a��L��;J���D&զv ,�|3:�9`Kzw����<�P���3Y�{���T�N,���A�n����>X����ӳs!�z�b��d���gJ �J�� x�p2����N⒔���"��z���, ��q
��k�"��,t��69�Ȥ�iO>Zb���K�ZD��X	��d��6�6^���i�Hw�y^Bq��Lx֭�q�猖6�U�)�����">�ݡ�>�˾-ǌ�^�6�����tA��;E'�E\�&�8�;�RcWR;��m9�����k��t0n|����08�'v���u���{��U�Ŝ*�Dj����7z���+�J�l3pX���n�8N�����n��)n�-���;�9a�AM����<T�f��"�c�)&ʄ@��0�����xʽO�V�׺�NG���,��m8!�u��N�S��:x�!�עQW�:,q���/8�(�]���S��OV4�H����ũ��Q�wAK�1�����Y>O��W
�"���Vϝ�{p��_�#b�O�gkva����t� ���£O��� Y�cێM�+|r��I#��u��nz-���� ����DB�,�7�~F�*�MD��|�N"����6ҮXyz.�ǡlrXt�1����sC�qi��]�T�bj��ljG�_���h�ӈ��4��/�}9�'�p�qy��]��~��/[�7a���[���1���,���e�~8���.��R�h�ڈN��V��ɼ�����V��HM!h� \x�!��r��'"�.��XP�`�W,ݮ��X60Lv��X?�*�XR�Ƴ\�U�D���g�P{�]��S���U��p�g,�u������*�����F���2U���S}�G0���aM���E��í��~z�̀�T��D�����KdռR�� �������)&>ꢄ����d�,�S=C����\���(��������s��Ȧ&OJ�o^�#�-�x�7�x����Cbr��e��V�����L�{Х��2���|L������;��~%p��.n��V�;1��f1����i0/b|��x��M����4n��Q5߾ @�ʧ�7j9gpx�	+���W��O^���t�AZ�{�(�ālRʨ��G�&����-��矸�]����\,�2k�Q��K��mm�t�s����^�k�ܓ��^�r�̸�t��������Mj2��~��w�[�X��FGi^�^y�&ØI��� ��uw֯]�Jg��x�x�� 2�}��Z���j �@+}c�F$����8��/���-��l�6@&�����XU:f`��0���m2�]�*}䗔����`�U'F׶A��0��am
���z���$ڟS;���s�5�[bo��
�'�MиH�.�_�6;��Mj���QU���֚�ϓj������W���J�GI�]�f*��?`I��,��y$�^�k��c�^H�����m�Qak��"u w��^�]l c[s5�v��a|4@��6�?I����g�������
�չ�3��.jP����f�~�]\V�r�_B�d��/$m�o����9t�룦�Z�0Y'5H)�F��*�5��[t����[z�:=x����h���	7�6��=]�)ּ����`;��+�b9>EK����q��yQ�@�~��v@Q�T�(��h��e�1��Fse�	)��!05�c�(F%�פ`�JƐ���
G��,���CI�,y��~|T�<�X4�r��6:�o��n?Q�F�ȊRmv�|����K��\DC&Ur-hC�i�����m�õ."�:�Q>�mfZ�%��/���R��H��Ũ��	�e���*�F6}*RՂ��wc �~g[���(���fuAg�Y��U{!T@��nl�5����o���ڨ��(a�IL����-�V6Gs��;�~�g�d7J.nK�<�����
������������53NՅ)H��ҏ��/�%z������(��م�˥���!}��z�.N���i��h�r��~:�ߚ�EA�xH����4�a����Ole���A�i�����>L<�t��G�S�߃]��1��  �3�bг\_ʵ��GA��B��Q"��r�p~��O	�mL	"aeNפH�!%T���}�.�|�>�Z��n W�z{Υ��A7dDdS�\Tuq��$���h;e=Q�C ����[�ra?Lj�3i�&���#]Xi���
7�D{���fw*j������ �N*JUrtO�F�w�>uW�['��8���N;H1"��Rq�N&h4$m���d�&�i�B�qJ�|�:H��k)ɼyձ������?�В���k����_�-u�N}v����`�$tD�\���^&��O�&��곑j����]ft�4�z�2,������̖(ovù
��֟�bM&���.|�JD[������90�m�:(��qP/t�S�A�hX���?��mfr��8%��j��9V�� Jq�>��R\���'k���,q��F%ا|�x���Y�����;����tK3�rɝo���q�Vz���!s��t��^ �Ԅ��]V��	JB"���w�`����$�3�IO,��.�����~��]}"WL���$����˟f��zu�'�D�ʾ�̈��䴞q63��W������qA0}½X!?�nN�N��zS�&]� ��)�^���߱����^^�I�Gm�ø�\���x�"̭��ݕ�V�l���4y����h���}<�H	#���a��U��
��nj禐F�!�U�K�ʁ���sd�sBS�x���(�'�,Npr�����y+�Ʉӝ�������%O��}
f.Yw�l�jo����l�k(��Y����:C�ɏbM���]oON:N�8�o�+3v
�K�_[Mʰ�"m��v��CN�t��2�E�:md<a�Bb��"������5(��x�+�j�
�����B����ׅ+\���:�4�<�98�t2)F��y��h��ԋ��`�<�[Y ߡ�E5ўO�dE�\���a�)�Y�}L5o$c3�
,��?���7ɝU��>)�e��ݾz�m��Ǉe-Ű%�����g�>l�|}>0�_@�Ix�S�a+@�{���$mOJɦ�$�/�!=�@�-�A�ZC��T'���,>���d���)џx1Bm^A��Ŭxui��VbV��,��.�	�|}e�v���AA̬7{8^̉�t;<����� ���%�af��"��Ԇ׾L�ŴG�5�|�,�Ly���2�-�q#_�8,�4A�`�.*._w�$3��yNz�FN8u�$Um������8b�_1u���쎭��=��s	oƤ�c.w��3��~3�ϒe���3�>�C$�����e_dq+�M�'���Y�V�B������b��PZ�7�s�uV�:� ��j���G}.�����Χ�[Y��\�/���;�,EEk?h��re�ѡ��gU�J����'�g|��%�E�kY���U�g6YVD/dɨ6Z}t�[N�������C``�A��O���h%(%�\
� ��X充{�;c0�+:r��Xn�D��M֕���:;5������an} �X�"�6,D֌(�j��h��&��0�	6ɅB1j�mk�g�4��7�������->U����O��}+����*`�of<Z ;F�G���C[_ѹ�f٤�	��;�A�����N��� �* 8����Ӛ�.�fK5t�Z���1͠4��?�Z裝u2�����ƹi�N}������k�(���:�%SO?L��/�R������~�ٳg�|=f5��[>C帬9��^Ǹ�`��u16ǒ�и��Q$4�:K@ � �����a��QG��?�s���Wc�B�dw���N7"m���8����g:UIt�K�x@4��g��"�8�ȇ۹�u�mu4��\�'�\�Cy�C�ݠݠ�*>0�R��2�	2�B���3��F�[�5�
��F�e�{n;���_��Ĳ�Pg(�
Q&I�;�/�-y tONA���(w�~�>�sȡ�\�V�-R�(��c�eG��gh���E�Һ�y��O�؀W����%.��⍚�LB9Q��pHɴᤌ�P��՜����uH}��j�d#�k���So\5���ꋾ~C�B����:6kW�YdS�4�̞NR�(�����_E�Jv����ji��}8�t��Ř�MPL��pV�~Ҳ�Ѕ³�I���< ����=;�dP	���ٳǱP�үJ)��l�~X�:���=��g��3�+�����3Uh��rx4�Y��D[Q���&�LL�>9z�s_���-]�w���'���ƅ ���� :�uT�嫷�%FOr"���Т4��fiM�E�$b[�5C�{���R�.P�~��0����I~��[���z:mD�ݨ�b�(>ݜq�+pTrX��x&��E$�f;���V�:�-��E�*k������40�ȉ�j����\�vx�''Ĺ�$	�*S�t^�6�����%R�.��ӟ�Vw���8:�1��Ĉ�I��Q�[D!� N��Hm3 �[�q��Bct��ɅRP��@�ٳBa-���y�8%}>�~��?;{�kɽ\޿���n	�k7\⫻����D��*�����FƟ�١>�k0P�M���޾�����)�ts��w�V�<҄� igq����7q��� 'ȉ���Z�j��������������U�@5�}\�p�Ӱ��Ҥ�_��֦���oĪ�E��\P��iB�����7)ȇ����-1T��P}�O��<`�2�+�M�ɚv�:�p���媥�A��E�q	�6�&��.��3X�f�[��&�#��Q���h[P�E"Dc�n��X;��/Cm7�v\�Js��ԶF"l]5�ۉ��(���'1�'T$�{22\T�����*�
�����/���@�qK0�)��I1���v��-�4��b�ۮ����~�P��dAxIF�9t�(��%R��|�t�7�޻���D�Ɋףl�J�����G��2Ѯ���miƴX����~g���߈��W���]���=�B6��p]S�� J$2�r�:Y��GG(�{��"e����,i�����Ӻ�A#�7,=w�?.�gS��l����j`T�iF�5��k-,E�9��`��%�]VQ
(���6���p�lK���#ѫC&������i��ha�ǀ0�58�hI�����I�M��p�h��f�$�2g����;�漑�!բ$O��M{��u�Aҷ:��iC�w�G���Z��sl��S��b׬�	��� �:�2���K#�1m�rD{�u�$�}Q!�c�ϭ{���SJ�"�hʯԍ��� 3_��?�7M���sTA[�9�X��"2��UW���{��@��ɴ[����l�݁����kϛX��x��*�ݑQlv�nm6yʩ5�ҙ� g������uγ���J|�c4���)]�k�*+D��5�ppJ}Ug$s�G[�k*�>����pCsEPL��x�du��y��Ji�t;f��T���MM�L���<�}�(��<[Q�Ě����d
�;���eU�c�Ӹ	~Ձ�D��p	�bԂDDu� �n�"V&��I�\�>��ΊZ��:h��;�EH�k�U�	���u�/f�~g}�P�x7�3i;��3�hn/<[�K|�u�����|��õ�ۼ����H�2K>�y{�*qae�!�"��Tpg��~��]���:m�!{_�Z�SISE�XnN���*��+��Q���)��AĪoB.��x�&�x/I�����7���q-^r)�	�$>g�*��b@Xl��r@��3qO�|F��.@:��@��'�X�F�#��ݠ���ԸS!�� L��X�J{G�ʊ�k�ݝ�B�+B(����c�Bk�]_~M}�%����I�Ӷ�T���Mꛐ'�v�6�������I����d�S��Y������q{��*�PdX�&��FζG/+Ԡ�0ft�,�%H�C���hDW�ZsWq�7�רS��w~����c���� )�;�f� ��~8��G�d%�Qp<�I9>ɍ�t,��GT7Mj������U'V��Ǜ;3�#�{=������U}O�̸�[�o��Ӓ�1u��G�{2H���M��ӭf���	�o �jo"(���.:��9�6@��ZH�b��d"�����Y���'�C���hL���M	&h��/�fO����nڦ�22@cu��y����ܡ����zپG�ESַ�m�!3�oT��d�]�����k"��ΟM
�ۖ����cS��!���qj�`���T��}���M ��:㠆˶#��d:4�R9p�ؿ;*������b���8aH�O{ɲ��2#�Dˑ1�+PDſ�d�}����y����`�k���SeL7\"�>��#�����]�?�+xV��B��m����L���̤�"p�{�h�I8`I�6��/�m��c�B�<ZP�T�FƁV�P<�q���>�c:/��N)�{��0R��7b��0���;�E�h�|�{.�TظW#�q�β��~T���?��1�τz&��zJ"�[��rUK?Җa��]3[��e���4Ʃn+�.=�)���ڌ]x��N��[E!�(�7�r���]��.���&ޤ1ـ�C�h�躭 P"̺�p�~��y�㋞Hi{��,��~-�`��dK�?윸��T*�y6=)�����������Mx#{�t���t�Wk�M�v�%�Fn��<�Y�(zmʷL)�����ݪ�mX�g?��h�x�,7���丸�%��8�P�Q��&L����-���H $5
�Y!�Њ��&A!#�?��/�R$
�"��?{�u�0�q/<���V@p�6F��0��<�f��Y�$��+n��mo)�`�Pk�8��5u����kv��3;B�~{x&	���?H��}����+F1mZ���;��ľd�Xc���i�)�LF 2V���Q}�!�.�7�8�Z [(N����Z+�l.q��Q'�)�Y��o�u
]~�^U���]Cl3��Ң �>M�/�����:tt����B�C�{	_��g�&r��F_k�7���y� 4ا�������§PƂ��[=�s�s_����=Τ-V�_���RT���Z���N4�d�Tm�މ���� I��C�*��]QbU �>f�P�	��ʅU�Ӿ�!U+��s�u���a��=}8{�Y,ֺQ5�!ʤ�0���s��-9 O�#�Tǧ��,�v�i��HC�kA�(��,��D:6��m���G�E5��mF�xˌu��.-0����g~E��l���gy�ż�/��S�C��9�}�n��t_�j�tGX��ltx�d��?��H-��L�̄�����a�S9;*$�G)(�0�=�C�˻�=�F_�+g�������g�9�hQ��ҙ޲xGܽ��J�O�#~;R{����*�H/��h}4�8����O��x��-E��Ha�$�І
=@yVJ��Nc[���8u�y��N���>S!T/���j����,X[} Ԫp��c��ҝ�m4��z�\���⬔�U@�) D��#��ϴ�S������+�i�g	������LĪ�]ç�t�_�n\�B����rYŁ�Ǭ1�=��O4e?ę��Q�ޜSY�>�f�x�I�l9|�=�E����*�ʙ(�'M�If0��
-�@>:�0��Hg8O!�8����~�0�u��w�8:)`��h*���$ᾕ�M�����
-������׈�g���:;�n�����{d�|��R�>[�R�h{?��%u�x�jw����	m
���Ϧ�-��\��+P��'wZm�d1+I���
�F�g�~!g4���(�Y���Я˒��[՞�fC��؛�.>4"/����l�R��|J7���,�x���0�#�ż1�g:�y�ì�z��j��TiU}���5��Z�aߘH}�R����@��
�&;TI�_�F����#|����ڲ��|���h���@��,���8�sD��>��ʼ�����u�̳��qJCM���: ��5z+g�WW��W�u�~�X�B>U�����:�l�jv����k'L���&�Y�[�G7�"��� �$�����DDt��X��2\�b��
� ���g3��e��d�u[�<p��h/Z_�=��#�x�w}�ޝ�.��j]!��x/ɐQ]��*�_"q��d�������NѴ�f����lx1` о6�/R��g '�	�Z�0�6�֝x��&�^��(�M�|~���=��"��d�u��VC�̓���w f$�eh �^50H�G�Wޛ
y5�T��)!�;5�~tֻ�+_�=N;Щ}��[(%�{,�5��7Wt{Li�
�����I�䛛�~|
����=��dNJp��������^�rq�A����h?�;�ij?��5���<?�a�i���9����m]���/'�����JOj�d�'��8�B�קgX����8A>��#PZ�`��NI�m�V���
���$)ԧ��Gq.��\㑑	��]�{ב��FH%�<�7k��o"�G/8upax����w�,/�k�1�m/�<��!�
F9v���ttIt��D�����{�b�{J�7��	�֮ȍK�I�[Qְ�FP�0�U���V�[|����0��_`�9\-QB��|�2h�\����D46i�d�B�g7�cM(���a��K+��~׷��
�fBk�3�q�����(`x���߮�9���pV��b>j��5[�V�ي��J���J߂��$cS/H�s��RK�vM&lw³��i��8
DJ��$��uLHhy|
_^���97�'����3N��ݨn�O�ܡ�
#�؀�6�%��6�O�q��V�G0��	����#����UP�S�J0�_ferh�Mkx��@�B�
��4/ɥ��������j3�j-�� �r�#�z�z��`]6Ў
R&�F�و����*��� hk��9� ��/��sX�l��K�T��%g��ʀup�+���1/j�fÏī��4�->_�)�"���)m!Y:�
r$\�C�at�G�Y���Lbn��!1��T1��=�(�/ڏ�ؿ�ʣ�D�Z�D���|zI��Y�����*��9�&�I2��i�&�fmk����S7�(��Oo*�p�\AI�h1�^Eƴ�Q�F2��ƀ�9�f�!���a�.��H����I��O@:�$��n�b�0�r�s�l<�x%��_jC�cC6UY�����T���k&f\o���>yC������L-�;z��ݡ-��0�=�;'��8D܈@�y�爉��ݶ��������IA�;O
��܎�2�!��}(��ǣ$�x��$��� ���0M�\���E���{��(G�+b
j�(h�g�Ե��`bFJV(Ye�q��

g�t��O�r�Prbn� ����~��#q����~��(�1w�Z�^*M.1d��9����r�`W9���>"��p\��Z�v;�η�%`d�_C%'Ӻ����U7Ģ ���I��|~�>:��/�L�s���c��k�2�p7#���]i�:��T��������.S�b��˻�$�C�7|y.k�(?�8"/3N������y�S��KZ�şʫ\�6r�a����{�3^�w	���6ᙡ�Smo����ș�<E%�D���鷷~���%.�����A�T$eޗ٘&��	���V�P�~�"f�e��8���p��M�D��fy�fS�ّ�<��W����k�}`዁HS�
O��x[��bYX ��G{��htx%�+�����=p�����U>�8�"�0>�#�V��Ot�8H:l�r���;�?RYj������bʿ=�Q��b]{N�t�e���q�'m�0B7��6H��5r����(=�`&W!
L�c��:r��D�V��Ͽ"��<�YI���- )��!�QG��@II�����u�{5�I>{�Z|r�F�|�sQO�Aw�{���7m���ţ���Xθke�8�J�S�ߜ�1Ʃ�(I�|
���#�N"([���n��+�a���n�H�`�g�W]���t�*��,g���h�n�I)[�i�N-��/	�5��{jBp�vt���bz(��r����2\��O���	� ��]��z�fU���6xzA�H."���b�5Ȇ$Fr�>�Ť�I�{騜inL�8\�Bԥ�x�q+0��d�:)�L�����v��|���qʊ�V��x%�\�4��-*=�=6��E�]��r�uv��@��k���O�`�	ɷd�?7Ĭ	��O�9���y�WwG7��5�o�H�~�v���Ӷ:�����.F�iW��Ay�����J?=p��������K��ij��E�����B�.��\ye���'kw�%� �?Y��Enp�C5���t�^�W�)X4�=k��{a�B��_?yP�W�=�^���f�;/����Im�0*zܼG�O�L�J�<I��Z𩝍�x�5�-��fMڮl��_'Hz�~�����\8q��l���<b�xN��2�8X�kTcFa���S���h2Dmƻ\V^8kKG�Msd�87�YI�be���(ݲ�Ǥ4�@4 ���s���.mW*q�3ݢF�� ��dL�v�9p��X9�q�:g@8�Z�$�P�}���Y�:��J4H�6��Y��f��3+����-������_b
�����8�$��)̣�Qu�y���zƓ.��H3�`�Dґ��RP���/��*��� B���ղ��g��n�n�dOC�k���lk%V�/�f�,���A�%�%A���s��gk=�1pj�����u'6E*�<H���d8ښD��1�*n�T��u�D�K�"�oƓ�F�D��(�^~��mN�W�%E��ȃ�(�'+��Ml�F<���U�./���ޣ+Z+��G�g1�y�d"���SA�CǨX���#�Hb�����7��<{M�;�[;W5����h�z�į�E�ά�I"�����j@�"#
��>2�r��ك�Z._u?�ע*f�:�l�!���e�rg�Q��"��"ѓ�}��R�h{k�"�l�Q���G�W� Ќѧ�l�e۠��<�'��}U����D���# !58^@�sq4 ��]G�$���{ǡ)�0���qqPb�c�癿W��x�Uk����5۪�J ���N�X�E���84~/v7�V�W�ۏ*N���)��,��v������q�������"�K?⳧	��ՠ�y��L����|�K�%3���~#�P�{�,�����)��:z�j�pm-׊~R�m�N�$��_��t�I��*o��*\>��L��e2e3�+V]����[��6&�כ'��3Y����P��I� +u�n/�������1�0v�*�k�:a�����V�'��v��{yp]r*�&/�?+@#��wI��9�	�k3�2���l>R-;K p��4�Đ�*�ICe6�e��:X�t�*��'�O����FĒ^��W�E���fP�Hݼ%^h]{-r�V�R��c�:�蕶�,R$��R�v���Qk�vHeEx����e�t���3g�ϔ;]b\#@�l�Ms�)$�;�~��*��밖�"�����wStʉ25�p�`���-��.# � �FHdN~���@�ɯ�̲>r �/7$6w^V�\r�������7�:�8^V�Z��]���͠�͈�6����.C�̖g�b�'%8�Z�B�
+��~�=4Km#��nD���t���,�R{jh�{fV�~*��C�ލ%ԡ�P�����S�Fh>�$L}o���SY�����=�����O	�x���.I|'+�4#1O�q�G�ӵP���0�m���O��WT��q6��lxU��NSH���h=Zw� #%���&	��~P��i���I��џ�)�2q�y��4��lr����R=���^3Pu���.N�6�?ē]��;Da�$��ME �Ao��rC;�S2��~��o�L�}��_G���i�D_�����s"l_�],ۆ�����T�mځ�����'���Y�##FI��b6;���ó�-�ў�if�����N��w�>1S�!4N�:S��5΢��be*���ۼ�~��TV�Bդ�9*:lj6%^��o�f�8|x�:�ǫi�ͫFvƟ_j��Ȱ���&H���]�p��
������������p(q�@��h��IFoa�|m����^m�rQ�2�����Bh�9�э��L�/M�f4��[4�m������������=`�Rr:��Җ��Nnp�
����}f�U�G�. _�Gy���q���%�C9nX}�G��Yy�+(֗�#�F�#.M�È�u�(⤃tP�{�G�~�%��-�$�`��'7|���Dv�o�#a'-���>	����h$@UnM�f�s�b6Zp *���Y;�YSg��mTjX�P�nc5���&���SE���8�B������d��̤4<������A���6V8�� ��56��(��.Õ�v��#a��J!�ٱ��`����:��+��]���;^�&��5���<����[�f��������3�Y�ǀ�R	\�9Φɚr�*Ps}'V����a��b+-�W��8�j�>�;����t�X�6�z/����"ә`��Ts0�2�Ky� K'��j^K����G�VP�H�/��RELV����w~>xH�{����o�Jg~��,��TE��I �k��$k[���
�a6�={��c��94�}�Z������S0>@ĳ-��@V�Y��ߘt�=��ޫߘ�y(���	��\��an������i��%T�B��I��e� |�q�OY6A�d�j�k�-(R�oKޯ���ɻ��u�&�#`4hC��7�yW0�����V��/�N�wǟu�6�D���0��@6N>w���	&�t����:~ �>ʿ1���*�4�y�?_4�$i-�!$�Py��s�7i7�O��<<���5����!ي�� ��~����g���o�eA�Έmr�Dv��2��O���L���N�8��Hab�n��>D�����{)}��Y�Of�q�����!vp�8��JE���+��[� 8��z�"�?�FGyR�pR�2�a#���ᓀj\f��������S���I�:�,�`�o��N�P�Տ��ӈgD�"��Δ�&�q�$@C|�+LѪ����TBF�����T)��7��`���5�wyP������>�$ՈL���(;#�K#'h���S�ȝ"oU|�e33�x������&.���mK��u���o\V���j����4f�VG7猐�����ۧL�H�5�Y+�s�4��8�2����Eե/�u�=ģט�+a��,8�
yL�^w��^�a�B�G+��g�<x�ad<l��y��%tĆ��C;�-p��y*=t��m�\�����^y��Dz4`�����:jQz��+�^��O?1wK	��W�GU,z{�9|�>{#߃9<Z4C�4�6>��R-��P�ʃ���&y����p�rώʲ�$�|sg�a�k�{�v���9�m�<�V�5�����X����t����\�ݵN����\	M�R�����m���5�!$a0z-A���zJ����HZ-b�>`5d�`TF؋���b_��x��=:#3[�;V9��ațyo#�Wj���69�3*pS�	8��	,C�G��{V�	��/�@���P�l��$i�I��<�[�m��'�]k:��m0.C��X'Ee����)�IgPf݋��B�3L�P��7�4{NؤNmd��t<�LX��,β[�Nҍx�h�ctX�l���iHť�X�{·�(���5_<�2�6���\4�g�!��SQ���*��a����[�!w�[���hy����0p12p���^-g�s�\i����}��[Ky��'QӞ�~�&w`�8D�����\�\P�hJBiU��EQ1��&K���ɘH�����Lv=�}����PD��|c@d�(�&�1���r�u,�u����#���?� _��ɂp�4��9�Z
ފXF�'n�Yc�"��M��"��r)��.+�k�*���]	���(��
|R��Ǯk��J=�U
=&@3on{�u
�/No7�&���$�QB�B����O�߼�Y'J�ژ�=n�w��,,�F�mЉ�'A��(�|��i�e�+���_�F.���b�AU����z��L{{*V��K��b��H�?Ν$��(�R���4_�9��Q�́������&�;�[�"�b�� \Qx��
-��d��e.H�iV`�7��s��6\YW7�m|�|5��aҦ�Ż�9�'\W��FoS�A$��*�i�U��8�i),,��v��{�~LҶ q���8�R&b�����}����������dȿ7N�W���Ut��=	�mK%�α�Og9hPp��Ň�D