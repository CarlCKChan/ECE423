��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�+����Rq�����������+�nS�U�F7&���S����"�M ��U���@�˴�5��.� -;P�~�oa|
)k���BЖ�@�o�v�4ߘ<��4�l��D�4Ak���-.b���mC*��D�i�M%��%�k�~&ʳ��0!����nY�qe��3��ck����o��z"��,f�ը��%$���|�;+#�0f�UhOǃ��2刑�Lc�����|��|����Q��Ol�pf��\�4Y�
A�Y�a@��qnNAz�pד��ݮiF�?��'~&{�X�v����H�	���Gʲ���dӤ�>v�� ���K�B�x��X�[#s��W�V��.��f$�n���:Qn��24"M��<48�}[�� �(�5��t�L�6����ئe3Xa�|=�X$nD�H"ď�Vl��⼞=��5��n�Q���6;#٬"I�L���P����/P=�}�㟂���C���?�ZI�r�	5��]%���ē�2FTC�Sh��Ds]鉬�@�0:�?"ܮAۙ�>���?��i+c��$�vf�:��P����LX�Z��+�'��Y�}�G��)��q��ʋ�X�]���ۅЅ�aڴG��i����(ް?	�P9���y�
�����E==6�iS��=م�gU����!��8�د�§���g��d���B�Rx%��E}��8�!-�U��@=�R ��s�/�ǥ�;,'�f��|�<�\W�21u�a���{-��������k�����@b��G�9SK{[O��Y��7�vb���yS�����	�63ǲ�Sr�,B�/�t�(��� bc";W���"-�����?�1\�ؤ'

`�x��4Q.�H����E�l���5��S���kd1��{+Hڔ�խ8�|$�������؄+����)���gn��+砯y���>3T��Xw5ӗ<,�C���   ̰�78ys
7�s�m�MO���_���t�3���d���*�۱�)!܃�9��-�J���.��qkT�*)�
0�Fx����t�g#@p��s���(��ܐ�q��U)ײ�Zƚś�!����qp� }�̚ޒ��	�v4�nMg�c=�^�u
����6$�|�Ct����ogaZ�U"�3ׄ�)�~0*1X���vq�����Ւ��-�d{��*Y��] 	Fy`;�������K��T~|�uw[�����rw5������7˕L�vs��U���yvo���x�vR����fڲ;�^�+��P��o�-����ҹ���J����Y�C.��@��O����cd&ݯp+L���
�F��Ҋ ׷���é��s�QK�<�i�B��K�T�*7"�\��<����0M'�K^��A�Pd��,��o	R5oj[Q��\_&LSrXMJ���#�aq,�$�1y�Ff)����zP����ᝏ
�ڱ���Y��ޝpB�����V4�>��b _���FPKњ�ث�(l��|څa�l�>��P��t�e��ӛ���ȩj	x E��ML�zB��E��]W_���bj�ڭ���E�Ŋ� \�z�<I 0���1�:p�\&U��� �������>�"Gb�g����Da�Нjh�l����^���ZY\V�2SJT�"�7s<b9�[��ƑQ���K�'�ጠz4	��N��Z��fUnsV��T�P�L�H�ˢ}!@�KGZ��˝��k.	��#D�$�t��Ƈ)Oŵ>��> %OK�\Z�w�B���=.�[e����-rqr���?�B�ށ����NA^;�cǎT�m��w#I|��M4�#�o1�W��3wmN�j��6���e�D�]���oz���Mm�R3��U���ȅ`Qol�z0�?7��G}��Gm��\���[�vu��q�"kY������9���]
�	���ߌW��KK�x��t������	�"�x�{�:�ѱ��
5��xҶ<��\q�f&����C����?�5��~" o�q���[�[Q�Ir$���O��������+K�e�M��6����~�!4v1�)�b����1Z����=uMg=��k:�դ�̥ �#����pb�и�W�l$h�lJ��ć5�Ώ��Ѳ�3�����Ε�W~��Bt�����ߙ���G�L������>i�*��*>���U?�����٭-��_�KÄ�ۭ�?F()������[n{mF�|Ǟ��of"O�Q�wV�V�,P<wx����_��!���4�+�p�[ۧo��/��\{&A�T��d�Z�� H�"�Pek�g�T�i���>݆���J�lrk^�bPQjeZ�'��t�W^��%��j/��Jb��u�;�]ZOUT�5�:�%'6h������иIկ�`_%��)V�8����%����X����q���[�����᠛%��
�j�p3�Ou��`ȗNU�џ�b�g:[d��l���6h�`r}�&q���]e��^���&�$7�c�qn���A��9�3GIkiS$qf�"dt�(��Ly����p���?8DOK|e8y!c�u�}RD�y�w8�fr\*:}���H�-h�Z�j�:�ސ�};��h^E����zI�Z~�va�(�y/ʚ�]p��S�5�1�Npk����e!aݰ�IĬ��w1�7n�s��[y^�}�҅~�u�em��ǺB'-U�Lv��c�La�տ���޼��u�z�_�	�� �PO�S2�/`�X�-vǖ�'eO�#�c-&�F�s�;�a!�ߘT2͜��A_|c�������}-ꀍ&V�	-����.�u	<�TL�a)hкQ�q7%G��\�B��&��h ͞ҟ��ĦfIaO�B6�*נngx�t�|ݲ��{�~	��c��c���%C�p��|B�;fk�W0���@}45����~�i蹫i�%s&i��N9q	Ѧ�*�0�I�^��_
]jXM��ɧ	�&�bApS��abi$�c1�D��:Ս�eT}����	� T��w$���EK�O���\{�ΟGb����������K���L�CX�	��C��$,'rL�I16��0ۧc�-�s���2"��V\n-~k��Y�F1�Y��sj	�ni��y�̑����v%e�J�}v�� 2��O��մ^R�ֱ�C������W)�tk��*����d%S�>?d.0x�Y�^GVk����uF�B�,�l� ��z������ĥ��{�M� �/������q)MW�|�ģ�}��/�qw /�vz����:�¦�.db��du>���
 �䜈]�s0�)`�*�H�F�`����v�cˬ���:��E`V;�D�r{�_��2��/��������c$��@�g1�������(��')����Я ��c`�~.�.�Œ.%_ٌ ~0������D�S���R�y\y��g�c2 �D����LQT z� ��������$8�8c�	��;.�J�q2�hZ=�'��%�ծ�vѷ��8�m.�1���QR� J�߽�T.���>�mMi
*kS�I�l�t�t���o�ha]q!�#�Yp4�\�_↛��hfF%�oj�����3�K�:�����05��Y�Y~��~Z�w�3DE\�r~��1�����z��H�8��|�?.�B��^W:(������o�*N�/�X���9��1tϬ��?��5̀:�"�hc�vq:�F���@���Wnq*=�lk��Iu(�|*���1x���N0	X?�)D����q����t�{��7�_2P���L๼y(�"�C���Z=H��p3ۄ���o�GC[o�QȦ&v��#H���p�s�J`̧�?�]l*����"��+I M�����^����L��j�X^�C�d"h�J��m��n^���`v����:킢��F�V��0׺�0���9�t^D�*�c�~�l!24� j��ňEK��E�)�7d�W�m�i!����+�β�cTCnU�z�%�uK���� T+-��Dz8��lW�U�R�X)��FP�-
�HH�$�c���0��ck�]�'��/Ǥ,��N�*��/�ߚ5�s3����x��Wñ[C0�%�������e��b8{&à8��/�?�T`!����DbȦј�p��l��꞉z^��S�5�R.�}�|y*�9����E��W PfQ�� ��@O��k�ܔ=\���h1+��y��?�`H�)n�k��vlrW�(����Po�G"ǰ_�mc��ŠL cӳ�u�Qi���9��/�x�c�5z)�keЊ�V��~�2��=��鯉^�Vi�����h�s[���d�f�Rث�)�2��L  #� #�医�J�(�
�YWK�$ 's�p���)�h�Q!�4�IR�oЌ�.���Y�M���l��$RBSP@�OE�-����w��	2h�w|�ӧ�^N��m��N�Wz���������y��f��;��IU=h�������Ʌ<�e֨����5����8uqP�Dz۱ ���+Y�"8��4tA��Ht"E�r�
��:��p������3.ו
 �Br��sv+
"�k=�����$�5ب��T>kj���H'/� cܰi-:pHV;�@��F~����!��s؆Ee��wd>y�D��%���#�f67Vů��ScP1�yDH��6B&�]�`O��u�N���*�ޠ'Ӏti7FBPNܕ�g�c_�16���MA��D�#4�s�+ҙNïx��|'30Q���,��[v��)
L<PL^Z�Hw���U�J���!�ަ��c��͹$*���nx�y?����8�������+��K�M~2���h�i&�nAu���i��j�4�o#�����6�ThQ�G�>\]\T �{�o�qF^B=8�Ok�o�",�H��v<�����e1��u�H�� 9��"�N#l���d����FYO_�~�u��ύ�\�D󃫝uO�N$�϶�za�=�.»J��gy	���j�|���$(x�BAvyU"q��CMtnH��&�J5��P+hp���P�W\�Pl��c/)�eݴ�7�-������||����=�GL�|gv�>C�1U��3��b�c�
o��i�FU����S��玹�/��xnْQ慥��G)��aй��F�ߗ�t�[�7q��;ݬ�� tZ|�8ns�� �9Iy���~Gi�Cazf]%p��g�H����aA��˾�&���=�h{��P�B� n��|����c���3�8\6��a��*(nPO�.����öx��7.�q�G�Y.%�DD*[o���k���I��3�4-��<�-����y㷕�� �7c ���2^�����_��-�4>d���Y��w�%�.�<fZ�M��yI�j!��m$�ܳP����ǚa����9j�T	�K"��\�D�1�V�D�,P���Հ_ލSh���w�4�����aq��K�W��Q��b��M��wƤ-n:�����#@TN�߾π�KpU��p��Z�x'��0!i�ҙ��|���S���t�͍t���5����YhZͼY������0���e���h��ϱ��t������)�5�ף?�pX�]aV��W_��Bl[���\��p�kN�5rr���-�`({�����~B�R��C�⡼y�<�c�Z�/����K̜֔6�<K�p��$X����
0�c�=�|�ŏ­��S��4>SbI���Ke�	AP����C���j��bȡ���C �6�Q�LȜ3xvqr��9G!hn�C�&
�M^��,~ ı��Z�aR<�v �_5� ���~��<?�:g�ߪ�1��5�)��+4P�X��c�$@��B�f��Z?;(�	E���˧,���d"����@Q�"�?88��B���\��΢���d��^�Ճf�f=~
k׊�*�ƣuσ-���`܍���y���C\~ �`�w��c�8�,3i�0l�B�,.�%On�ʟI��HZ?��&�Wo�8�$��3���ȫ�T��3�Q�f_a����(ﭓ�I����@a0�5Zp����AϚ�8-��ߧk��7�A{DN~��z�EM+Ϭ�{����*���b�n,�@�?	������C�p&T�b��)��v�Q���r���?�je㍻qgF�2�;�3,#�<�`�)� ?QO��V�C'}�y�#P D��JT�����P#gbF�O���J�� ��֮HI샸�rmFz��c��M�PRD���	<�����c*�Е��վKl�B���o�Gg1��3��>�eN���ũy� ���=ۗx✕����BgW��T��!�8/�<�|������k-+��!�*�;5����6�OK��I#xA*����1ϴ�"����.�XgÅ,�`�j�qU�HG�>8i3��
#0vX��>�Q3]��� HTѺ���s��������5�Fˈ�@�G2H��:�kn�Ď(--�4/��Ƽ�1v�+���e�b���@�,��u5�̑��N�����&`!�eG��t2R�40�~�W�X�V�qMz�5}�% y��C���!��bP���6> �U�k{��KP^�fϠr�Ǣ,a����sd-P�We��=�%���a,ٿ�-�W�::$#�>=�2f����O�����59t�Cz[K����R��kޭ������9Wӫ�ҎR9��m��s����7ǯhg�]�r�#�K0
_10�("+`3������J�&1Ӿ�,�V������$�=�>�_'�ޏt�P�NK7�q��6�歲-�k�_.X�(�a�Ù�	(H���*85����(�.���߸y왂��-���[i+�V`�ۯ����3u	d<#�_���a��0��d��ӊ���Pa�?24QQ%o�mG�$��w����d��H~�a"�do|Vj?Ȭ��֗%�\ u�v$B��v��\����"`�W:�l�&�[��'�~�I<�[=����Z�{������C'��j�����W���@��8�
���潩��'�^f�{i.	�2�������Z���<F�q?�;����o��}��Wģ�Oڰ��	c�i嫨��bI^?;�BE�b ���H��"�bW�h�Ă#�aȴ?�b�;G)z�%|�&�HJ�R�ޙ�'�ap�	���VS����K3��(�4����I��G���䴻�����R�ΐP3x���ep'R�Nj�8Ph���g��$)���h���逦2xP�n0g���N�,�j�3i���	���"�����w1��-� �,�b�P�c����%���߿IOEj%�%����ñ�T����Ϭ�.�����#��&+�y�<6���M�eoϕ^�7k+�U�C���p9�d �bo=�N�(�0�
�7\���J�4���4�N��j�����{�ĠX��
;��B�B�.t*�K�\��ڍDI������X2�;�ٴ�d�z�X����x7��v�Ro��2��y�]+�N��*i�]�qw�zC��t�����!˅Ĉ�j��f�f:�T<]"�>UKn3�g���l�������c���P+��vȌt �4���1��9@��O �r�5�ޚ�$����)�W����[:y2p�ް�f��]�B��\�Y4�e���?��}�f`\;(�+�C�����j �<�Y�}0|���0�zh�Q���afECE�?��|S�݄�_�.����0c����Ԥv�>�L�'X��ܭ3��c���EpRN=?f�_0w����99����%���楀nX��D�
�J��h��+^L������L&@.� ����MZ�ˀ
8}��E�6���(o�r �퐱-��1J�G�r4K�	]�9�oѭ��3W0y&xy��Ӎ����D���!D�6�E�q�Ł[t�#+�X�j/�,����'�wW�{�߻�k�i��-. ��Mck!�7`�?)����}X��@ɼ?�ՙL[pTS���Y_;G��c}��ިJ�#��eRE} �^�}݈z�gL�|����aE�M��<Yn*3�k�S�� �"�\�H�@�zj���i�9�6'�+#Td)T�~/��R�� ���
T�-��3i��T4u���4�>�چQw�����K@"�+�+��a�Y�䈘�D�*=�Rh�"^Zy+�_:���e2��T����슿<�Gs=f�n�!}���}�d����!9\��	Lxq��%����(�+a�*�@�x�c�� f;	���7=vol�o�}�Y ���ҘU�[x{W�8���n{Iv����aS�cg�Y��r{IT��zb_�%�iR�� ���+=�{b�Z�������k [�f��h_�m�ʡ�@������V�����W��E7ЯU�� #��M���A1L�	�RR��ctn�U�@5�v�@-"�G��|I�<�!�%�L�L1��W��./x7��������o��t	`n� �~:S�٣n�7`�bN�L�� ��(�n�t��x�v*?�.��S{��[���Ϲ�O�#J��Z�x/����r�X�,�T�-5���p� mg�`�SZ�!�z ��)+�T���~�7ضGM�[�Í��8)�a�Z`���ݷR��|���
�	q��%�W�T~-$��}�?@o�N�[���Z���t�)8�\�ȩU)�v��osQ�L��O�i:���^�~�ԪC����{9����$�-�5<5�Ix�l�`���k"=�������ɐ|��Wv�|�+^X��l���������DP�A�'�ˇ��� ��C��WxT�L5��~R��Z0���n�Jq �լc*is��G|��
�����m�IBS
	�R$�eoJ��| ������	g�Q�6����RuF��kg������m�5^'�-�!�T�P���4a}�εLN'�6�k��G���rr'����G�Yg�2��pp���js�����b;�c��6�F�i���t�RjE��<�79>1cPn�d]�n�߈^�d��N��6�P{zL��xx�F4=���t������[�	_���ԝ��4�c���L6��J%�|�'��V@b�M^���"��e��*?UL6�p���@A~�_�*ܤm����tHY��Cg���'���B Z��ğ�삪gP�r�HP��֤A+��=  O��L?D���]�uF�M�o�{� �aԅ�e�Z�Z9�ȶ�1\���:MJ�=8|z�_/S�A�	R߼?lg�Ή� 2ȉ�τ�T�ow�m�T�Á�O}�_�Q�� ���M����.�s����eK�wo=m���q����V�_�
��0�w����A���N�z���n���h���cp�Dq�����x�O�n\&�jaSw�ݍu�J��-z�r�z)��묊���_�$M3��l];�QP_5���$b��ӄ��V���M��Ȏ�g����T.<�7���C�oRx�óhC��^`��[�vȢ �,#���wC�Q�$k�۽#�K&�IN��MHUBC���J�􉺌�Y�ʤ����DW���LR��;��{O�'ԫc�J�����<#���.]zwZ	��ň�I�+���.�8��L�l�����+ۤ6��Xj<������֝�7Dd�E��h[���K!�<�N����<�:RuL-��5s{GY����P;7#�.�$ۮz�� )A(J��n\���*B6`
!G�F�C.j�H��Ӆ\;MZ�j��	�J�ۺ\V��ts�9�(��͖$��(> �-�����V����6�%G����yC���ݖG ���a�\V�տ1�}xo�pؼh�������$�%��~t�ƢK"��ܞP��a���~��U���C����j�2����i�؜G�>�0��p�1�ӏ¢��9Ȩ`�!J&����ܥce���H��+�Z趃>����z�`Ĵ�z�3���s�+�$ٳ�8��!=5������R�������΄���N�~�̾K��Y�������!�qn�W35{�U��Sz�ņp%I�Z'��+�P������M ��@a+��)�E��5o�M��-�:� �NL=/�J�әs������i7K�2~� ��cH���k�1�@���(�b��w���߸<�	`6�oz.fa<���=�?���N>�PuD�x��G_��oB1|�,1��7����|�`�.Q�C� wk�'��Y�g�{ru�g�MP3K��c`�U�l9nl;o��Ӣ�����%�PE���)V�S�/��yu�<��J�_�ީ� y����jE,�1� 1��"� ��*$r4"���Z�!-��ֺ�U�2�RG,���O��-Ti�#&+���ݵT��#�^l�b��O��Co����y�Q�����������%�T��5���J Ă�z���w!�A�=�qaj�O�9&*����x���Z,�=W�W�r�R�&F-8M��\Z�9� Ÿ&��3V����7۵�!�_e���ͭ�f[���F�",�#qz��Gé��>���?5�<ǈ%��u4���b�@e�G�"Ü�#yB >�	`e��n �$�S�f������3�p��Yuh]���im�Eؑ��V>*[��.^�5��Z����2dne�|8����g;�t�U9袛'-yRy�˗����j�P�v<�P���@n��JX��s7C�*�U�qu�p}
(���b�PW3�*K���{ p�NK D����P,�ug��I�]U�y%�@�2�`�ȫ
���/��_�d$n�N������^10�Q���IM.;���T�f1�W\��(�l<����4�F�A��u
���ԛoB���!��p�JR�L%2��QKOjע�/ߤ���w�z������}����y�Zb�:�Lk����>�\��a�&ݹ*���	�;�t:M.�'k���ח-����O�FMOV�Ǥ�3�d;� ��:��K�Q��T.��_�US�� '/������i�AnS�����$��E��	��pA�od����;�� ض�@���"��s��-b`�F}[#���P[6Do3�*��Ѡ�Z�MȂ�aQ���낺9Jp���w5p`�7�Ǧ�%��U��Q��A�T�#�oY៼�1t߰�W`�G�ڸ����{�O[㮸_rP��}�*0�Ai8�}@��>A>����� �a|{	�͙���Pi'���|����c��Z�3���a�{JS(>�j��I�5��-\E����*�g��y��X�^��j$\sFA*L��zqka�=m�;�ɯ%���;|e߸zv.���^N~"�jsR�-�U*B���B�fT��/ �!��䯅,Ĕ�����iJ����9����
�A8�?���ܾ���.~��_뺈L���=~�����c��S.��C^<Em�?t�jP
�;u_wJ��������j8��(��-��eę��$��yp(Է�KF��b���^��V�jc����=fE"�ŋoP���	��ǭ(��__(<��Z����n�	�dڎU�:�*�U�t��F7<�["	�Pf�B�Ao�{�|�k��m�>D��x�HF��W;��\-�=���Y��Ԩ#9����'��8V{n{+^�gd�m8�o���%� 7��^B?��@�.�c�/�l�e�7�����cz�J�;�֏���$��@*;.�R ��ojf�I��&�#\�j����Ǟ�|��L��6k�F�C�M�:�+�Ub�	����o
?�;אS��,�]I&JI�����&���
pt��;͆~�Z�+�d�e�)���9S���p��`�hӊ�A�X���>��٘�a2��=�a4���\�Q�X��o��*�D�G�ŭ�_�N��iR���u^���v��\h,�>|�p�-���<m�U~�
�J>��Dg�ec=��.
�v�t;����*$�46,�`qi����g%k��i3}��R�/Qő;��$Li��HԈ-�# �Z��:h60� �F7�����S\�e�J�ܜ������K�L	�����lg�z�T�"�U�q���؈�V"�u8E7�S��y�[8b����@����LL��
}�p׍�?2�K:I��$��P�*UO1���e�N��?N�
�Vst�;��:�
�aL��ɦ�h���p4sO�0yQG3?bx�� l���J��-hK;��+���4�*`]�.���{g,���6����_G���k�ȼ��U>65z�3�L��WÜ[�T�~{�k��Ƭ�-ж�b�79^V0J?�򣈳\X�-�������m�Ú��t��~��O-�޺�Yu�:�c�믻zX��C?�6�X��9���
=Zs�Zi.����Y�n���n(��e�`�޹�M�(�H��?~�P��)r�A)sDq���ʒj(X�H(4��/��/i�9#][��0�/�Ǖ]���>�Th�c�ط�t������S�����[�x'|�/~���
�dԛ���O����T4&X!�j+zҡ���3k
G*,�Ά�[��:�'Hx�}��h2�.��h��.��݃��	��vb���?ߛ�N
���Uo�{��`�i=��^��T�J�qg_ن����)�c<s|���z$�����n7���Ȧ>D����:p!�g}=�t���by�wA�C��{�!Rĭ}k�D���Y��?������+y}����z��f/�Ju;�o@;�����Ǧ)8|8즛�A�aټ�<sbyڵ�{�&#����%Bb���6։kY���[��m��n=Y�%s��L��񇎋��� ��,���(��J��:z|�����?���=T���s�J��0����=��p���^���oyʘ+~�e���Xr�K��O~ R��_�f�ۯօ4RV����[F���ln;��)>{y=�/�B7,ɦ��n�x��p���'�SU�uM�vY�үu��am��!��������W�͠�j&�X�R�ҍ��-���֞>o�
�S�y�sJ>����?Q��9���6�}&���:Ήh�]��*�G[�C6**�\.8�.r�,�7��V��(/�g��,��2�AS��<��Ք+�-S.p��{vP@�=k�':ae\]N�,s���C�۶R���O���V�n���=��c�0(g��R���q��G�=�	Joź,��6.<-�Ru�y�z>����aA��F�v�����
ʐ�8y�\�_��Fl����\��$�(���y2}J:ZJk5:�ʹ�c$?����=.�Gl�-�D٣��> �|O��u���7���c/��gX�"lB�;�I�y��O��Zs�������G<��5��A5�6���bp�3 N`�)�.��Ix�[� 9��nX@zQ~٩�d̆ ����<�Ͻ�_�0ǇD�O���$�kj�
/�z�|�Y�R�C�z3 O)��?�O%�p���6��~- �LbȒ��:*�K��ۮ�ECƈ����Pfs�">ک��ՠ�W�̔0��{S?�����$��'�^�D�G>�e��쪇EX����2a��(�㢕��	�ebp��D{k�[�;ݫ���G�a�ME�T�"v\�a{��Q�aޥNt�z�p�|{�"����axv/�����&5V��u+W��-Et��yf�ciي��������	z��U�X�Y�A���E&�����z��jPA ����堉��u����g[,�I���XMN�@�`��Jq]Xt�3�̣�=��迖q' 8!�S�J��\½9# ��R�{������
|�RQH�E|�Щ!ܺ�dnv���+�6��&�av�{��0�=��7]*�PqRҙ������N�������?��e������'^s�|�=��3o����@H�f��1>��*�\���ZR.v���zgt�W�Y�\�����p���(0qij�{a��ؘE�IC��[~�I(^{Ta�����Y��^�S/�ו}�nc���Q�
�6�x�c�,�b*�\V���Bd�����nB)�ϐ�l� T����Ĭ\��E���%�]!�?�\r�{���v��ӊf�rpɣ��Ԭ��Jz����*���
�bړ��3�J��R�D['J%����2�s����d�EfG��*.�E����xJ��+je+%+�<2�\]kYa�zCwY�Z\���7�Z0�q�9{�9[��#���@i�,VĐ�6�9��#�W~��;Ҿ�:[��pK��fJ�������r`���:c���U����o�<O��v�r�$���S��"����Ve��e>�{BR���U���Ū��"���ֵ�c�RB)�Gi��:n% u�}�dk?�t�@����?���<ˏ�Uo� �����xTJ_���"�<��|M�\O���&��������G����W�)�h^ﳁG��7�����&ăק0`-�O �>j<��4v�7��v]�:A�d𪧪�����㚻P1�p�Ʀ�u��>5U9ϺZ˫�$ ���F��;w&ӧ�n�D�����$�F�ۮ�+�!��w��	TGו��8c�Ґ�luەD��%[I�P�z��B�R�
tQ��҈�p��k�]���@C|��gi�����Jzzd�J�E/����:�V�F�m���vS�.u����9u�w�vS��q ��q�q5�����a��'���Qy��fU��� 8ɡ�G+��ޠ�^]���!�@i���{����*2=��>��U�0#�vS�Dv��^����o�JL���bwD�+����ϻ�t�7#YG<���\��].�Ì�tCZ	��l'����}6Z���ͤ~#$!��yޛ!��Ƥ:9�c�0�F�V���O�zd�w�w�]�+l�_Z<D� �MG���}D4H�L�,W�#'�y�f�@�|Cb���4��{��t�e����[1�*���(TJX�OD���l��{��E+քg��r�h�'��ӗ~MS�S�����6�wK�.MP�p���s���7@�㭍��A�2U�|	�c>)���S)x�tȍ#�p��3
��Z�@܎����4�Q���'�G�t�م��hv0��Z���3Y��7zi��c�O�e[�v,���G�$�0 �ɑ]ă�գ��г��Y����N��� Aʧ������s�lqhm�W�=�B�yC8@"@���=!:o�5U����꫶&�a���c|X�ULy�F�ֲ̤DD3�9Ż�����&�r͸2l�)��ĹI��Z�hk��/w��	Z5�zgwmJ���9����8����̝ Nh��6�o�g&�xȑ�b�rP�]�yE���-O8���҉UV�-@��-��~�����/��9}�r\5a�|q��0,�]3x�<�I���e�x�H���9�q�)�}sq���v�yvv`z�p]`�܎i/����HAZ!7��A�FV�{�>OO�l]B"!�뽀�d(I�q���w6g�Dy�$�ru�T�{���mI�(f��D&��ܮ�A��+�7$&��I'�h�8-�E"��Ru|S�Ó2�vM��.x̀6�L_�C�ip}�)�X�}��{�4�������D��M��E����q!N��b�燹�^�%b7���"��ظ3�9N6�H������j�H�q�ux`�Yo��&̆!m���h�x�����o7��aHP��Z�j�Z\s��ߺ�,�z.����"H�3j���Q�%T��d!|{$�A*�_^��L�]n�E�gcGs�-뱅G%�q�[С2���qx~~�~���g�_[�b�,H��=���ҥ�^x=]�����k�f����@a�0���h��Q�`In`j���~
3Sc%�("yN�%/��{�	b2!����j���e �YU���%E�X�aEf2�[)L��1�V��9x�[����{h�_�_hE$�Q�������#.&~��#��A���<�VJʹ�]�G�hˋe�t��U��O�����۫]p2�{�^���on6��t?#^;a��."�	`���7f�M훌�S%[���&���P�[����kx
A3�
��nǣy�a̹���4�pa��BEW�| �B� �gj�ƔJr��yf�*0��h�k%�Һř��G���=�e�L������{rƚ��$^¿v��֮����b����>�8M��ϱ�G�j�D!�@�� tU����H�O���.����{�#�=n�.e�@"���`z�5���u� �D��ʐ�چ�U�.x�&�Pkr��",�f#,ǉ�A��!I�v���V�ÉV��}/��`��}!�;��L*�dc����&�~�a�����.<�}Dy�f��oQC{jO��b���=��F����ۍ�A0��Gޕ�8�Wv�eXw��K@�������2�(A��L��m���ᑪI�u��#��[��?;B����#�kH��0�Z-��y<���2�x㇩d.��T}q��h�����Ѥ�)Aͫ"��b�
��%*V��
�q�t�Q�d�=�o��)1��pH�|���.�s{r찎�Y�1	0҇�4�}��:F��'�X�Q;�ի�6��S77';�S6��8k$d��ß�_���/�S�������EZ6��hgI�Xl<��s��D��߻�����XEY�5S�3ٞ��f�*YIM#\�Wp��h�}S�>�x}�ݬ@���k5\o����T�fShYs�:�I��tT&͑�r���X�%4}���D�2�fl PUM�b������F��(�n\u/�F0@O�j�"L�r����J;�Ǚ+*�YB�o�0-A�R"�1� �	��1�j5��q>,���ֺC���c�EH�sT뻟[WP���@��7�%J�Xx��*�mw�,VR���Ĥҋ�ю��1��FlP������8Tp�ZD�|qau5U�C�U��xU�T�-o�=RͬАx�H�6�"�
��B�؆Ҵ�����`���!i�����&�P��H�!�'���D��qNsK0J��+^cy)�Rֻa�$\���Y?�MX�/�w�ۑ4G�ɇ(�f�e�\��E�Z�E\��p{N��'����3ӗ�� �K��V�G��v��M؍BB�j�J�h��� B�f��k��l.��qZ���I�t���m�R���{m*�j�|Օ�yݍ�t���NI*ZñZ ��$��~�-��Z�����'Wj0Q��:T�#B�9a�t�9^a_pa���=v|p�����|����s?g���"tt��O��y����M�E��������E@M�a��[7���n���7�a[%OQ���˓�'n��woz���jڀ�V LsNW����Nj�Z's+��Mܷ�7��n^;�B��~݃񼣲�m�G"��=����_'*�C�G*�>2����U��..�'��F�pl�p67BN��<�㷴d��"2l�0��m�mv���`2��7*]�9����F�uR5x��i.����}1��q&Yae�5��Ġ�_�lš.۰��7G�g_�����`���t�^��g	Q5�D;wi��h��m���>ٻ�e���..u;w��x��X��޴$�Q12ZF=6�y�����p-�����?4���V��F�DHR_��h�oN@������9VAy1�mo�_��9�Y�Q��6�xt�4��H�j�g�3׺��S477|��>U�V�3s��T����F�B7�:p����=�<���A����� �o9���:+�~hzP��*?����ލ��ӯ_f�AH�|��jh�a$U�iu�x4*P*�U��r/��+�|���'�Mx�֖��^�L�@�ƺj���Ʌ|�j��w�|c)��1/Y���D���x�e��q \s���L�
����I��(�%\���S��7��W�1*��^�^D��[�(��}�
A݊����7�8� �ddO��4L����#hu��9����;L�4�ze�,��.�?d�O(�D����c�5�Q��y�k컢�=!x��	0D�<� dC��j* �k�k.���N��'�#��\�R����=!�h���§���FF�I�����H��u���;��w �F�dg� i�,Y���u�]��Wr�`���@.z�W��b!�-/�=����?$�LI$oMd|�A���ZTG�̢��=hr����	{ ��d�kѐ���:׷�ԕ�,)�J%�x'7�Y� �^p'�^�Zp�?c<B��4�^T5#���>�Ү����s�߲$ta�B�������p��Z�=ԓ)�w�1�z/�	:�a&���9�H�l(D�(��Fϖ�^d���|X�@��FY �<���W{���� F���vI}�o{!��à+�k�A#Q�qT�̓�g� ����/�J�y�N�fj����F���^��2G�~Ե�m�b+إ�a���
�J������V�ֿ!������P�3:���vH�ؿrB�&]�6\���Hs,�d��\)oS�� �w^G}Hm��q��%S]�Ps�#1#e�:\=
�`�4;T{X�G*d���u������~;�.vm]��?���-��pL_(�$KV��{9�;J	�8����\��@2�{�sٵ�����i<�x��zA�v� X�1iT�v�3�_�z0Q�NqL�4�6*�2��(�J��X:K.v?v�Ѹ�sNg�S���FnC���}��J ��y,A*�ƺ�<g�Z|d��E��o��"���wl�7?�S�ͭ)D@��<�[�{�ִ��[��|ST�ֵh��=��FrE�;�p�����U�4d0.rm���x�u��3�S6a���Q������k���Pf�K��v��	2;�H
]+%yn�c��W��	�_�I:#���Kiܚަ�MA*��3u�m<f+X7< 05<T�������e���/?�rBy�T�|(�������Ϧ�H�����(�tիE�sd�F7�����n7Q^R�f-��K�,���'�J�l��+����S��(y���f�VĔ�$�M^�6���S�a�Ѹ�*Ez�4V-�:��MڛR���Y�'.59J�����"�ȩKǭV;�*ȑ՛T�3�=�U;^I9Cx�h�QB&	*3.����'��#�+�SbGX(��<m�'�Q��70s0 ��y`�櫬Iu�u�E�q���m(�ͻ�M��5��j����V�L�V�-�c��y�9�@��fē���CK�sgv����8�H��^�n�^����%�O�|7�?g�(8��EsL��8p#�ɲ^Ե�6�(��$�=4/l�Vb�b;T�����ppF��IOI�$>t�׸������<|<��������!�)�_�+���[]�鋄� "��
�.FD��v�M��/,�E��@N�p�7ʅ��#8�C�֚��:3���$�d�`vb���}���Yr�]W�\81�i��t"���櫊���@��(+}�� �j��c���7�z�J���Yj�uC��sj@�?��E:YG�&���@�BSXC�YH�d �j�|�S�lZ�9>@�po����A�z򜧇�f͹k�4�&[��yg#;C4�v�6�+�5Xk���u0%���?�f�ؙ򉌟��B[S��)��Vp�3�����܋���d?�����g��m�Dt;������lMa��X�P��R�)F��=��DvȄ�NgsU[ .���(�~0:��{C�%�2��f9jI��<���ԪX�@�УV�����m�ᜌ��4���]�A���,��/�ڥ�c�):^2͗���y@u���Mg�W<�K��C�o�~K�7F2�!���q� j�lF
^�-����zU��S��"EF�a-�N-��bI2�����)s�_AUSp�dQ�c���@��a�g&jn�Ǻ^x`��X��C��A�^�}D���n���j���N^2�j`�^���|��m^���G�DSeGI/=�~�0\;�*�����LOa�P�=��¾���)}&FNnʥ�3KKT�)	<�/� ^�P�UZ��%  hsώ�V��o���SyC�c��S��)�yWn��N _H�'�W�J0��XU�)���l���.��O�
�& �ȕ3�Ft�u3؉}��_��
� ��~E�:!�-8Z����k� �K���X���%�˘�7�|�Z� �TA��Å�"�s��d��=߂��-{}=4��l��14xg���щj7?4��^��]�Sp<a�KF i��<�'3���ݮ���r����(��Y��W��et;�^��O2���T���O���v�Aa,*GG�K^��Z^�XE��%�^=�f4��{-P��X�I�HB��`Th9�d�ω+����Q�Z �mm����E�w�m��fh��J�:���S;���D�:���ô�����$���G����R��:a&)T���QO�n���k���^<B?��?�V�ǩ!$=�I#"����q�蝹��� �� �E1����Z�������J�p����ڮ�������8dj��b����>����M�����(�?P�gM����T:�ҏ�;�;�&ƙ�[nM�CV��V<�R�'ā�~�q������dZN�J�|A.
��;���� ^�H��������;!�휽��K�>��z���/���E�~�Τq�Z�CG��}���T�/�l9���sƪ��=X���%%	:������or��RqZ~?;*XUV��w���)�"	��@�Q����3�Vkw�c ��%U��m�V�/X?$XO�ƴҟ��b��/�a�k)�M��ۊ0`�L]�y��F���ow �#[X��#8��P��QAԦ�;&i؉[xpD�>��y%Ҵș��L�c�+��h��}�V�9	�ԍ&4�IE\N�<|UFԳ��������x%�T<��)���D8�+�G�1���R"�;���K�p���C����C��}Z�v\����VV�
A��N�f�W�S��!L��".'�(x��2�hy�5�0 �x�0��o�VOCL��l7��*n��sف��C���� ,��5W�K0�2���6��J�Ʉ���)�Wo9k�Wa	�eqS��lT! Y��s��C�f�Qz��K�#'N��p��0�l��y�}̅6�j�r>o7���v0c�$���s�0�
�}�����<�\'̵-U��/���őOc�/��.�sE�=p�
wL^-�U68����)�F>�?vNE����=���^�	�n��\�}B����M㛙@��~��,�h+�~�"z0{��4 @R�E��Ztɍ$Ce.��ͩ�T�c�J��@�#�@���Kn�a;�N�߄�/�K��cs��n-{���1I<_��������Z7�3���&L�bh��?{��wc#{ۭ������xl`16�*�>�#��|���;,�l7qFO��8�z��%G����H��ٮV�U��"�7��1L�*s�q�ӎ�O؀���}�ڬUsk."���li%�{^3��&������ԙ�U�d��@�"Aa9oT��>�)����KF.�?��/��tYN�k����kf�r�L��ޢ�^�5w��_�U��q�إ����N�3u��0���C����?$HU�(��$
��1�n�V$]���I�W�������cG�G��u�`��n�X�F�<J.{ʃw��n,	?d5�q�#Q,������Q����Ρ����" Rp'T��v!1\����(��\~�418T#Jt����y�*��mi�[7Jfr�:��[��wp���ϔ� �PV~��BxM��HK0A@�����5��W��i�X#�CPH�G�nZ�Ҽ�1��&���@7�;�NK��Ye��/�܍���`S���W��%���b�4S�2�\m	X��^���v0^d���rlp_=3/���)��*�@ ��HV�g|��-�� �9jd_�B�=N�LI4� ���J��M5��ʍ���Z�ꁏ��4n���lO��_�={�Ł��(��But����2@8�3;⧲�i;\b2?CC>z���Y�!�_'��u���9nP���Er�`�a�������zי#�eJ�p��7���\8��so`��	�9�Kp�Ό,D{ $�5�Ӫ^�7�T�߂�e9��n�X	eSZ�+3\P��~[��A=�͠gw�����'�J���%��8�Qז��Pޢ���t�jC�]��as8 /�f����������\-�� ��F�J�{�p��o���}4.0@'�H����g%Z32�}����ԯ���,�MUs�̶<��̖&|`���6|��]�Kz��ƊLX�htU�0$:�����)��Hp�B0oҮ��Aiq�9^'�i��4 �A��lE6��ۊ��o��<� D���2�A��
�G�7�]������t{�(Yl��\L�C�b+�i�2�wI�\���X�R<T:��[�_V�"� �-�$$l�����+��	4�*V $Rl��%�j�>�;(ܰ�l�/#
��{>,=9.��~�46�kl]�����:���d�L-v������r ��nD�X��ɓr��4�?����(�6W�9(\c,��rГ�i�ы�� �8Ԟ����O�_����6z�/�+�Z�
�p�UW�kN�H=�u�V�m-�����A��@;,��'�{*��V�֫|��j�C�%����f�d�z���g��6�X����ڱ���/�.g1��.�(oF�m-1����{�kfa��I[Y�G���L�@��o%��	%+j���|����e���~΄ľ�{E
W��'a���n�\2�<�����ן��Lsxig�%FP&h��A\��s�5��������iz �b	ʻ;Inv��`i�O�����H��vH��<�頏����q�U	Y��t��t}6�ޚ��<�q"#�D��G�8�Ҟŀ��tN~����suf�1����4�K,�&'�m��wy�U"�%G[u����pu�j_DܡwOni�w��Cu؉%�"))����U�Y���A�Bɦ���0 �q��]Yx��<��`�ѷ6�;K��*�J-~G>�:x9J�Ƃ	"��J���ڏ��M�S�Ȕ��"i���C�)�.�s���w�h����<���V��8�S���R�������=�t�� b�ģ*��h_D�0����Eo���+��*�*��9�'���4���N��7'U�F�)BV�&1�LYh1bE���\PHR�~uz�@��zqq��{2���xm��6R�
űvc�H�˧Ӎn��U�9c&������3�:٩��|S���7[��aۀ�Z:��:y$O���:�v���p��Bʠ8��Q�1�^�q����v��#�׷L?o��w$ZKrm���8�B74�����Nq͓ 9����
HxKz\\��P��Qî�]ˍ^����F�{/:�1��_=	�36��g��zsh]���.�L>M:��C˺Y����b��og��Bzپ
�m]�م���K��$�V Ǒk|��~·
���Sp���o�j�BX�h�iU*`���w��VR���m��ZOV��6������:mܭ�GZM�f�{�?��>Fy^9T���:w8����ޗ~��`wYL�Hݲ�n_;+m!t���ty��'=X��/���Y��\�?�Eˆ #�q�s7Kh���.�265|𐃼��m{��p�Qu�(�2��)m���\PX_*]&�F(�&��W#��Nm�t
��ۡE�Ґ��<sx�;��yh0��L�UE���f�����ݒ �R+7��#����hOc�弎8�O��}��.o����Kj�$�������n9��[UsA��[3v�K_����(��eM[��yT�6*
�E�&,@�G�5���O���b�#e#MH{P͖�m�=y���1�A�N��P�G��job3�MT��-����t[������~��\���H�nz�sXOJY�?#�W�ID*NE��=k`{���ʌڳ�� ��ۗEʮ�q�*_�pƇ�)�tj��	�s����o*.�%2���ʋ�3��/X���i�)����$�'y�1�Wx0�̡�vYI����}_G���&�ȵX��^��q���\^�*��4�j]e���#z�
�Ї3!��h�Z�z��C�"�	Q�\A��̋�[71s�0�Xl�CyWO�������h� fcF�����Y_tj��=68攞�Rq�B�^�s"q�f��_���~SU��d��mū�(�n4�;*C�R�'x[���'�p)�V��C*{�� àW�(��p'Nέ�G}!��΁�89�o�$�'��Gl����噧	�-4�U��� %b�V�X��i7�\�e�Q�K��*�S��{D����O�ȯ���Eq
����D�I���I���Pe��v�0����=�A�KD��M�x����R飯�7 �a��Z����*�^����4..>\3g�T�`�`�V]`���RA�x�g�Sý$�>f���T;vL#��-�'�]u��+�j���5��&G����Q�5F�ܜ}�o�]����C�M���r�9HC������F	���k'Y<�S�%�$�Į�A�����ܳ�>��,Tw�� |�壊���8���JbT?�aү�R����pZ`���}kiR_���й�vr-S~�y5X	q;�ek�i��'�
���RFޟ���m�9�O�b��CK���^��!63�5��=���e��k�dU3�5�aq6���WfTl�bt����OZgY�*<I;�_�NJ>�ye��`�khxuZ51S!��X�B��m�ՅM���<qe�^�*�ɠ~k��g��iz9���mM��m<i0�st�F$�"�w����q�S�֦�=e~��2����f�QYZ����{ⳉvg�����'�X�cH}����G:)%�c�_yt˥bO?X$���1�q��G����h�4e�L<���'�5W�=����곆/�1G�}T/��T]���x�f��MZ��Çt0�A����D���MLi�Z�d��]�b*i��n�R4��������3����L?IF2��D���\�Y	yY�����sjT�!�����*\��yӷs24�^�ܨ�T{	1k��������x�M0@��B�x(_���S���Ԏ���o������P��TD�S+����q1��-.�2�a]tH��Tz8 ��Qy�u��Z��<s��[⑍7*��l�|O��l��:@n�nC�Qs��;O"S��0v�N~�B&n��b�Á�#@zH����w�@��-A�|�'k94�z�V�\^Z]E�B���N�,˾q�"���5N�=�%�vQ
`���!V`�o�A��W����$�Hu�����L7�Y�D#�r�\?#�(K#�ޮ�#�D�+�H<�OE�E���8����;
��<��s�>�<#���@�Xd��\ծ�Z���q����(�b�w�j|�k��̹>_�j�of�7��P�0��E�[DJ��������U�ѲO{�.�n(S��?�L�#����	=��f~Nc�h�<��Rc�Z7%�(%����k�kE���;�~`��82�Ȋ%۝���:���@��o�F�_�9�K�:K~'��ω_>��}���u�˵�[ӒEڛ��ث�*�&� ¾/k���&,�a�]6P��y���o vk��I�޾�/y���yʑ�6�S��p��%`��rn�w�[�ݐ�f�j���߃�I���?2h@�gg��fX�IAח�DgB��ԛ��������k��zPƬ=cx��4,�\Ԕ#�KM,��c���c��[�������V����/eb�׳�Q5}e?�ݧ�5K���dᄽ<����>����.��L
����U�R�&Η�g'R�r6@�>!�t�G9�M^4ą N�h��عAF@.�`c��F�P��X���
y����]	&�6�2Y�-�!��7mH��?�0��3z<�w��`�H�,	q�7v�]����ڥ��J��/=�a����F
�p��>��9�{���qv�xp6Ȭ�#é��]L�p,��&A�ܸ̩yq-F����ɫ�U�Braն�D&�?�7��DP�v���S�վ�)��6�"�BN+@({t�-^���8h��x�DWr�{�Y�����+G�F6�n��+_8��zKeJC��&سxqPU�G�>�����Qa�Xֶ�s�G�"��ӻ�E͞��Y��M��!�w��Z)���L(V"g�n#�b@���BԿ�l[�)N����m�"�5�;�����u?+��x�(yX���N	��QUM�I�ҍ>��u��o�tg� ��x�e����D���͢A[��6(3�*B�
s�ش�?��Az�����ʑ<���i^wU:%�0��R驟��KU�{����Wj��^I�C\Ɇ�����.��G�|/ю�S�e���=��̛�Z������j�X�7|5�s������H�� e��])�g]Me�8y-�r"����h�O��A�m�R���0��Q���i�/4|��������61������bS�>�]S��s;�_�i�ӭ��� 1)������/_^���%p��lMV$��DP<A��P�bTƼN��y������f��"J%-�ԏ=m�Gۮ�^�� ��k�r�����g����*��@���*B�v;*C����Jo:�<����V�J�莂�44n#���Ps����Nw&��$FG���09�+�|�h$�zjyޓj)I��-^�Z�I!��QSy���������X���ax�8���j^���c`������hkSk�q�H�g��*K�#�zkܓk��|a7�
V�*$���<�nB��V7��.�Y�'��+�N��W}wD�y�|C�-]4�����J@co�u�A��M�P8ҝJ���$��8�����ƙX�d9��%@��/s�4 +��q[��	w��{?�WHs� �"3#rtiϚ�O���=�=U=!e���mgcA��⿠b���bA�D��d��b�^�j����f��K�g���nc�m6J�ϧ�B�k_�Q?��u��(Pқ�.>
��r�Ix�d��?Ц�X�B=qC˳?̙���
q�"~c?�6�[�5V��RjΫ��9�Jm�>g$ ��W�ƍ�?����|"��q��ʑEs6�L���1!ok����`F��.G�cOD��u�����/%������w�Ƙ�r �H&�u�U����%�m[+�ƴ��夡��]O��D<h�I,y/{ؤ�Є�XT,��\r�;�V[U�r0ٙ����rŭ����m�.3}�~�;�B��)<��f�Q�ZR4����珁qBμ�Ű�Y��?���z�)ƺ�{q��V�Ϙ���$�ޱ���	��������ݟ�T�o~��� ��=�^5�. ��DW\�(:�m�D3�îZ������lyQ*���H1�ã�&�A[m�8,R^�����!��a�o^���4��N�^c���ζ�����O��� x�h��֤�H*�����rѯ��s�X%� U2��c_N#���s�zsKK�;(�'\V�����J�(�cѥ������R���6����z��z�wே��I��C�ץ?=~a�F�~�7�&�/v�y�������X�)({zxZfֱ���U �{Ϭʉ�J�i�n���}�+�9����B�f��ꬊD�v�&��7D/�GMl�ė�=[���l�fltW��|K��M_qҳ���8�Ŀ����Q|.�|���J����o�Nax��œ0m���-����`A�_9ކ?��n�"r&,��C�����]���\��$�ih̶AJ��7���ܖ���D�Cr�e�̃�ް�O����2I�j���঄_|���JG�W$������
�� ��`�+�7E�,{&Ν�!��_Z_̍�����E�?(>�.zJ�b�t�5v#�mX+��Wqu�
�CtI����{&UL�>0t��ظc�nE;��C�6x�ʹ�K�Vc"���G�U���������M�n=����a�p�x��D�5�)���}�,��a˂���n_�PJ���)_�"E-G�z52{9�W��枾$/�������8oX��9�T�t��iSp��~��͔P��83m5�~�ޝIJ���Ò"�6]1;8_���#�t���~�*�j����u����U$!$����ܦZ��
�F
<8�
�
:�9O5���i�s-�V��sݘ�هC�fѢ
}N ��SܫejP�Q{xϫ����N�Ʌ�Ĩu���%���8��Q���\H�F,Z��kt�������v\�M6�{�L��XԎ��s��B��_6�w��d�����ﭭ�-�����X�C������Ҫ��[�wA�va��j�������y �lfK�F����O3@ˢ��������B˙-��w����Śa�=HKMT��D%*�����U�C�Kҹ�D��]d�T.��ݝ����2��	˳%�1�b��C�t��6�80UY<��*?9X��9�+\��� ���T�9�|>?y�j���y��H��S'[�G�`fZ��"JGI1�,r�q^�3"���1�Q����ڬ�=�
�+!�*�z����K�P7(=ۑ��^�2Sc���KJVŋ.�x@��`q �Yh�Mit�	�{�zL�����J�:���.ғ�&k�����Tς�P�²fm0߮ל�����Q�uVS�S|.��Roՠ�Dj�C�����$�~n�'4{�
�,�3ZބM�J7�/}���>����Ð{h+�)�d���^���_7Ú�1dA�V�/Q47TA���R�`��t"�Q���}����=R��J�����1V�)�
~X|�/��G�p.k�pH5��x&|C�W��g�O�mM)�׮��?�q�NQ�uv�,Z��n�e���ȉ���<�'�S��
q&d�d*������4�{�~�v��e��i�x�%m��2H%�?,[�]w�{�9lz���ƛ�+�yo���_E�Qg�e�d*t���l��[��c�lY��8(������ݑ�����B'<�?��<��x��Ҝ(6���@�r�1���X�,�%ݙ�H����S��&��G��	��0]X䁛���	2��I�
�y����1�bϙ�̶%�w萌�tf�v���'���w�Q�Of'v�������U��]M�@i���QOA�¿�d%M�V�/�F�V�
���VvbV�L��dv�e�z�D���o"���0[��9�c���� h4�Y-*��������A�Q+d'�J���\��I�SK�>�`ae$�w�i���:2@IGe�(Ah��g�O�����Z�5��AXӗ+��[3G+ȩ�g���W�{M9��CYL�t �E��~O�9�H������+��7E����F��&��ۀ_Es�;	�Hb����Y�_ٝ�e��~l*I�:�߯.9f�ւE�̠��|��^=С�0K�H�_�sXjW�$/����eVcx��(�1=��@GxeQ�T�DG6�~J�ٿi������Kc���EK�K�!I�qX�?����C��v�$�^��I,
�6x��Q��8����/< �I�ԫ!����4���ۿ�����Iy���J�<���e��l�o/�*Z��E ��OoU�6���7v>^/�Dtez�/0�'u�ڧ���琛�;#�v!�QDw��K�:3����5$��/)L�k�C?ם�F���jG�LsF�?/�A�#�lG�Y���"�<�>+�d�d���ڴdg/��pԨ#8�[L�$��j"M;�)���S!����f��AJ��@�lk&��O��UU�;��2��a��s�Zn�t����pU5Z�ރ��mPL�8)��z��0t��JF�����(���m:J�
{	�Du�+%�0��ZH93h���Е�F{�1#?�r7��Yk�H,bݟ]�a�i;7̪����뛙�u�'@f_���
a?,jB���cd��m}�EN��0p<eCM�k��^d�l�/�-���փ ?�������`L��٘}Ǵ�pe����';l�ݻ<�.��i����*�$�ڏ,xR�k$�����0 c���	Ŗ^g�rVh��v@�*��OA��S|�b��Q��J{��}Y�R��)�V��.
��z\"����+��J	��CE��w?x���,a*+�[eш�ݦ}��}(���T�dzS�mv���������i�2']�"�p�kU����D��w�$q��싒ZX(��N˕��4���+�)Q�X�m�D�8)�E^�-��)/�`���� ��t�Y�<p�22�^%K�J���0a�"�`�ͷk*�(^6\
;̞q�Q̨��n�QB���-B8�k��}�D�)|+~pD����xB��-�Pk	~3.\%r\I��m5aW�����6��j�r���it�v*�~}�ήNd��y���K�M�ɮF�6�?�2L�T�y6��S��S�xn�U\U�9�U3ID_�ܨ?|^V�`��YO�c1���I8�>��\�v$@B�RH����د�v�1:]c�&A�1ys����CJ~
�&z����d&�Ü�FK����u��b>�I�]�X��Q����ؠ�T,�>Z�<�[���P.��V�X64��$f��؉�j�1��Q���hP�6 q�1Z��y"��ERF�taW X�W�NX{�5������޸��/��ȷ���Yp�#����L��i�Nw��6@�΁8d狤NnF]�5�����$�������pX`�Ω�����@��΁}�ި��'@o�J	�Ă�`W�QB��$ah�\u�BRU�I�B��փx��g�/��a��rSv�2n���S���K��tȼ��;n�ܬt�J?d������+?ѫ�7��'�?���[��;rr���t�],	t�w��M�b�GN&�H{���f<�:>�Iݙ�oZ�N-�(�k4̪C�)�;�t��I��d���e{�ɪ�ϕ\큍�凑���q:�v��h3��v�^="%cO��w$
��qs��/����e}G��E�[�E/�K�( iF<�_�:�����~�j���Pe���bJ����I9�n��5c�Sɨ鼆��r�!!b�B6@�P�T�M�{�p�Nc����ky�lֽ�����Z,� �Y�l����>k]����\�|�X�[��C�{��:����z/��h�4|cLF���»(`�M^��	{>!3�R����ܨM��� ���Z�&A���R�0[��6Zq'�����'�HW5�Nh�*���4�Ӝ���8�T:�Z��/�ٞ`�Ɠ�ߑݖ֋��5��r��Z��\amM��+���X�q_&��-ʠ9�G� >�S�����n�I��3ޝ0�eJ&ӻxSP,�������){��4)�L���lʶ���H5Ɛ�>�{��M:�R���-��X�K�ԯ̲h�X���´���X@����wV]���]�9;�L.t��y�5Au����r�cǐ^����zEs�Q���1)�B�`�B��ө����с�v�$��Ba��AoP{�{.����tt�")�ƌ*p��n[r���ab� �y�]'�_u��,'?�~q�������t�n8R�T8��]��qI�Â0;��&��^��ZjG�����8N����A���N���w�2��3=����˞^���Y�����؄�0���e�T��^�{��O.(����q��:{��a7k�zs�Ӊ��"�w��tI���L�*�]�ԃn1����D��*x��b����O�]�h�Mv�i�Ԡ�"���[�)')/y�QY��G�ݹ�u X*��\ɀ����q:
+����t(�hoV�@�p�I���sm�l�,�m�B�8��I�+Z�O&K�1��W�Vx�)'�1�0J��k�%�t*��UKc��݅@B=�'}>��^9#.Ze?JN	Ȃ�/,-��8&�2�C���ha8�j|��
�r�P[ukh�$��`_��M|&!�=�ۭ�0�aҍj��l&��0�J/ ��U�������N�XAv9����Q6�,��<COq��a��U�_B񔳣;�4��S���T%]��x�_!/��m%D�w��4�#���C��M���ާ�ӣ�\g(u�ޞ�����?���b��c�fG����C���is	���Lz�\�>�^�lR�u�/�a�)oq¬�~�8X��S1^7��t��z�����"�Z!��kp���b�u��=sƖ�YJ���5r�m5w��4���Ʈ�Q��?Va��s��n������x���">^�������$|�ԨSg�V(��b}�SM�fU&���0+��%�N#f�Em�
����Yɨ�kX�`��i���8�b	�d"�|Q�::�g]!D�x*��Ya<ܪ��0ʢle�\��W�B�v�csl������c��+/M?V�bԑO�<����M^�-2�����w�"��%Yw({��O�U_WX=���S�l�m�\������/s-���,X�4@��	gj�j�}�d�gܔ�Û	֬��L;���D�͠�!� �(� G����������iF������D7cJ��ۡ"�O�ܔ��9�O4��yEG2��wE*H�R=:j:Q�ٰ<����ho!gObV8�ֲ�yh�r:v�v��
H D��~��2��%H�����u��Բ!;����W!#�NWAYp\9��E��E���5�F&�]@0֝�����ҩ�g/��^]��*��s`�����7j�]�/�5?%�,�����g�]��J�l�wNRe��d��֭��BƝ�n��W�)�ޤ�7���4��1a��=��7Vv�٦h��+V���iB�ZcF,��l:��wG!}�����Z�^�m~�������o������k=���S<Ԯ�ʻm6}_�L�.6^=G�Ϻ fO�{$r���O��z#kV���d����dn�/7�'��0���aeO��U��C{~�y1#&��j������N\��H�6N�O�F�<u֋�%&)R)�#������G-�fA���xS��L��0h��>/c��S���cߒB<z9���ꗜ��>��jܒ�;,��r/e�6��}""V�Õ��C� ,Jz�M�s���I���fWщ�2Z�P�J��v�	���K��Z�>5�pF56%7�3��]�/{>�L���,`<�y�RF���C��4эڷs���1�;O�A�jG/Z�V�Ŋ�Hh�.p����wmf�23o:i��͢���m��.Z���D��l�3�ӡ�����wcێ�G	s��!\�+� nC�P��a^O�"�� �/��X�9�H��=LS��T�����{�U��F���!�I�*��6}r?�}@[|A��Կ��p{�K#��0x<�n3��a�����[��p�5��j����F?���E}�S[,O�b�w��1���Ṻ��4�GF �����L�i�[��jΰ�O�y'bа`!T~;�QϿ�aմʟ-=��K$��aeo�
��l�K�Q5M9X���K��P8}@uq �H�����s�/n�G-`��4���z�Ŏ&tx�)��
�_�l}l��a���a"�h*Y�}FXe�̶ք��I+�KIO�;<�+uH����'X�g��a阂�&�ǳ�������w�V0��87/��"�8�GW똓�9�J)�s7�\��������!�㫩�&�eX]�BY->��ٮ��*i�Cc�;�1}��Ϛ���}��vh�"+q��_	�m�~��@��4<�s���#��D���̀|�5�ǁf�Ht�y n}f������y����ԋUM���=▁i�7�-n
�5�B�Ȓ�0/��ؖ�&�)o���r�3%~86�nngQ>u�zڶV�4R����wNj�Ûz|��n=g��j����=���V�gމ���Q�.F�k� JZ���)���Eࢢ�Dc����L,��_B���U�~���A�b��mݘ��Z:����U����>-��)}�������ʽi�ʌA���H,�$8�HrH��>cpQ@4�Y����Er�8ʾ��UAz0nQ�{b�9*{��[�N��v�Q١N�d;@H�9��i�ņ7S�����(�Ύ�C�L���*��9q&<� �� ���0�F�5�q�%~��Uox��j�*α�SY^�����Y���򯲩*payoY� ���V6�����,)y�/�R�fZ�y��e�f����7�6���lK4Q�����k,R%,*���{|ч � �$���*r�i� 0�t�_�Ct���0�Te��Vd����?m:���$QS�cX� E�\��A��ko��n�4�c���tԫ�8|���";*����b�\(w�݁>kW�<��d��z�T/����R���o ��C�@qí5��oK� ��U����G�]|}jf�{oC�80����{���L��_�P�~�J=���4U�f?(Ʀa�/��:
s��c��k��ۅ2��E#ȥ��`���<KfA�U�y=QH9q��uъ�i#vXۡ��&��]@��Uװ-�5��Ym#ܗ��G>�Q���Q��%[{oIX�CǎT���vOdK��bڠ_�x�����.sk�uU�ܕ�"F��݄��#v.�D������$�d�Lj�X��oFZl�6�3�����>�T����u�ZY��?I����Uo=L*��ŵ͍^�FGNz-T&��㢍l��~F	�ʬ:���S+ê��.���H��EڒA�\5���Ϥ[��f�����6�oi8�x�/��,�$�j�]q�p��[��t���紑q�o�kC�b!���@��7���ч|.�:N�r
t��{���8��H��rglc��,�9�wO����S�����kR��8բݘ��k��G�xWU4���2>��=p�_WQ��<�`�wq�x�B:���p�2g�ȣ*P7�M5@�ۖM6.���2�S�����9|�����y~w����We��,�7�t�;�c�%3�
�Z�u>BW����k'��1��4g��M��8�j ��b*�h˾Z%tuR�UY�E��ᗡ�j^�|��'�ZS\ld!y���Y�nK�5��'O#��{������=��F�=i�M���"��R^:���e�.�!�/>(�F�m�!��4���ІL��Y�.3J8z���j�a�\�������ب؂`�aCM�������M�J�e��(��3-�$�� �?��)��J�4X�q�gx���S��lM��F�m���1�c� ߳�Ng��� �d���Q�m#.|8y~ ��tY<��WbTQ��7�Pv~��F�g2���G�|4x��K>���l�>�O\��!��9�p���ٰu��M��I/����b�r�v�[wpY�'يqX�=�8D�_j����T��v����E�5�ެ�J	�B9�t�x�G�'�fT.@� Yk������p}7��ڥ8�+�]z�{�ꕱ5�"�f�og�aJ��R�6��d���}Xl_��Zo�KX��b�7�$`	�}Uʜ t��f;T��.=>W6ѯN��rbvם�3N̋"A����g!��;��?"lE?�KA��b.���D<��s�	.���� s%cD[�Q�W�E��Ӝ���p��v��-���y�7o؁�����̕x��p	���!9#���y��#`/9�����T��<]��r��'�ІU�ʯ��3�2hB��@-NFD-�N�_E�0?Z����t/K2#iz���J?5�0˽��Ik,Ү.�o�Lg���� ��.�Q�p� �.p�gf^$ʪXvRǑjh��wV��brO�W��}��ZȾ3S롴S; ��o� ���WZ��D����$��(�T}�f�d��()H��-�;���(v]烕�Æ]�2y���w�m"���ۨ`[�6l��Vs$�~0�9���� �Y��,��:)�l�
t?��4�9|<c䰛���B���z�����!�jLT}�jv�L�x�d}�]K
���ct\�C%~��h�&hg�5
aQ_�"q����
�,qd|�-ƞ�8����29��6�`�w?��[��0��[��(���X���r3A�mf]�L�n�Hc"�S%�Ib0gt�Pʩ�����I����UY5e�g��Z��%B3�0�7��C�ʎ�28�Q�˴*˫J��%D�uB/z4������3ؚ��c��ں� f%���H;ܻ-k�]K�L?�=�s|�u�X�^7�U��M�<#?@i�|�U`V�+Lz�y9�vM��Ҟ�$<��tۚ��UP4�Jr����IOZ���vcpV�A x��2G��Le�E�zl0��g{8��]ni㻊��#|H`m�}a3��8=�i�q6_8�;�}^Ɍ,��a��6�2����{GQݰ��2S�%O����e�$�Ug�v��t���՟Bz?�����Cl �(ݼ$M�x��|a!)����-v|��"��� �6[94���.�P��	 ��u�6��,"/6��\���9���XNY��h� ��m��������D��R�|B)��o�WX��@ 1���oꪶ�g�q2m�=��`��(z0��LxO���L��%{�M Y �t�sa9Xu�{ؖ@I���g��H���9M~	���I��ۅ�	��C�bs�s�=p&3���K
��ˤ��V($i���@���k�"�e�0E�_L��,S�� ��΀"�6����v�u����T�H���'�CP����s�vd�$�c#����'�Ij�l�(�!x��#%��y�NN���i��=T|��G�n�|q�i!�a���?X��yR�\�D)S�:�JuW7 2li�ph��H`��	o�e$���JL����p�tJ�}�,<��Q"�K1�9��[ց�/����W�O!����w��3Sz��Ql��<,�A8�~����H\�@ΊbІ�V<'8�I�]3�����&k�e���r�ƫ~��"
:�5C��6*�?�0���o̗��S��1}<ڭ3{>�nD>�%�vrK��u�Ps��?9�\�dq9M�Թ��
T��r\�8���r(�cm�Aп�e�MLs��#"Mm�� �R�pߞ�~l�cƹb/G��!b�pO}��+ŀe���f䞱��K���3����7�o,hl�I2aW��2D�%/ˊ�K�^�];6&wQp8
/6z�I����wY6�O��d�|�����t��$̡`3
�w��X,��ؐ��~*�� ��"�
ZoT��Uv��b_���Q�����m<�s���[�V3x���2^�[s*1�
��p��B%;�VmK�W���*��@��~��o8�m��������oa޺��)��Q!O�wD�J��u�K��c�[���b�5��d�,#�݆3)�"�� L.;;
2�Iq	 �֫q���W�=�}�T��JK��ypc�iu�0����2�F�Kކ�#��i}v��/���n av:ge�_�&;�7+�	��R�1��e!ȟ��\�E#�F�R���͍h���d�٨�y��)�l7_t+3����~�@�!���W,*a3b�I�$ת�[%G\츴�'ҵ�Sa��9%X�~7�;u l3��&�`��#7FI!�G�G
�Kw���A�����цU6����l�w���S8@\
�J5�-s@�v�ר�%K@n��kO3M~��C�Tϐ¤MOYIωa�+��u����C%p�O(�KZ>��O�����\ls[U����`�Npڂ0oܯh��?i���٥��T-s���

��(%�אkX�3fW��̝lZw^�Wg5�A��u���q���e���ux7���~Xw;��Ĝi�ʡ�N��Y�e�o����Z��J��g8��(8@�˳�B���Nw\�^�`S'��!zYP�����2]��0إo�oU�D�$Up�^O�YΨ46h�"�E�^X�Z(�e>�3����� ��%�>��"a<�7�x��� �:��/h>��q���\8�i�vf^��4]����n�~
�����q��5S��iz+�Qb�%cm@�%H]:[�˧�p�,g����-�q�#�A����%p���G哮�U��A��kX쌦�t �5�ڍ�s3�@�3�[�CK6��)%	CQ��Żo}�S]��H,�5)� ���/G�~��x��_Շ��W������f���[�Q�u]~/@�[�=<�坛E��n���௾W���'tz25V��
C��c�.��V���kN�G;�~�B���(G��� �r�YD��/um+3¹Pu0�Z����y� �_�A*�ӽ���&�"x:���#{�4�!�jm���+$x�Y����8��H�����I�-����K%B�`SP6��3��y�����Kdy�|b�P��7��ѫ_nǁ�
���3�o ���ZZjC�*�}
Q�P@N�J�ɿ�aE5�\?�<r���$ٕV�H�E�11��+i��r�m���c<��v,1{٫�L}A@�=�^e�t&[�LP;q?˖��k�E��7�X����W�l�o�Ӎ䢟��+�I���6�IY7����aOA�o?��|~�D2���� xcP]?��"�����>}�XE���_/6��28eŕ�3f�x��>(P�*2K4�Q�N���q+��K��q��DeNJi< qW@����e���n豾�YN(�����f��]n��ж�Ɗ�|��)�0�N���9�Q�	N�a����*14.2j;�Lq�"z���P�`�(�����_��N��@7�ے����x���\f��!�as��uu�F$��V�C@�
"�E2�
Cv^���5�B��rQ�@|<��F�1	�ђ��M;ZZ�%��h�ҋ�;/������U�Wm�c	_�I�0�F}w��dMQe!<x~B�O{�s�v�0�D}���8Kh��z�!U�x^q�H����(t�摷v�}��f�- W����*�mړ�q�"��c�q(r/���ħ�ك尀>��r�=���)�T���b�X�v��l� ����p���a��6���QK�������W��p]>��?�Vn��c7
�GǷ�ත�}�3`zp�M�UnoY�^Q��z�4>�����ik��t� �>����ɔ_�����Lum�%���*;u�	iQt��Ph�P�(9���ojpI�p������FW��0�=!ҳw��%
��봗{�*�q�1�T�gr',��Q^� �Í�� Rz������t��*|Ӡr$T�ZUӷ�̌&KL�]�v�����"��C8JƧ����~A�߿U{A	�1}lFdŏ����G�q�&�=�Q���-o-&ǝ;�7U���<��vK+Wڒ�#&�L4D�!X��B���1�m0H�b�{i�ɫ�*z���G�Z<��*���sy���֌A�[��n�5#C��q��>�~-�}"�M�M��9vB�MC������H�P���n4�(��2�����s���oڻe��;@��5IB��(15)��2�X�3��g�!У���d�e�V�N#����x�����,|7�3G��d�ˍ(��/j���p�ɲ4h��_��T~;��d.�l*��Ǽ��Jtoې  �2�H/����ŜIҦ'б�9�Q��z~����=M�B�3(����Q�%ND��3�&K���<�� �Ug'�C59� {�V	e��m����=Mz�������\��2
8k�`�����&U�=@�@�gW�������0Va=GW+B���u����oU��� 6Ǯ�ۨ\GCB����ͼ �<Zk���6��jWI��S����eMy�0�j�L�Z���n�V�b4jS��*/uP��~ʢ<V�ޘ�+���s��1�1=�G��p�a�������
���A� ��͛/X���|���
S�4)�:�M΄��,^_���"��]l�,)޳��88�-�p�L�}loܬ���H��1e��E7��	��=dt3�D:*wf���}�[�M;����o�/��cy��tb�E��R�qW����-����3���^����u��o_��k�il�";xF���#��g�С�g��+Wgʝ?��Ǡ�(���ݩ.e?���~��It��M�\�PO�=���ǅ��U�i���6�^����(}�y�@oY �z�=�e*﯁"
&Á��f�(����2/,Sʝ�w����(Tt�Z|K�L"�(`�p� ���h^��q)���2�>V[F��0�w8A\��M�}W�����)�����ဤ�̼je��'ə˼��80y�_\67����+h���i�06�1��`Dx
E���ɳ�:�Y����V;���`��	{kz�y�ܛI�p��\n�3D�ӽ=�(�Uݬ�RI���MK��J�L����9oz@/��Ɲ�mVAN&7g�����è9��fC�b�=I�k�#\��n��j=~��ϗ�lWm�zW��$��&����)��������W�1�mq���
2�Z�޹�!�S#��g/���F����]S>�����j'1�>����JI�:�Є����v�lJ�0b�`D,�n7ֻ���<[V$��lR���w/\����BH����Kh�������4NW('��r�?�ַ�{oy�?X�U�p�f�G}�$mA^��'����'�;�;��+����u��AZ�M�k饕_�:C1M�)�<�2"X���eL�1N�"�W	 2�D9�PT�"d��6|�u��u����#M�!�	�.2,~CJp��u���>#�f�<����
�c�P�ԓ=迱Gh�2�ԁq�0SX��	oE~��B�\��S�����a��}� ��pl�%Ȁ�.�����a��G�S���v����pHW��++e�)Z�%����-XY��g�rÝKie�V��H&H������|'C8�i�7����t�n߈d�:��3�����6�z<�y�#�~��c��B9�9�H���9��W$[$�*j�L���K��X���ԉ�����l|6��(�grm}ID�5�J�9[��^��a�]����?�~7�P����*�fU����]}K���4xޡ�֞��EF��e�9���m���f��OF���`j9�6a�<Gp�+�Vfd�G��ʖ~_�6ԣ����f����|���?�
��G=�l�Bv����!�^re��x�|S0"�~�A�������C��$O9��ܯxC3 X��� ��_ӬJ�LT��M��?�����꧛�h� �#s%��Yݩ�)<	@���P!O�z&x<E�*�R�0K���.X���lۏ�u<:��4��J�X�N02x	��{�~�h�������jWV����w�4l-%Ue��x4��ȓ�������G$�-b�N��h��#8���d~��c*~�+ӹo�Fm�>n�TN�éc��[�W����[�<'��Pp�P^7ٗ�t����v.,ⵀ��ˠ'��v)p�U�H@��J}1N%h����;�;[!�ي�0g�ʹ|q<~x8��g���^My@n���S*�EQs}����}�v�.��(5a�d"m�J=d/.m!��"�3·k8���z�����d�Kc/c`���t���Au/�?�
Ιz�Է9�#'3�������CT���
��Od�P�:��:`0d��K�������I"卢Kf�n�4�E(����Cړ�� �L;��i����w��dM�&N˥���A%�m|�-���pW�B��p+����m8������ɄHO�*��Ǚ,��un�!��8y��b�x!d��&����J�.�D3vqm8�7�}��Q%�=����W��´���*����D��jy$�hB�Æ6N�M�w�Ot�a������E3o��%�����y@)ڂE<�H�<�lsj��T��p�U9�O��j��q��Ě��F� t�v��A�r
?ψ���e��k�癈�=�n����$�`�{d���57��4) �C������S��!��i
����n�HչE;��3O�WpPE��p]�3(P�
��wV0b����%���?��r�%c��#mn�W��V�R�@Pz�����?&����AN��-�:�� .I�F�qqZ�±H�B�V���A�F�-]���~*��K��DZ��_-(oMJ�W����� ���m�(u�SfF�I��f<�/@Q|,p�y]�_�ł��C�n����;U��	��dC���1I���v���@�F����
��q�"��W���3�������,ʆ�'y����\#�V���H�����1��SyԸg_�x�*}�)���F7�ϟ�#
tQ�*I�^�;�sy�%�q;��̹V��q��?�T�X������!��1o�L	_�Έ/�}I�c�c`
�a�3���ūp,������f�l7� g�a�����C����x���ǥ}����]9ub�ᅻ�a�3�[��2ߔ�2�*F$ ���i��G�z9��T0
�i�|��7�
햭_EȨ�x	-e���A��*���'v�Ӳ@�Vy>F�P��Z��L*�~���<��h7��8�3�Ǚz~�X(:{���hiM�W�a;��|j��8w�e�` Y�F�f\\Z��
�f�}����!P2�v��Z��z1��A�M=��$F.�_"'�oѦ\j�F�g�ކ��/�8�N��wET^����L����t���0i�����*z�"����W���!XξYD��-�H��#<n�9��d��%�0�K�L��eZ�$@_ey_�}�ٚ_W���:$�	�b
��䧣�'���}����ʑ7y>�_��qYql�jrGa���8��vʮQ(�j�@�Nià5|-C��]؋�X���Z����e�5 N�4��d/1P#���%���?��re�JN]�P#瘷��T'nK��d���t��D;r��Z#F�7�M�E�6^��u�yT+Q?���F4��5��U��v5U�i�V�P��v����Fdj�fd��+!ރ$.�x8ml�<�D�SV�l�$ѩ��E\7���$��])W�?�z���� "�J'+s���"27y��Aq�����es ���`4UmJ�;��}��Ѧ�$�r�̭��� ��7u�A��Ǫ�-��M���i��V��	���@'�p��ԾyV�p�h���+-�Q��u�h�=]|��A�R=�9��OFR5�d�+�~+c��c@��U��Tu�ƹd�����¡�����W8�B�L��}Sڄ����	��M�m--J�'�~��iC��ۤNw;�]�.,�>����9F'#B��闍��v��h����,,�����DP��]V��ؔ���߁j��,���� # h�@	!�r=fw9R�Q�8AU_ ��Af<������H�᜔W������YW���P�,��@7UԚ�����1.=Ǎ���@.i�&|U�^��ڣ=�_`Μ�IRЙ��Y�C}$1P��ڈ)��͵�m��Th�] n n7�
^��y�i�6�L|L�����j�v9 �C�VG�{qT�b�nOn+�T~�~�a��|���WpYq
[ �;i5�u��U`+ĺ�8�Z���k&#Fsi��)&���O�Cs+�	r���u_�>:�3ȅ�!�7���}�C�⊋9����F<?\s���K��jd{fwI�]�ײ�ř�.�Uq��x��l�N�	G�� Cm�M{�g4E;�U\�-{�R�Y��-Ø@�o�|�q�m�7�'2:K���"�x��Z�����l��A�5/� �vM��B u?"g�-�w��m�4{}���ھ�p�$����)gD�	)F:R���I� ���ٌ�>|t���c�uk�����nt�~5��؇����@	C^`����6?��}0ۯm��3�gl�Ʀ�Í�E\�fr^5MnO2 1>pt'�e���k����h���Z׊�7�S,�3
{�� ̵�,N�@@d�?��V~�_�#!����I��5Kf$�j��:�䧮��b+��88����t�e@�٫ ��m^��Z����0j�����~��Ӡ���5p3�X/:����Y�u��Bi'���'�(�Q��֏,P���Q�U�5��,U�%q�Lq^��!����P\�x}A�$O����폋+P�8�W9���o�=h�����Ug�#�3��M#�;Z:���M��v���;����"�<��uQ.L��2]�,6�O@�]��砃wJ�;�-OV@*"���Ǳ�=o�q��8LܶF�������F���;��ũ�(^C[��
6��
K�,�Q�Jp�о+.^����K�sy\��=n���V����b\0P�Ys+~0R�9G�㘋���T�r̞ʧ��Y�8�8�� 8���l����dvI�C���z�df���'/��$H
��D(�9��o7� 3���D�������*���"O�)����%���~&��\�otΉ/`��Ll0��3�s�V���{%�/�oԅ�����>��b��m*�/~dŕ��v�l>��O�Rl���f[�,�๑I� �{\��UW�K�}b�t�лI�R�/��l��������gGv�^4�JM��Ŗ�� 
�e)Aܳ�v}��j�'%o���B�/�"G[����F�GP���`p�X,�y�]�^n��S{~x4�a�� uS�eh*�.CO3�v�*6̘�zb�C�ܶJbY�>"E{<�����HO _o�e`q�N0��v�|�z�.i��B=��?��ѰU;�{���M�l%m�X��b�m�B�����B��^�ۅ�X�y{��W����������Y{����儁v� �T��9�!�'�z�J� M�`B�4�>c8�����/���� ��)dz�;�mu
!��jW0t�6񌔶HdX�9Gٻ�S��(ZI�;>�6��eSk��)3��>A�}�����@~�� B�Ɓ/g?l�b�9w�G{��S��2N��u��>��	\sOm����ъ.p���~-Y��-��v��\M��8|q��>Y
���h4���),����3G��0%�4�dz��8�
�\�U��2�-	���S�aKo>5�xc������%z�zS	�l%��o�_n�X��ay�$�/���Y`��uh�GF���-[��;e�D��]'��bFR&V�6=�fاjB���3JFT��9���EÅ���|���2o����)�Ju]�/\���`N��S����U�����A.q�'s{�th��f����l
9�����'Mv|���1����hp�$�#�wEh8�J%)�?X��s2�h~�!�#��ok�r�@�I����l;������CK������7� }k?AB_��w�-w�v���?-<PC!3�_�m0��}��E�	G�oh�7�=�v���I�'��rn�*;*���Q�BϬ(����t�?��$k|56p	gF���I�%r#0%��)�pN��i65dV��ަP�|>ܜ��6���M�R�+~��I��T�#�XNϰ�E��16'�;��.*���)}����Yj){�7V��1�E׸1��a4n'�W.>2���t�W��a�O�[y�_������Ҍ��Y|�-z���e?�P&Q���?�t�B�6f�L�o�V8�	A�fN�A��jQ�� �p��)N8�&���}O+�=�c��z�<�t�����3�h޳)+j�k���C�� �Y�g��}�h�wk��~3�{� g)�d���A�Z��2��Q+�;H�:���~�9�+��(�8)!}A�E ����!]	QbvNs����U�p��m7�_�R^�я�44���k:=M���a���=~��e��ө�C3�W��R�5��ޙ��>E���d�,2�J����s����k�6���R��j4 �2�����+�ٸ�����[A��k;����_�������D�CK*{����s���of�X@��S�ь�ߩ�A�����Q�����q�>Y�>���2�i���p����C~8p���M���
�=���YA���6
N�S<��@�#@�}V<m���Ɠ���P�~_Xz#:rØ�W9W�1���wDH;-|����Ld�28!�)��6����%*���#��v��B_����Qb)qgDG�a�'`�ՠ�*��V㈮�ij�É��� jB��a�����&�ћ�����2���߫�{���w�5�`e�mu/�mG��߃}"��`���v�%5��֧�vP����ˍF�eg�4 .4�1�fwjD��������0#�"��s��t�E6�~�>�'���8@H��>r��*e�x�o�!u��v�kS:�6�t"d���3X�v�����z�� �6�h��0����#��DfJ\,8��{���s&�"�Mq��-��@�ֲ�&$Z����u4��
t�3��C�A�+2+���W/?wXw�����D,��f/,��'����|K�ўՁ�T���$1%���^WV����B o{�4~n���(ަ6�Ꙥ�"ĕ�`�8�ӯ��z��a����$�фS�Kd��:��k���=e��Q�Sa���)/\?:O�v�G��Й_�MGa�,����7�sPI�Ń.�*U^x$�WD�X�P1�?&��7��Xd�8+��k�����|�1��Q �񎳻�ʇ&ײj��DAj��mZ���fu�������v?LRO�i��2]Q�+#[k}*0k��(���T��0�7���$w�h�K�5�����@�9"��m�rR�'j�i%�o�8-Si$p\Iҹ�C��1�?�+/ޘ��e��%���W�5�ic�z���*#�l��X--I��A:p���V�%��`?~b	�����-KlH;F�C��koI�s�)�{��I<%�n�wn�M�zd�}�w[U�1�:|��\<��,w���"Q�<�5�9σX��O��fz0���wooW�m*q6�@o�űmN�=��2f��D}�c!�x�n<�֭y���N�I��s"gi�|bD�m]L� �Q4Ss��2e-���qy}��\^/�(Q��YQ5K�����}������nlە�s���~��*S\z4�F9��t�l���*��뽢.Ԝ�_Ѭ��[�S�.��v�o� �.�҃;���!�t��ƕ��8�����$a,G��Vf:�IT`q��8�ҳ8���ٌ�3)�h"�����Ц�ׅ�o�rƛ��r؅ٮ�I7�mZ>�5�=,p�-Q�J.[��@�h��ϲ�}NnK#?c-�hћ���]�d?^'9,@	/ �J 9��A��'�ra/#��H�T�=��SLM�J��J���eI�ٯF(���g�Z�	F��h�;������\�QM!��^�Z]���\	��{�'���X��m�m'�)�<Wf�@T��;�E *߱�s$$��0���L19�(�	Rc�Q��1t���VF�b��6[r��5��3z�t!cj���-0�}�鼵���H|Üi����Vz��/��<Ec//��Ȣ�;.�]����a�V��ݽ���K�	w�t��8�>oC�LRŕ-l��-HMQ�!���xX(�{���edl���Ϣ�vC�$~�>T�?`;O�=�8��EY���"/��W��7��5�?�3X��Z�~��j1K�)|��Ӷ	M�º��uӬ��W�@�;��S�h���"��Щ{a�]�N����g�f��5G�" ı�.u�>��U�`�W�&��5�|,m��%�^���Z���D��h�p�i����U5�ߋ�v�TrgP�u���� �d1�m>`�"�N�:�|C.��`:�qrƤ̷���E���c����<s��Ð��D[��y�������M�R�U�@|��g������I%�N���#���7�j��RT�pLg�H��u�u#���c�<��&����&,�&���N � e���\�EX�P6yJ2
�i2��~G�G��$�w��\/iL
�a��no�-�M���Y���%�~PK��;U>*\���B!j�$2v�3C��fX���*A���<`���zE�&
wk�X��&���mҟ1�
yqH�
��ݎ���"�s��]����;���&'�:��]7�aҲxP�Q�cǥ�@�Ƽ2N�����d�I0zhل6q�r�`a��)��s8|���7Hg��v}8�N�v����8='�WL�kj��J�P�c�DN���pA�hI��o&y��X�ss�t�|�����GU�L���2ѽ���A���.�/u�0��G=�0�rM���CU�Q �>�}��Y;��!tiژt늅�˩��z��}
i�W�-�rrw�Z�%Xѿ�o,�.J���2P�=p�>'93J[D�;i#Kl|�j��	^J�*�1�cd.���>X�"Q�3	#�R�����煲���XGԴ�dpU�-����5�^w��6K�x���Ԭ�w]O� 8c�sÊ�b��t&{'���l���Sp.��g��@�,f���Lܑ��BB2�fR��17UZ�:!?�R��āy�z��9G����*���՗RL��h�\��y�V�gluz}G<��QJ� r����Q���z͋FM�rך%�BP�ؚ x-�I�e����M��*�{{{{ދ���)k	��q������.M$���5܄�u�J3m�^v�sB�-E
�� �EV�j՞ry��O�3�ᨘ8�rӝ74/:%j��w���#��G���O�����N6����>`�d[}�o���k0��\h�NZR�'�F%��Ϋ����(KTC����Ɲ���Z��F�	�}�u��ۊ�}�Z�_*��&������Fz�wA���@LN�gр8ՙWA�Ң�:����vs����&�z	�S5�Cl�na��w0�~���b��_����a�G�y¸39�������Ӡ�e�0n����=�=5����(�B�`��X�D�/7���s���|�1��i�3[���$RP�����C�O�wC3�'Y���)S�v��r�"~����7!:X�J��å�>�.rx�J5�m�h�N�>�C��}��R����>�������j���X9$�,���7�z��j@���DQvh_�A)Q|��*CΈ�#���[����n��}s��h�9�SIj�-���"���|��5%�k\)Ʉ��8>���>�A��vPRn
4>����&�$���c���L-�P)#���S``��^o��T.�N�eq~?#�D��Ww��d�N���r����i�1�EWq^_�U&/6���g]�!�X�+��Z�K�į��r~�X���P/����..������NEmm�����͊t��J�Q$X&�Z��&��c�ھ���ye��*�VqP�~��s�*�?��x*0CBM�����b�.�1�y$��Gr�J��-����cEwe��Ņ1����%ȕu;̊��Jxy����@��)tŴ��]D�s���f#q�E�a�$@� gy����=�&�{S{X\%�7���@W�]ece�.A�Պ�G�j�%����*�Q+[��p=mo>�Nh��!ΈcP�����|��56�1��y��ﰩ��^�p�˟��Z�����dR�P8�גY�� �?!"U��[�,]I*hɃ�6���Ş�6SR�XUj�)v��i�K���AZ-3�� �=Wv=�[�z��E�"���9��na�ߨ��t�����/Ձ��"��b�s�������sKc��ej\(m�F%-v4ɯ��Xi�f�|cϷRl�@���	��F8�1���`�\�<�dwo��\����N։4,��A�DO��!�U�0�+Y*���͞$���M�2(S��9;�U�	��%L��7�υ���G�0�S��_�OL�b[{0�Lfx�H��Xxq�,g�+�a�A=���*%��?�cO�b�9����W��乥�l�b��V�����y��<�'�|�����@�E"��,ʡv��y���Z��͛0)DkcLN���ӑH'Z�(�K�I��YIknc ��i~�r�Wے/{l�[L��?�NE�s�#��5-1q4E����	UY;�ث,i�HH���2�����-�s�ͻt����GF'����[����aк!]��.Wyɭ��%���E4��'�Sy�Vݯ�A�ab:����$W�Nc��Z���ߏ��˿����&��o���}{�@������BU]���H����N����\��q�����ֵB����v	�;֎�0�i%?8�+<�K�6�BE��4nZ���D��6z�T8��],��>?���4$K4&��W'k2�i��ܐ6��.u�3�;A�Ń�x���?�W`��q�usR�=��m�H�(yN(�,�-�0w'���a
1^��A�
��GL�c:�(�5���]��$�6!��)��t��-qdż�O�T�����_&w��-���o���t���[�Vd��x=S�r��i�GJH�৥rt�C�-��$��t�|&��nᴔ��Iɹ�	�Z��_�T��pñ~[�b�U}8�?{�f�2y���}Qtx���ևa�)�bP"=j?�)�f���ʞn�[@�I�`d�k�-�C?*y�_��-�fR �����0�z��}k!p����B����	����'�4�Q\�z��jm&*��[���6C�ީ|Y�iu�nqR%!m��fW,�U: �l�f�7&�kk¨��S7Vp��J���Go�F����^y���URm��B?7�2�_*�2�m�s�y�l�Զm2)}> �P�_���z�\c<�iG.�����|�XA�2~]�S�k'FHd��y��DE�6B��R�RH+�.\���p�ѐy'ْ��r���Z��;q���k1^dNg	p���V�g�?I8�fp�"R��Х��N�J��?���>��d�ͩB��_�J��X�O���]b�z�����#�4h��
�@#��s/O5���q�r٭��NE�����:E�
���@ Q- e' �+2[K���\x4Y���po��f���s���b	��!uw!�g���^j��8p[��	�>�����K�c5�>o���M�H�ps���He켑��$�=�KO�A�{���8N[e�}8����O�_�JT3-�f��U�Xwh�bw+���v~��@�hl������ի�dL��L�`UdqM ���w��uF'~I�y��Hx��3��Q����c�0�Ǟ�a��>23�
��Z;>������oZ��(���N����0�~�y#�~\�T��b�����Ȝ�ʈ�^c�e��j`�3��'��k��
� u����!�)Λ�j�C\=��jSx@�X)�o��2�b�(E�G[�L+>��9� 
�'���O������|m��_'��A����.&פ�8Mr�SY[�?�C������wJ[R�z����U�Tx%m�WA����	�GY�1�nUn��ї���~YLU-��W����_7�J�SN��,^���c��	@E�S��F���u���K6�����%?���?���	Q܅��ң7��gV%g�R��S���+�~F�8��L,��Ubs;��׬�W��cRr߮��b�qe��k̵q�W��48�"R�E[��.UG4r+Y]>
=�]�|�~'�@�P��퍗���g����I�}�eeb�*4 YUh^�q�D�n\��<7/gG�&��M>������g(o܌�ct���lzw�l�X0�Nȉ��w�}�5�D=F����aw�c�毡�A��"�b�>t�#��hgi�ۉ��P�����c}?j�|�Y�b?����#I����QBz�o��	������xJO~��Nnt�0�X��?��ɂ�W<�Ye'�X(b�,�/���f� �PP���/������3S?�UI����Fm���x2C����/�r���36�k_�~�9�0�RA��=	CSX��=h�7˧�_T��&�s������sDa��m�9ގ�<F�X��?ٰ�α�,��|ir�!��jh���FKiG����ֽ���&��^��D�ފ(��Ǧ���3�p[~��aEA�ē0t~~��-�4v �8������m�*i�b5�X��ȹ��HlJ�TO���s�_����|t<6�s�EaEƌ��֡�ڝW߆Տ�S`m��A�N��b˿����V53����p��z��w��S:�h9��!�*��]Tk�
�&�o�������7��n������c<��Ʈ`V�dg����P���dޢf3����B�k�H���;N�r���O��/��}Y>U��4����6�r��	�Lp&l�N����7���࠰q�;r�
-�qg'YH':I`���eLK��J�;�ĤjYOoՎ�<�)��H��q�d�J�]0��a��e�x柙�|CŁ�sתd=2>��b�\X~��{��3�x?�A<:� 
�+J��zvB�B9-F9�C��h��!w���#�͋p�����XU^=N:(Q/��� ��l
#�O��^GKq���xɽ=tZ�%gY��g_�(��C<���"�/�V��C�{;�*�n@K|H��u`h�����3����DL�qE��֌�A3���&؜�<R��h�G����B�+���rku�{ɋw���:׀S��L&��v+(����.M��EQuV@��K��m���_�Ru�y�s��O澸g�;�&�@�I�~W����{o1t��2�<�D���� n�?��k���R|g��['TF������L!|�� ��.��{��*����[��At.��>�+����r ��0�V%h��Ҡ�
��w8s&�:�Nn�o���aj��P��s��+k���2���ӥA��@�.���[�/:	�VBj~����EР�y���`�W3��V�V�I��N/zC�t��;����r�g��/�t����q���H�<`}v�a��N��jُD������$�N7�������%����	M�$A6�	������݈��W|�}���e��f�M�1F���l_C'Tj���z5���y��mN�]�h��M3�+ƴ�G" x��@FB ��R��w�Tp�?.z��qLy�$�^��;LC����(�gH�1*Vx��9��7|��~�!SO�OX�K]&��������EE���'a`�6Gq\+3��Z����{��p��2-Ÿ���3C�E%�ڛ~H�����
�YsT"j6�%�%X��L]S�M�Մ�9K:uQR}͆�̃;J -�pR��m<}�Li��f���Q� ɇү0�,(-�P�~:q�A$��P���i�8��N,8�N�+� &fAƝD��3wH�Ũ'�-m�0��ˎ|���������j=F���N,ل��BC�T�S�g�o���Y1���,����������>'�z�tȢ/�4�Ο���c��
�=5�Y'�P,Z�'��l�}/꭛�(�W������~E�J�"v��聠,�"*��d�A	`�3Y�4`
�l�&*�:
kw7}F�������)ˌ$�`D�k�-ݷ�#7F`f@~,�P�A�r��շ�{ �&�Sm⎺מ�;��sOR������b�����9-b$d��a����r��\=������v83.M*��hDKq}�M����;����R�+���1���#���#��;�����j�b����Hy>�1GD��"���_�k�  ��h~��& ����g{�_�q�����H���Tҝ+�y����xӖ��R��b:-&}k�����-oӺo��4''S�������g���ꥬQE�0��1��(܈tv+6,L�Q���(?�&��8�5��N������S+hZ5�D~�R}��B�3_��7�e�@%@���FS���Utl�u�C`P�׉��^P��{�|:�H^=���]��fe͸_�t�6���0_�����B���Eo%�6��U�����v�k��{��=���_�Ѩ0�J���c.�Q�$.&�m��4@��( �O�yT�����_��aF���BE�{ę����^��_����5w�v�j������L��0�D�egD���� +�*d��e|�Yn�b��6?^�䰄�~L�U2X-B�f����d��	?_o���ZX�e�͍�a ��n�K"��ܥ)�/�Z�*A�ĠV�o�4N��CX��V_+��Ni�3�$k�-<O���W!f�`t��o�*--�+/!�l�u� j�%�ٖ�Wj]^B�����
(�WG2�?��W�ĕ<��8��g��w#�?w��av)�;�)IA����G���7b�EpV,c�Zvn��5D�U�8�f_�f~[�
�p@�ȁn����� \��L ��OL-w@���%� �\�y;�p��2I9ٜ8WB�,+�LY���,	2L�ܩ��oiR'���<�Ȁ�ڔ<�0���;;�qxҡ"�;n��h�"+�+�(�����E&��f�n��n�1A7Mw�9r��կ���D����L�eU�����R9�Sa�~�p3���T��1��$=,@!�s���gI��N?���{�M�5z,�\�D�-��7�4���`ث��.UKy��������((�됿� �gF���A���C�>�QPl(*
�ԅ�j} ~�M�ó��Ө�~�F<��|-$s�����nb�#��"Mm�쑓OVr����\\�?ڞ����~=��s�_�5ּ�W�[�z)'4��`���2^�	B���6�D4�z�ˤ���@�d4��f�1�.��������/���P0��ݣ�^�a�.�4a���b�!T�I����A��!�S6�u�M�MA�6s�+���Nrd�����і�W��u�3Jmm	kY'���yG�L�ˣ	�0x��$�j�A@.�r�+�� �?�Rz�h�([f���N��C_痴�B��F�}��D��W���̷56툛�B�ϴl}9���7&F-9�?��i<�ުǜ���,\)~T�|5�h�m�_�ه�}��%(Vn$�ޝ2�dM��vI�9ψ3���T��Z����L�p�yu.}�R8��r�%�����>�4��[�/j�C?/����ϊ �����.u�^|A^�� �ƹ����=Hs�Q�QMf�u���bX�q�y!�i�����ZU�kV�9T�E���^����M����dٹ:���r���R��G�X��]�m<�˻���PO�u�5�����:�*zw��w��=������С�р�ɁU����K+Q������5�Q3A4�w�ng=��o�!?�i��=w��.[�X0қ�F�d10��'P�K����� ঻�g��l�2�(}_ c%ck�Z[�tHۚ�rp��۵͐!���#�Od�T�W�{2���n!����A�,t$]΁�͜��J���$ܞ�	��^N���ť�sv�C+!�Y/CXڣJ8�o�X��Z�����o_����
�A�P@�]c���f	�v�=d%2/�}̚8%��Yi�J��7}���Jwu{�Fܤ��_zf�xƟ3�����f G�ù�]G���uV�H#�!.iB�0:�zw[�a�Q�_�]��,�hX��ɣo�_N�1`�����\}Fo3�p)^���<��5w����f ������d�P0�t���.�-Z����(��]�r�y���s-��ƃE[� 0�ĸ��r��[S%1��	1p�����g-ν;��~����x$Չ�zg����eZ3;1��=Y~��-�Nxm�f�l���k�QT�`ꯈ�A�(5�l��-�4q�$�̦�T�r�;�8+盳�q�	a�c,���r>K�~>���2�T���1�袇�I��GֽPq�1*/�����4�A��F|�������x�-׶IGA�D�Е3+���J�>0�Q���p���Ǵ�O樄6[��t������ݺ�Ė@4^^�h`�R��t���XWGj�F���D��b�11��6��Y�EF,`����EaN`�տ�t�}���M�.�u�*�D���Y��[Ş�&D|�+�w���.x�#4�euaO"��ǦC���a@#�A���-
*��8�3�&�:��Q��H',J��� ����~p�T	�q������[y_?��!9Ԫc6l��!��Y�%�}���o%y��Ě�s/Y�j�t!������rw)z�&�>y�$�c��,��n�.���Ԛ�(Z1֖�F�C��I���/5ݠbd��	�`)�Q�������ۋ�U��������dV���<�As�i{��º�D\`:�G~!�|k,
{t�y-�8M%A:=����[cV����g�a���c������G���8ƹ{p��=)�C��ds9z�А56J�Թ�ތ�wx�7౒�\!g�ץ�Z<�D"�]'��#���f����|�t����.���&Q ��l�VҀW&B����A�=�@Ovi>�	����A���X�K��l�B!8��E�j**L�	�NT�dϘ�����DkU�^M�P������Ew��N�݈%��M��[���]و���!�O:�֋
�PW���9�������.��!N��b�`��潋���*�#����vX������7�qU0"���S���c����4JD<;����Z�A�6�f��n��2��~sm9����P���q$����6�*֕���gGQ��������7n��PՋn�u{R�����1�V&�u٪�D��b�U�Ґ���1<��~���m1���SY�9�����@ЦR���t��E�c��[Ѧ��t\x��$�^�%����YC���j��ЄXZJ�U5UEp�>^��������sw�#Q�t^h�iκ$m�>�i�n?�����,%�0#��I�6Bg��5'4z�ܑ�qti�HM�p�~zT�bj��L1|~p����e�{p��X�pᣑs���$py�x�1�g��	���kb��'�$WO�k�My���:EYǣ?�'h#;g�D�>��`��]�:(g���80��O��WSW��m�\y�JN�b�.�#)�w%�&�~m+�)o�_h#����d�1�dԟ�1<N��`/֑�j��U����F�YW����*
e���y�V� ���`�� �鉤lK�[o:2�1l�t)z{� �Y��\[P3��M7�m3;C+�.��4��k`9���ö*� �->���W,n	)���AoZ�����l�g�{�U�|���Pw:��S����4�	*�Իo�gkb����K����2�1w��A6����q�����|��&� ;��R=C}�B:����r��ȸQ�'�SO0�k"�U�X/��i'.1۸X:1��c�k�K��a���k�?����=X}o4� τY�`��w�}M��X^�>�ߥ�� ������n"+L0\���4�P9�,f10�C�_��D��՜|� J���ć7K���o����RPߤ�W.�����D;
�v��'�~A�Pǟ|�SZ�����(�߳�L�' zO�ٶ�L#�d�j�ީ8��(k|��I��X� �u�[Ll��}n�]�2d{���`c0r{�Ŋ�)�Zn���9��}�!����'-��
A�[rV�+.u��m�;�)r�Ү�u�>������ZG�Ϫ�-�6����b��Z�a�:3�I��wx�@׆�d��,@LƘ���ߚ��?8�)�X�q�m�������_��������r|��m^:a���{��|M�_�\�lh����w�wUĊ ��M!LCo+ݴ���mX�96v�%�t�	H���Hr1��Q*����AkEg7��Al���ǽ�I��c\�����\�x8���]�9֊Wk�0��4ʙ�/_,���e�&�0���#�Q-{�%,-��E݊h��C�36�g\�r~�cOR������P�>�r�!��r�:�f
���dk�S�?�Qw4a�%m];9�_�Ԛ�d��;G=�x�����H�$�:*��	�.[�bP�
�km�d��ɒ�.7�/� ��H�W�(˱T�8�Z�]����dO�7d�]��h$�����_��j6�yi�N� Yo<��S��+5��۴�y�v�	z�P�r�5���M$ݿ4��N������o1;���z��k�[�����I_@$>��T�z���Ȇ�Tl��I2�0����k����T/A�1���|�'+�Y�Z��CCz<V��!5\�}�	,��bY����\��(���M�[��׃0'Z��ҫAν��͒��s�x�Xj���?|�\7B`�4(�F�a1=[_�(�*2aw\�R��)k����:H����@p�aG��niAb+D�&-C���5[�e��v�ҷ�rH+���� g>CJ��f����uZ�q�9m.��[X��U�[qٹn=v� ��#t��6`������j��"�8 ��jFw�C0:���x��'Nj1@�_8��2�Ԍ`���`�9�m��i�t��4�Ŭ=���w����W1c���~T���C��EP�>���5(��M�n�zJq��ρ�f[����Cg��K���l�O�z?Jd��F5�[U܏%'�x�Z�"�&��p�K����8���w�����&AR3�t�T;B"�=+����ۗ�i	��bk�\�/\d��U�k6UF~�)��8a�q0CYq���N�r�l #Q��8��J g��w�4�o�܆�ն΢�:o��)Frc�V�T�L�3�;��+[�%����^�(d7V\����tx�Q��~�PQ��۳6�����uc��Ҳ�M�9�pSoB�9@Rk}���~G�|Ó�W��G�R��.�[H���s� /�2*п����I��4����Iq��#�)�H�2����JN�� ��,�dB�x�������O�bU��7�Ł�M놹*8g���:2S��9����R��6*��)�����mZI۰6Ić�`��y���V L�Qh-���2��s�W��4�L#�P�O���)Abq�-�~��2kv��ql +>�j�CN����/#fb����Δ>�����vG���@qr�N, ��C{���f,ڱl�[T;=M��������8�ʭ��˛���H:e�}SE%p��+�x���*���KS���7�)s�k�>�.s���,�] �;)��'�f�TK4t��������D�(�*GC;����nM�wS�]�p9Uv�(��[[�m� ߀O�t����5���Z�:V}�������=%`v��R��YT9c�B�Y�U'\�1��6B�-��}C�%��d��Nf���Y��FJ��ȝ����LY �nhQ�����`�|��m�4�#8��T�o�����$�����������y��B[(.�:i���n�1��auc�QtPr�Z��n�^�]�J�K��/�&�e���c6��j�`����T�S���q�&�&��gl��y5�N ~�WWI����
.\��%rM�=zG��g�j�c�7ԉ��W���j���_)��^�/W�hn����=����8��XZ{\�s�m�y��wʇ��p/Na��m#F~5�"n�`p$���@#_On�;F�����%��N~�ގ�/H�	��k��\U�6ai�$v����DZZ�>c���v�k��6MOi����'�R\�"H݆�ޡ���;�������gE�F>4R�I�c�?X�u��'G!g��mgV��tp��$���E��Q�nA��Q	�L���b��*�LV�Ќ͹����h�9c�~A�}A����H��{F�w5mz��>�\?���/9����$-@��m��ܐx��:	�Ƭ�٠Kk��S��z��k7��S�5�����Aa�"iv��b��ukK^���ϯ��n��`�IZ��.kɾ������()��"�mVb��gb`)#h�T�B�n��ˎ���wƒ��N�?���F�\�^���үo��Pn2����|~G9-������}�]9?l`@����'�5ƨ��K�����RFzi�K�H�I���ϐ���O�ۛ�)�U�x�`3|u���h�)�K\
�6�ŝ��O{7������C�#�2z+�v�D�{�׭"jW� Jn��K�LՅ�a�c�plE���5��Y"��Cc�v���ƨ"�Kv��J�B�J� 5��mx.<y�~���<��T��kAD$�V���^Nw�e$+�,�ğ��Ŵ��#�1m�KX�a��QN$�?��� )$Q9���9�������F�`���17t��vw�l/�"���9�T��o�#+���d�_!���[�^�䛿{�Fn$�'3�S^aq�Z�4;����ZX�����N1ڷ#�f������( ����ֽ�2z�@_l�N+��Wʑ�$	���U�����Ac���w�W��/�4B�VYY=��GBe��K�yhFN����]p�Y&��*��Js�Ε�G��C�!+����m�)]�3��pnFO���"n��B���Q,Qh�ő�ݎ�x�Ы"冩����-LE�y�EV�����2�w��*׉L��x���'��j�9���Y�����7�F^����b�+ ϲՊ&�}���.��n{��+�h�z����X���@Iˊo�>���ZM��7�gIށ�ө��.�����"㠼J9*��Ȇ���&H�m ��d����� P�
�G:B����M,B��ڪҳ�M	�1t��[J�f��ȵ�x�s���=g�ߖ+S�ۚ��P��"Ĭ�#Q�YE���(��V��L�+�N�D�qmȈ���ݹ
�G�����:O�	�Bs�7?l���Ef��,�Tܦj����"�vj!xt2��G�o>�*�e;Ma&|��A�	� �<ux˃�&�m�~����s�H�xLϩ�Zs�+� uO����a�{�8+m��H׀V���>�AC�h+K ��A,Do����	%%U�]�'�������т'�@�����O˦��*��}��7#�'SLA��6�m�kB�?|���1��eEeS��5�۶�՘= ݻ��I���!JW?OHf
����j��թ�����nSnu�Hj�ȵ
©Th���d���2Rw�L�֞�i��^[�k1�������y:�13��h�Ť���qBuA�A�r��Ѡ��M�!����#<����x�k�P���߯G��#��a���Vx�f�[�a&�K�i�!��:���=�(�(�}z���Nx������<\���µ�6��4ל��=��*e�_G�����s[\�,�%y��m'�	����S;�D�7֮�
yq\�j.������E��RA.&}��5E*6���5������Hd뇨A�YJ�������VkIn%�0R�ygu�#�FO����u@\+�K�҂���Vos)�Kq�RX��� 'u��zKq_��o���iȅ����j����X[��s��L�'pzth{�eI�,�dک����Oj�r��YCk�����!��>惉&����8��o�|tn�&�`n��H,�!]b/���V�ǉFV�n��[=�Xʖԃ�Hg���58J�,��gr٠�7���Eu<aCfYgȏ+u�F�l`n�/�%9��zp$�y�ֶH*��KN�t��Kt����X^�~��6�\���C� ��X�}?�ټ�nN��ՠ�iT3�&�R��d����7�z{��@\QO%r���6��:���p�s @UL�����.�{��A=A+f�{�V��ҡt�Ѹ������<ӢdT��)��q����yaT���6@ۣ�f�3�B�%��u�v�J��~e�Cgu�@=&|p!��OQ��X�!��jn�N�����zϝڇq�+�<&_%,uZ)7s,��7m��܍�p��`�ƕ8L>6;`� 9cAz͛�v��V�n�g�rO��r��T�yS�a�_���?�cF@E�s���7�śٕ�����`L�جR?�m��]��}W��V�?�� �5�Sì��4�ePS��5.��@e_��Ψv�k4���8ڼzE�J���,}�n�c���=��4-�J�3��R�;��m����~��}���:��w?Mmvr	��l~t
R�>��5����Z�峳��WZ�Y����
H�gN�r0���>�r���@ �~�w�t�_7��R�$��u�*%rD�1j,2A����[�����s1�Dֵ��	�� �)7v�.���A����r��w��l��96hĳit��$=��x�t鱏U����t�@�יuu\��B���5��(���8��,w��/\ ����n��6�ԍc���y>!��.c�䨁�����z��{���q�e�e�7��m㘪��	�Mz��j����!=ܶ���/��\�&�<Ȅ���aoU���t>����`�AϭΠ��ls;�x�]�L�Ţ�v���K��@������y����ݾ%Z������J(ɰj�����c:ۖ���$���~���f�$cp�6a�>1��Q�!�j7���Ƒƅ9G��I2�s�t�o��{��-,C�ژ�Qڤ��K]^��e�-,FO�U�MG���9ܸ8|���?H���O���E^����Õh*��c�T�8<���Uf�>���GU�����pB�U	��\P�x�&q"�\�D��������Q��l��2��hC��"2���5&�p-��%z��g� 6��q ���z��CR��7���,�cU�S���h尗La��@OÇ�Rj�'��L���S��X6X�2cU����s���j��(�y)[T��KľHWViGi������O�Hx�
�]������(Kv?���b��L^�(�����! TE�?Fy��&	�;�[��'w��Sf�S�v��5J��C�,�G˅����K����vw���]}1��&��x�ܮ�)�D�6��_!�t�@�Ep�e{�=ͳ�w5fww$�����K�RJyDG���
�̘D����<�n��
+��.q� ���ž�[p�۩@�J�6y�'b2��P���h'���[�|�mW�y}ި{3�����[�`����r���*,��wތ����~��ا�j�����VX�#�c�O8z'�k+K�Z�RX��x��{�՗��OsA����G�4�b?a��`)Q��e���M: �S#�+�6Y7S�ia�'�Z��ɏ���e�⣚-L��$sx��e}�x�?I:�ګM�
�� Q����Uљ�h3�h���2�j|��#�X=�ќr�A(��v�#_�8���"��@��O�e�����d����3$l��W�� ���5��,^���8��%��'�RǇ͵�?����]h�41�?���[�.{`_3p4��e��g0���n�&ͱ{}��U��g���W�QM�k�����u˯\�j���0�=�u��Ѐ~g�i�|�^�^���Іu���
�ߋ*��we�Y�W�\���/+�N��{vMO8���:��6��|���ǭ�e�
Zw~k���M��镔Ɠ�jj�I� ׄ�1�Bw��7}Q��G*5�:O���fѶH�ɨQ�zj)���'˝d2�/K��ʬ
��X�����Jg�U۠`�G��v��(�	d��,��J!!1�xx�Ul!�	���$ʐ�o���":�F��w�۝�3�
���RkPƢ��j��K�Gi�׈M�8��L� /fL<m��ʚ�%��������z�j�{��x�fr*rZ�d
��M�AK�NT�dB��^Lbͼ`�
���K��+�W�$����k.����G�o\&4��ch�2�*�v�21f�L�|��k�O�i�0Cc�no `3i&��'�*����sZ��\:1�WP����4�U��� < ��LK���w�/�U��T�F�9꫱ A1E�[��p�h�K�"�OBmJ�>Zv
�'���0j��4 �0���SN�c�&i����I�9E���<�`�V���m�j�_�H8.#P��N��"�.����8ۨ4��Eqw5j�'��+���D��>���,��K^�[v�t�橵�a��Z�V����VH��G�]��C}b����_����v瘝��MG��`4�Vq#IYq�U!��l5�*W�͛�U��P]�Ԭ�����g�%���6i�X��=�{��{�VSp��X��-�S��Qo�6���/�_Fo�=i>-n�'��a��¤kE$s<���/X�9��ɂ͠�L�0�7��̱	6�*t=)�Pk�=�G���Py�t3A�/�\���}4���P������)��>s����T
*��_t�u-��B�M;₍�z�Ws�?u��t?{&������L��T#�����w����i*,�O��o3�~�x/��[�v+$���juzաiy��3*����l������r���E�fB� ��Ng`�R���69�+
�o6#�<?�g��J@Jk�=��g���l�{�xϑ�d	�����j7���!�G���p]��s*F�B�9������1s���J�ĉ��;����c� ���xB	J}+��Ì��p��X3�/)�P��i]�.f9$'��Oa�o�qk���E�å3%�bfAp��|j[�:�>ɶ	;S���!����t}�
VeY,��!�0*��<�l�G��������Is'�|Mټ@i]/�D�H��ncNz3�����ݜ�^�Lв�|�[����@~-�-�}�vX%�p˘e�,�����r�"6t�f�?KCR�D\�}��N�"�I��X�sf1�C��K����r�o�T�P-���O�2<�f%@u���0s��gpF�t7:[w*Qc�<�X�ҩ��.��.��ן�m\1�DG�hse�;m����u���z�-�����{��En�1=��;80�eU؅]"F��R	L�lt,Ȁ��K�	��|����������'!?r�L!�p�ݗ�=9�K{u��H�N2�2[�N���e�!اz��7��,�_��Y������ۗ���蔿+�+4a`��0{�Z���~����a,h�]k+M��3�#x��J��B���Fɋ���g��8��;s�}����I(�5DYq��dw��4�m붑�]���c��!�El��X��4���ƣgG���Iވ&.� �YV�yՁ�RQ;'����E��l2����66�ळ��,��[��3�ת�ٹ{zPZK'Ic��m�<���]�0P6���g�ŵ>��!�r��gH�s4��}`�p��By��DP�j�:�"\7ߒ�������:%XG���a>��CCNt{�x�u��y�kV}����DM�ݢ�Zև�����Ӕ��:H��0�8��&1�Z䉈Ì��t�ۦ,)Ƞ����3N�v�{+c[�ҵ�G1�!�	�Q�Rnd�̹i�Fk���.؛��Q�6�r�p�J�ȸ���いi�_3��SoC�\=��⅚5��6�����aL���6�wm��Q�j/��*��O�u}�y�kC��P^	��{��30����������OP�{de�G����bO�CN�+h��c�p��,�|�Y��('�������w�
��U�wu[/�����㚔ʘY��X!XYp����k��'�%��T�ðn
[GGѐU��c|:[Z�*�cє����t[�'W�f���`�L<��01�Ϗӗ�إ1�Z��z�kOY��q:��IĸB�J��89ޑ��[0�y���"вoL遴D٤�&��	D��t��4;�暴�CTE�D��4�񱠧�M�a=�ď���:����+���a(Ǽ���C��%�IP&�k�W�B��^�[�Eq,U�l��8�+���%����gʫ.��d\�C�'�b;�.�J�l�{�q���/�N��\�OU亠4k��B�����v�"{$<d"�D�����Yq<��X�W	Q=�f�_|cκi$�N'����#�/s�i�q��lGII��Sc{i�3㮷L��o�F��b�ԯ��!\FD�kh�V2��9H�&���@��	��5w`����Em��e��C��� �h�V[�(�1+�HX�U�,Q�᯳C+Dc�A>��kY������?ȥDG���A��Z�1�5#I`;L�p%���
��ww�m0U��j��*&a`�w��Z�
Pס�vd3'[$�׳��X�|�"�4L��1_o�0��8��|����*E��a�,�\;��C��A�ZP��tٗ�X���_9"�l �}<O{"�t�%U"꧜��A��S&	�8Πp��mk܅��$���Ϡ�i%�O��Y���̂�*���������C����3����Ѐ�]q&Q���[���%$���Q[)� =�^�Z�p��䮚,pi�Z������:y�F�F{S��r/5t9�
��*�; ��4��ɢd�w��e�k�� !�LM�a��.�VR|�����]�r;M5��]M�%��N>!`o�ѫ:��YG]�/��P�T�kA`��j+�����K���{Ϛ���樂��͙�����~��X���܂[��7F�¨���J�`c��rQ� �R��d�9�ˬ��_Q=c���K�1�N7Җ��ZM����E`-�I�m��ӫy���|�W�W���xp?h2�H�`���_,62��J���v�V@@]��m�+�кӐ�Z(.�m=�BTܔ��!B��)�}6�Y~o�[Q9��;+�D����3����/��#l�0!,*g��S���3�FN�O����*A�� v9�RO���9s���E$� hY�����HlH��~��H�Ws���jqd�1:}ME�c.�S��<o�s���'�J�k�y�����t��N1W�}�|!D�i�a��i	�G�G����1S�Թ��Y
�Q8n_3�p#8�kL�DP�����DIN4K>�X�����͍���QMc)���k���i7��3�h2�e!��"��/u��1Z:x���SR(�ҵ�K���l-���XT��§�������B�]�i,��~kוN�c����
0Rmt+���rޛ�b ��a���ʡ�&GDX��܆��s�Ej0��ܯ2=�t��U��O� ��e|LQ�&���/�B�v�;�L�:aޯ]#Ť�Wwo�-�Z$9�0��S���$g�eQ��0嬖�\~�	��_���A�l��\�T�-�οK��ł+*@	?����Vֱ��ו��or���="b�|"�+���-p��M9f�g��u�+����/�_o�=	�l���
wm\%ptI�) �P1���
�XD�D��w�lXjPM�c�^�n���F�j��􀄋�,1NA�'0
$>���U�J�T4�>����v߅�G���YEeo��秈2�n�l	�F��ۨW ��5�A[lI
#h��#�N�XР��*=�v�.�G�۵�*$�].��i ����#}z���wee�u��۾���=49C���\�Q����}����V�����E� 2����$)��LV�V
�%�·�)�j:�d0�엃�P��	ȹ��b,1��X�3�������S�,i�U���C����-D<��s���J	<<sXI�=��Y{�1p��. M� Á�M��q�-WiD`L�o�b#���) gb:���N�AsQ�w��+"K�7,Ր9G���֊6�����k͝�Y@�?�3s�� 9W�NS�v���5���xZ�����_(ƊB��>���~����*`Z!�'�IQ3V�����3:�	kX�ƞ$g������PSxM2WV�ķ�Ì���d-}H9��aX�]���eXz�a񣕍n��`D��r�"ǭ���ǙX���h�Wy\�D�(�R2:3���F�X�t�m�.w��Y�3n1��o:%_m������]���g��>U,ǭ��-
����̚������,���bH�pH��V��Ql
j�k{�Lqծ���|ϊSy�A�ӟ�i�6(Z� 9�?�;�v�_�����$�Y�*�����aK$�DQ�d��g�N\��U���j|�����gd��c2�N�j�cd] �y��v�*���T0ڠr��w���6��V�ӏ#h��c�OZ��'�8%Sl�E�>f&rI�"�eQ�ļjo�q�a)��ւ�2c*����H�V���5�6�����W�7�����0�Sp��h]�F�UT��D��ХG�#"�?�0��-�}��*�yL8c�ܻ�v��G�Z5�!�m��g�T1��}�c&�'�	F��P3S"��Uj��x�0�p
�t�׊� `3�b��kE�a����کYq�0E��2������Y��+oDo�89��B,�F "Aò	��q�A�^�c��/N[~��k-〰�0�Ҍ��D�* �WQ� `�)�$/rD"��'�/U
��5ʿ�1�vt>�,��a��`y=���q���U����[@����u��C�G¥H9�/��$I�Ewˑ��C|��A�M?�SJ���Kk	�^�m^%�?zj4}��>c:���A�����%��>�|7Mꏏ��z�ܐ����E�
5�~�
\W�U�����"RWB^�H����JF��ג�1��J�u����pNNGӄ��cu�J����������n����4�/�"sd��+�Kr�h�\b�t�U*���������vE� ~��g��Aj�ї7��0)و��a�E��A0�����['��ȯ�y�ȓcɅ0~5��R�{������^� t��R��+��=8[	#1�[>���[�o=̃	u�����<���֧�.p7C�ͮV��m-���[s3doЈ�2�GRwS� ��Ie^����;>[G	�fA�:|�.3�H��0�����!�5q����{�ǹ�WD�Ⴀ��٣]����(9�j���8A���͢�FOKb�%(r��~���Z�ו_״ߧ�������s�њ�m�Bl�d��.[�Dў��0��"�ƻ=��)������Vd\^��'q�������
[�`�֍>npz���;�o��;oL�V�m�>�Di�1�<��{�$Q�Ę�`��!�{ax�Aۯ��lbgY$����O�Γzf)l�����oN����p�1���Ay7�P��n�Cv�K�;�@�1�C�P$��њ�
�|�P7�vo�8w2�>WL|�$� ?t���]T��c�Ģ� �dZ��KI�a�n)��")�'����y\�ot`�$�����gm�䝼�Ygџp�LCY��+I��F+h�>�Q�Z�<~��(D�y�8Yw������/p���9�G-�<zg�9L�C���/OS��y��+1�D���z}����;�Dl���C
fqݎ�H�^m���?���q/K�~���9��_������0�˯�Av��Xc�����+�R����#O�a��PDe�����k+�H��{t4��N����>��h�k��奚�V����Z_~���8v}�%�ad"ڡ`�RݲMm��&Ri��^s˟U�ې=E�z{/p�N�PKg��:�z���@�Oc���X�n/$�TiVq���g�(�>�O_���&���_��1.I{�wfD��5hA�b�|�l����6�YګN���Pݬ����Y�E�al��c�/��$�p�υ�A��H���� WZ�3&9ʎ�	!�|Gy�8��$�������_K��/4��M+Z_�ዯ9��OL��$�J-I5~���)ݜ�u��4|�Dk�e�����k̞G�X����M�]��������r.	�\8����h���O�'6�P���lp�L�A;E?�!PEn������{��n#2ï<��Zֽz�&2�C�~T{;�ьe����}�N#핢 �b���k�,놰�*N��Dʎ��*�K|�05��/φd�� wJ|�F��6��k���
�?u��G~�c�t[��s�|"���Z��\-Y��� �n!�����s�7|U�1d��:��>�bq:٘B\Y�O�j�
�4�mVnD�Z?z��B��:��q8���i,]-�|P��%!)�0�u߲��D���	�e;ZT�H�(�E4w��8 �ـeњ�b�Xz �.>��W��I1,����� �]W�Ir�>��>]�aEh���jі�>��M��z��)�F�I!T�ߕ�W#�͙�ڥe�0_���y*���~����ڼ���$"��uA��֣��Y�>�W<��R�ؽ�E�eygZ�o%��).�u�Ï��&y�HJ�j�'��sV祾�C�����!�c��d��E7q�6��)����4�A�W�>�k�3��mc�\�Rl1�!�U��Ĕ����R��[L6e]d"�N3?�h* ��$0����ܑ�ݙ��te���� �v������o?���ȼCSN��w�f�CD!R��6���o�D��Q cF�x����Jq�K{'� il�6��%�=T�)J�wdl�V��!��q9u8wC��l����ǫ�uq�P>�V����t�Dw�6h��4q6�P.�+�b;}mH�F���P��f#8��B~dT4�ܰA��j>	o�\�� �6C)�ݒM�#�
�X�����v9aM�\Ы�˄p;x�)��X�p��!�~������R%��O׽4�O�I��jH'�G�R�c�q/�E@�U7E�<�mY��|�$s��&�蜳�K�@��w��%x�qX��$��G�p]2RȴĊ�Z���g����~:���X:=�&5x�-[�#��8�V�m�$�G��Hڽ1�xƪ��%t�?��t���͡o3e�g�8�=�<�p�Ő�[�1�23��	�5���[Y�p{)_��`�6Om�mR�ν��,�3,�Fx�nݕ�@>�&������D�ҏ�o�j��ʭ��ʹa��k&�5�?9���Π�i
$<��zPhZܥ�O��}�q���q��q��(;?_��7�	eC���{�Ӹ��a
|�f�.���i%i��ů�i��BG?�7:�W�@�������ja镼�d
g�G�śk9a�
���Y��#�j�C�3��{ ��KU$�&��.���1Xdn\�����=�q��[|�*Xϊ�9�ϧ���Z��}�6د�,^��=�t�ڝ�+TB1���8�7�g��s;Yi�ꥒ;�#��:�
Dr摵#�W'8j���ݫϪM�Z.ɶ�6L�oA�@rTi�!݊�Ű��b�+�[84iA�Kl|���f%�v>��v�F��8�1�r�?�N!��ɼ��DF��䒂)��q҄�J_����R~5�S�)3��ͽgrd�5,��-���2>�� y �`>�-�.�RP�+�fs�_z+l7]���'و��"UQ���2����_��hp�O���<]H�.~����ɀcR�̼Z2�ܙ���)�f@�b���C]%�MR9����+����/���*~V�6j��ʧv�ި���ar�M����&�]��O��H�����JhX�����('b�V�@4��׃݃�����u���V8���\6��p�S��x?�� �5˱�xv�p7��W��k�Q~н�[l�j�h��K�|P�Ǘ�
{�\>ˈc=��G�ְ�����uz�\"i,�;!�@7�f�.��r��yU|�/ye��,�M������!�?-�#���쀥%�f�x���BQ>��C�>;�%nŅ�l>l�vr���b���Id|�,pX\����8a;U�
f�*$��BRX�!+������Q�?�����=<�BWM@8V5�a��b���"���F֤�����I*џ��?����^�'O`z���\��0�(Ht��K���rTZ�Tgi�k4��������`ʷ�u�H����Vzݷƕ;Ф�1	�[�u���1��^z�}[�m{�M�s�'�$��H�
����C�����"z2L�&���h<2-��� E�,�U/<�@!�[T��ȚѦa=o;6)��3ļ�������kڢ|��i����Y��w2�$˭L�qnC��&T���@��_U�G8L^w&�<.��f�zLs�Q��`n[LŞA��o%4�b
 ��%=�KH�QLz�n���<�+wrz�ֵ�$n(���>��Z=knt_�(y��Y@#���y��OI�o�}+���1+��1�����^�g���E�Ej�9Up�����ê)�)8�b�%��i���i�D�Gk�M��Y��4%^�@&���&�6(C�O�2N~?C�â.���4�~ye��A���z���QM�H!_dL���,3�ꐺ�B@������ة�[��f[�}��g�������o_aۃrzʒ�k���n��WTY��� l#��EP��1Le��i�ލ�fq�����p�4�j�kZq�m���4̰��{�P�()*YI�Y�"�H��Q�ʕ&�'.[\`?5�q�rG#�b%�b�����a{����D0�DXJ��۬8��&:�ýùt��P��Y��<fU���[�.���_6�H*��T^`T~o���c�ǎ���(�q����&�]ݯ�yAA��r)�[��f`�C�nI�k��F�s}��z��@*m�#�B�p��j$33"ylʡS3yj3g�{G� ���;
�o�&����ɷ��[�6;�y�_m�3��\���'j���'��������v��P7b|��x��]��Z�#���o+h��t���T�w�Nk�x|�	�٘�և���&�G��,,�W��q�6���]:V����Թ%��MYl��Ф'�:x�:VDn+�7���	 HN�a:+���d2Aּ}	Y�Eb$O���C��ө=��"�y������(Ģ�^bl͗���E�vi����+]_^~�aX.���1�
fo��|ǃ��rĉ�:cc�����Ì�}�#�f��;�%�qԥ�Ɲ�c�ΚFwUUX�I�������+������4���H-�Ն�i�,��sw�{*ǋ �
���}���y@׽�2��h�A9�5�y_y�|���������$q��gl�T��[X8ڱAZ���f�((�H�����rC:���P+ŋ;"p&���O_���0G}�$�5L�/pW�?�C݋�Ud�i���ŗd*&�@�	���vV��%�/o����j�'&a��N�+���O!��et��Jq��s�G�݋����7��ЍJJ�@Ȟ�($���S���t�Dy b*?~v�F�y(3'ɫ�ӗ �6�h���:���2C O�TiJ���~�wY7
0�d�������w��p�m�qڕ��� �_0s��Dښ�����p�!V��"� c_��~�SIp�^��	d�5�G�эd2�Hv��<��2ҙ�/�������Oa �~��/���|#vf:���6��&<�����&�Ч�~]�OñWB�5$�Z����1�D�\�Y�
�pZv �ʉә-���f�|� ���mZ+l �:X������q����1���l_�Eʀ,��@�$��g_��:�V,�)�	PF4p�P��^$r�Ϊ4GY븲!q�(k��gYf��̒�)W������A��ܨE�޿���}C>E���i��Ew�U��8��x�2S�ADfPDu�1[�}󇃨-��K
t�o��`�J��^���܉�'���.��Jv���##������~��vf��^�X�nl�\��(������}st�+
DFj�=e��#^F���j�ٽU�T�%�vK'a�nd�C8�fK�..�E��.�G���I�L{��ꢶ��j0<��n6�XQ�C��N�9s-w8*��U[6��k�UX~Ș��@���p_GǢ�j�=i�I��,A�߯0�!�IE����տ�����I��3�d�j���%Z�<�[��.+��I4b��:�2Ƈ��ۚr�O�KI1�����t���!�bU���j���vR� ��e��;�O����u.j��e�����}��V�� HM�+s���A�n�J/ӒW�e���%^�@�Z�5Z�5� O֬�%��7�����ƛ������������/�	x2c�ML��
�4��vԕ �r�I)���U�Ɖ�a��ZW��鈌Z�^;�W��ʠ���G��N[<+Z��[�&@X|�s],T�>��f#HNs�d 秪u�_v֎F��Q���n�q�g����q��12���U�����_��&}�hx��p�|�\�e�f��|��pԇ���F�^��9DT�CJ4/ޢ0����rŖ(�e�;�ε�n;?W,œ��6òe��؞�h����,؅E��,��UN�V�������H�Lff$p�q���fL��o�-����L�g���d��o�cΧ�%%+B$�+K�k��#JE�N�!m{���VX�h>"�V���}v�d�����y9�P���(�I���T����[�H��t���Y��w	��c����&�u�-3���Y�9C<W[�r�9)��:��F�w��̱��n��������47&��a�ݛ'%�M�8n{��7�yP�֯����E����$�$���u��@���n�U��) ���0OE��'��UY3��)�\'�G$*Xɣ� ��)���	mL}Ҩǿ*�Pb�Ǎ,ՊK����o3X��7�&��M$A��ty����G��<d� �S���i" 4"�ZW�Έٟ��a�mQ�qo��H��ӈ}#�v��˲����u�sc��2m%hn�%��^`����M�,YQ�A����<b�ZH��h+��������"U�ʥI�+��)��4������1��q�����Yρ�Yeh_��$Bp��Z��~o"�*�������Y�B]�2�?�#�q�l��������[�P'�,r�N�W�vJk�[���N����@?�Ȇ6W��� Lw|%8��ד�uߥ����Ў�(W7Bi%�+�?e�$��5G)�6��}��?������	@z6�&J�`����$�����;�?�[���,�?]��G�w�$�4�9�4��QK�m�>�����A�DV�Ax�b��q}�К �P2�1.�)l��1��~�H�T`+|�32CeSs��X�!�[�ɪr��Q�k�Z����Yw���ߐ�8^���M�+"+%�!���R�%V?��{���̲���t�D�ZB�D��=��.+�I�E�*%6<1�M��-�+ׇG���w	[8����E)���>��0|�+bUF�G�MUƜJA�K�);gc��z|��h��}��I�Z_w�W��8T�lg�r.˖J�!H�c�tG[��9��6���:ޝ�e����k]5�Y�wP�/,���#����ܼ\[{�Ѹ�KE�����1lb����Ls�[��$�ap�x�����n����榽����F�p^Z��]
ᡟ�\?`�pa'�\�Ked�ߟ���-�����Y���-]7�q��*�j��|�a@']��BXiB�/[3{iE�"�B7��6I�\��w-J؍�b��]���K�\�/���ibO�X�m����4��+��X�K�7�L���A��ȸ��GJ�,|��o݃(g�e���9?�L��0L=�bsq� _>�8J�]��E��*�Z�.!"Nj��%��%5�Z B��^��H?
�%���EQ���Ou���~?�'�1 ���[���׌��k�R�o��݌Ca�����+j!:�õ$[����y0�X)��|׊��-	�����a�.�1�GA�#�=�<�==c��������U3�-��S����%�QH�u����M���qf�2P��fj�_��Q��2h�\�z�*�|�{6/i���6f�89��l9NS��������c,��O��f����PW���X�ɜ�jZ��ػ�?�'�T��LU������o���|H��A�K�pE�/R��N08<��{
*-�\��d,�`�*y��,�w��d�N֚�����{u9�cػ��0aBTo��vM�4��7����x�T0V��}#�+�u��k�گ��T?ɵ�瓍��ѽO��f�����0�@�ӧ�����X"T���L�)����Gv7�fJ��ؼ':}��Ќ���#�Wi_�d�adY��$	R�/�b�I�%,i�r�Q9���N��8��j��$��H�y<`{���{2�[�N�;J�@�E�v�C]��v>�iG6Ygٞ;M`qG$e3KV{��w#�U9D�/;��o�#��.[��@�#�z��%�3rm�'!�(h�|�i�V'�߳�L�ر2��+a�T<���|�R�7@�@�8�s@�d��}<蔗�j1d%��X��P$:Ox:i�ۑ� _����V]Í��pb�Xo���ycyd�U�pic�W,���|D1���5�{�y�6��S9���	4���/�}��������V� 8ӓ9�q��~�2t�t�j	jkx~La��W�.E��D��68}�`~���O��/��r��<�Ԯ�F@W�F*�K�+��w܆����ދ�XKa��Nد�������]�:�������3J�(�H%�_�;w}�>e�]�	�~�z��j�Ďj*p��H_����qo�7lz�E��Y�J��^�����/`����1T=1�����C���n�V�s��ա�R�9���7�?3y1'����h!G�m�i��,p+�C�3A�ݚe{�8��q��s�����c-���5Ծ�����aM`�2{zC�I�?4K��>�a<���Uk���{\�}���`��́�ɹm[n^���^�y\�����,�2�b6wT�˘�B�!l.J^fS�i(͛��v�7��g�ϐn^KFna�R��?\��Z\�:���[JG�����.����߸�y0��� g�,�1�ſ�5��O��[SO�k�+?�i�����<���G.���M������ �U2��8�	t����E��`�jaB'�=Zx��D���[�X�@���aU�r��ͱ�'�����o, ��*a� ���C\b��E=�j��2�XO�)KaW
K�.�Y��!>�R��C�9n�|����������a$���͇�#��������b%���㴝BoZ��7�*yp���ϳ�?����r�.����FwM�op�T#�6RN��l�0�GL�%��P��G��4��s�̑2ͳ�y=��#}����c=ts�W"M@$�\})�Ԑ�, *{yv���B�i�+J�Dc_��L#���t��1��։��������{�|D����t;�֟�&�p�t��,BZ�vf�N0��n1�M�|�\�5��O�Ѷ���Μ�@�Z^����������N���?�]U��z���j�4�y�p/���.��U�%qbm퍞˂�ǋ�80�б$�E.f���7�MXY���U~T������ӏ����;���Sʩ����>�X+igP���|��=�6��"uV�8�5r(eՀ,�x���>`�Q3ǅYq^��'�ʪH���T����SH�;���S�I�K]���L/)�Q�h)۲�%4����
�aM�xO+�䘅��+j��m���p��tK������	!��e��{I�h�8�����l����t�)�8���.o�mpn��`2����<�G�^÷�^Ik�jծ����8YȆ��i��-]�}�FRg�O��/�~�9�D�xv�T7���R���G"?�>�o���8s�] p�����#��'&r	8��{�.Q�0�l2S�r-�V��h�x
�������BvX�X�,h�����"x�hB�m���S�"�[�۫V�͉��ǣ"G�WPdC�us��^��P��Z�67�	O4A���Fk4AjQ
�1�%�o��o��n����t��-ed4
�@x��֐U,8tV_+�A��y��D�"����7˘HD��)\�5�{��-g�.�*\?���ó��kC�J��RLlV�@��"����^��_���C�1���F����6����Q=P��i���nG��_M��p���֓<��z����u��$��,��\�*�"�5�2�����A.�\@t� ��pxR*��8�FaK���*�'���)4�BDa��������q�	m���a;��ʟOg_�3���Y�_�gU+����|�^w���=5��U�<�B�����և���1�fK�y�ȅ��5���]q�'d���A���-����(D$��7�`�ߥ!��\�]<�#���U�![�i���ߠղ����n%2p{]��+�1���[�{���Fc�/n���E��7s�2u��cW����0�SY���϶)ܙ`��9x�C)+a�p��3m��ԇ��?��L�}Պ��>Y���e�4�4E3LmP��Ѻk��m5���*l��b��IDb�F%�(��C5Ϙ�,n�~mI��Ǻ� c�"�%Q��NbF;�G`�	�~�� ��@�=�*���9g�'����-:�p9��5����, Îj�W����ΔxB/��8=,q���W[h��tT^��<�$���,E^I]��mc �|�x&d�^�Փ�r]�<�>���U�-/R�g@T!j��t�����h�g�"�������K�]�8:8mWO���#uN�����4 �ѺMb�-tH���}6���Yᡙ0^�9�a��b�2�ʠ� �m��6�;R[�4S2Z2b�"��s�����<��� ��D�W{3�&Q�� �@"2\���G�"B~�h"2�^�i�����/�h��S�e\1i�UG��L��K�cN�F�> r���ꕙ���L��s��`<� �/m>�p�XE�ǯ}d��$�$��3����`���e:�xT���{&�ƣ�V
's���?�K>W%�t����{~�j� }��@��4����`��.W�"?���>�5ב��@�@�r.���+��r�]�_;����D���	E�٠�M�RBҝ�Z4T�Z�:�Lz�A� 7U��A���!��@�$��j� տÔJ��	3Â��j~z�L�����e�0����__���j��UQR
~����gqkY@	3\��bp��M��d��	.��G��!���#�%�ikB����P&�OO�ʚ(�2{팭U��&}�tG�e'�ʾh��g҃��+�pk��qC�:���6�2оR�V�Z2/�x0d �,��(t�#ڿ����ք��C�υ;�YF��i��ա��	���;R6keH�h��!������g~�3"���|�YzEY�nT�"��n�	�������̱����K953G�[�"�	���Fs��n_�i�AM!�Uzq���:݃J�C��A���6M�C J���/��J@���i�����y̹g�]"���b��7��%/���\=�y��n�*��^�K�Е=rH�޶%$�%�����խ����Û+a��Bw�qM���5�-@ҟy���#���;z���O�B,uc�l�����e��ιnt��Z��Qx�'��\C�$��7���i~�)�}��Re�SY>��PC�=��C���"!r
�1��T�^n9����̙�����eEr��S��e���X�����}(0,酨����t�
gӝS��;�e�Ӹީx�M�i��i��/r����~^Mz!�~���c�.��v��P�^z*��БR��N�r���ĀE�Z?�Z}�9D��yL� ��|�<t����(v�@���(�/S*�w��zx]�~���ǈ:d�No8}�G���}��I9~�A��uIκ�n����vg�tE5�L�E�|4#n2�7@a�-�:��bMK�R���r���B���Ci�F�����+�DhTr0Z���nz������ne#�q��ļ�[m�m�[�`d���HԒ�C�2R�M�/���#���jC7�BM:�=>Ö����n,I@�Z�54��4��Ģ��LGV�X�I:�ǘ5��s͖�fo}R;A��
�����[�&BMb�������{�+1����7�V��o[-�
٣0)�YI�#�;��֚�y|7����S�w�>��]�$ֈ(�}�ҮR|c�;Sz�ȑQu�b�qu%YV5����$?�<s;vZ��)�-{���I虢�r�W��������t�t.٤Ҙ��U�$�f����?-|��	�4lNE��w�c���
�9���MeP�z��݌��P9!�K��r��ܰ�P�U.R°8e7u:���*�%�;�M�Os'��qߕ�iάr��7��+s��<�|p�DE��M&yx���G�������@����_?�B����_�ƨg������MfMze�Fߣ#���"FX>��o���dŅy8/��I��BKqU�&����S��+��IC�¹wn�?5l��P���@��!R��l��D�R}`��Ȕzn@m�����b��s��e�ğ����:���L�6嵷
)�*��^Z_�Ĥ0��ܑqb���0U����I��jN�����2_����Ge��R��Uo����R< $�N��s[Og��ԍ�?b6޷)��1���8��js�����=ۍ"�r�tL	�UV��+s�a��>�I��?۪U�8^��Wca6e� m�w����k��M��֝;��s�{�QB�q�Z�U�@ꚍ�L���!Y��:�`�bZ�?_�e��p�N� �1�����p�������-��%p��ԥ!�l6�
^�����-R�����(�}Y�[��/���||�Z���;���:�iƴQI�˄Q|5ށ>�6J5�ݴ�c�l��2�������.�~��:�^M韩x�nΖ��<�"�Đ~���㌗~>_��Ńns������~j/�ɩ܎E��	���)ε�a��}�� �~��$>�P��)��9��q������;�7�m���{`K��g�ch��P��/�D#�t%Ţ�p��������b�W�@Ws!�;'c��5â��Y�D72���g!@�*���)�){��ShBm�a�/�Xѓ�~�w�����ޚEꥒ*e�e�S~���Wѓ��?�RcW��F������%�>��C�k2p٪7�}�*�5����W�*Y"l�������!z�ꍗʛܭꁗ��[x ���<G��e[�!�%=¼y �Ko$��h���e�����
�%>�+{�moz����_��B�ʯ9�����.����ޤ���Ss=��%3�$S �눀T��3%���u��L����phA�mw��=����U�\��h�ث���4i�h���-��wh�2���N���o�wId�z�rDn�2#X���>�|�?��Tj;���_7�h��W�r�~gx�HnvX��x����d??��@⮚���2�U�M�"�ј%���~����'�!K���B}�ES�X�b���#�*0Qm��+���bFӍ�-+hQ��=��HD_"�R�.��X�� �K�	H��)`w�֓�CXE��%�ڧ B>�5���8��c��5��+!�c��=v�#��"��e��k�*��3�b����l�j-��G\�_-	��dg��v�b4>r�|��5�޲� X�$�1Bh�삢�F��O�ె�����3���V��çƤ>�f��$�"��(�2B�Q/S��x�Pq�\�v�)��LY >�r��"aSǞ)��G^!}�L91P���A`B]-��7D䜗t���QI�X��6%�?���Ɩ~/�L��޼�������Ϻ�y�W׮@}�9�A F���\8*�Kz>�� �e��J�q�|t-�G��?�~)��\��Ea�[[������/�T6��/��e��aD���,$B�D�;�`�=����6F�F��l��$ٹ�h��c�n�t�)^S<�8Ue�xX�OnM�W���'�B���[g�>o�p��~r&<Đ^o?uh��&�#<�Yw�6[l���CP��O� Չ����ϯa�S�HKF���A��=�P\�!��V�K���g���O�/ o,��޴?2���{V�22c!���_C�6��U�&�z��0�` �y���{�,�u&�r�\��OZ�bZ�8�_�W�{9��r#���ϐ�I8�l�B�������MT��|��Z�2�PD���y >(sk�1�B�O�3�uZF��y��4���L��]C��0H-�!�r�+�twGir�#=?&`��dt��A�^��Ϧ��^ΪB/�R�{�˴�/T����=5E��1}��B�?U�:-�3T������ u�n����
�P- ��2�]��9���a���,�ː�W���F� Q	�X�	K����7�]��CVo	;�}��s�U��.L�#>ܵ�ѣj�I��t��)�D<J�����cM�-4��@�u�2��;�'��pOF��.�V���ˣw����E�Pzڕ���D�N���힤��o�������`������
W�	���l7j�,!�m.�_U1��	�Z���|�`��X��L%P� ��`N�+O�d�s�� H����1C����򮫺�o��Yj��Ż�҃���ET���$��}^���R�h�����C=Wƈ�ӵ
G
�|$y��o�a�9%+F�S�^L�Է�c��ʥ3>�a�����?0��h�������"�h�j���"2Uw'C�`�v�����������
���h� ��w��
��2:!�m�xV6f���~��I����S7�֯yg�{����|���2����"�����4|=/�����;U]�z�{�Ψ�ֵzAg)�5��/y\I��{�&��ˬ�T��N�ظ�4o<���o�й����������c
�����#�x�U�����r
i1�_���M��%�b5��n�xؐ� lv���p�)��(y�DC^�!l���4�s�n,r���0���r
!� ��y�0<�u}��7���P�y�$B_�qǮ��������x�|��?�SFQ�©�����Ζ
ob���]!��X��J�*�FQp��8�]�R���ȁ���cn�EJvf�W}��k��!��Ωw���UY�G�q�+�m-���W����ix��ű�6�(t#���ľ�7��
ն�����z���,ˣ�L|#��e7�EMWM?��p�])9ݸyx�t����x�4+ۥO��~�}���6ne?Ћ����!�cx_�fe�LΒ��r=�y�<T�w����-�����r�Q
�VM��/O;K��1NU}�����lM����,�J0U���%׌8� y��O��x�r3���.-����#���i �\CK�*�9Aop�i�S����XЧ(ݑh�����IvחXC?���󌧥���|�bDO��	�JR�|�|�Q���HCdlshQ����<�f&��.�V�/Z�)�����Qe���,��Z-���u׉Á��e/����wo���Sx̂�Un�J?�M�ʵ�!�G�߱oO�#��Y���)������k�2��H(�iV�yovsn9�<3����P���o��{F����e� ��r�t">/]Z	~@��:�!^')�;1F��ͩ�C���&��ï����o3�D�DB A;	�F�`��M�&�@r֥̆)�6����q���h�	�	����Z�
k��|U��-&���N�!vxs���Y��4_?��2��z��=��f>1�ϒ��<[��[W?q�6�(��n��<L�(gwx�l�����7W�g�8��[�|򄃲X~%��>��ZevN��2�S�8���byw|��]��e4k����=MØ�$l0!����*�E����o�Q�#�ta�`8ج��SDM�U����G�Ê�/;�w��T!����!�_��]���j��'W�������؁�혐sa-����?{̝X�ʅ�{��vw	#P�NL�Ĺ����@�I502�t�K��b1)�c�9���'H��D�d9D��hi�x�!��*�(*���<0�"@:��?��w�N �����{#�7���ia�J�����F�ӽE$:�����8��#A&�t��'��_gn2.d�Xf����v�i�IS�r�LZl*�AZ�g�ŀ}��:�袎h*|��:%�_-GP�Y--����Y��攱L��J�N"E�W1�]�b�����'��Y�+,鼃|x����׮��R�lEwVYE�)_H�2��;�h�2լh㴰Z=�@^��V�>�[�I���Zh
[�2NށƷb����P205t�>���Y!�H��j�E�qh@�+��D�%}��z��V�ut�^���,)־�xY�
�v���,Z��ԲU�M��u�R�~�ӧ��9�2���7w/��bbRy��3���u+�#�Y���j��̜jv[L:k�p��g������
�g�@4+�G��z[��>�'m|��G����u ���Kp�~ү.?uĤ١����ǯ ��f���h���,�=�{
���3��/?���E��:��}��-���p��P�F���M`5�Cel �i�I���/�xj���?R��݈M���-ݵ�bkQ�U�N���@C�~8/�X�Б�tO����0ӿ?�K�3l�k/Ğ�l@ �jR��6?x�2#X!Q�ۂN �]:�v@�0���=F�����/D��)�&��m%E��8 5#��\��^��H�.�A|��rSP�>�$�� /�K"��sɚ}���'���.�Z��"|3��rd�"f����d�oi-1�@�Scw���=�v��&	�k�@�/߃pF�о���P!T.�I��ϙ��+y�	P�n�l�R���r��Z��]�r�:%bk����x��W�-.>������G�3�|G�V���u��.iT��Bgۀ6g��s��V#��L�����?�Y�_���k
�[d"�v�I��{G.��I?��i9��i��5/�/Xa*��eT͏��������͂�w�d�3���֏���V�U��$N,8��pR<䕵���`>�Ps��>zM�=(:O$��I�Á�RF��v]���2#�c�etYf�9(�K�;�Dt#�Ƥ��������H��ߜ{jX�K��@c�vܥ�d�.+�����ډ[�I�=��N;���H9|��{�K�tIHÆI���$���^�8 ������-F����MP��w� ~2�#7��v���]�$�M�������o���S-�
��`2A�9,KG�R�A��Twd��z`���LcMy����5�5����O�vÎ?')����*�Sڜ�{���#!�)�	���sP�Gh���6��2��D��a�C���P�È:ڪ� ��ʭ��O�!k7ZQ�����6���RJ�����74W&ۖ�?$�oe8�1CT=
v
��F�9.����e�e�㝉7�b9�/�y1b��FZ^�'��d�\3f��O/�q�opY�H��"[�
���Ȍ���\�d��թ:��Q���)��]N��Ia!��B"��37�����p��rP��,�m�8��㉎��T07�*\�!�qWJ���t�ۈ��X�ϙ|cN�8$;�<�Ǭ�\�>��\
A ��p���9�U�F����ڨ��%
X�ﰐ�Ddr6��d�|B��H��\[e�Feu�� 4j���{F� �5;ǌ��bCz̾*�4~G��D�x�� v�N{�gy�GR^4->@|�#��q�~�q�����<F��DU�Uor�e#Z�gniq-` 싨^�i�_�{�LdR�l�����ʺý1@�ğ�)��((>ev�V��n2�Bq։���Zg�^V��hKLX�%�ᴖ�I�#3����7�w��ӟ���I����E7��Yq,���S�4C,�2d�Ȣ������L~��E�Z*���U�/�<��G���&A��眫l��Z�-����k�%�w��N9�oe��:x�J���$���A`�;�t+��U�O�uk��#����DF�6#�Գ�io�9Fk3��L��trRϡ�~�/P\�� o'� ��ك� Çrv����Ѫ����rݨ�
�v���'�LQc����+�[)�ި��E)�硾�xτX(]:��?0�%�Y��]r/k�(���
�B3Cu�l?�N_$Ԟ�aX�x�-)�;�<q�bXP@���z/�\�<V�
��A-m�1����'1.TLtI+�L��2*���}s4O���_�[�E��8*��B��re�~�� ���+۟&T�����g �s��	�#H�Hx�%�ur(T~�Fߍh�)�w��w]��$��c���t�үtq��'T�A������J�d˟L[U�P[��%���C8k@S������BP�
�`BZг���F8]�|Q�_Bȅ���uw"�m����فʹ(�H���7�N��E\"�oDw��J���lثqn��\��OM�0v�f;��ጽ� ~,ei���-���L$��tM�I	I��=�.�n���xϢ <�P��_�� ���@R=�C��՜7�ܮ��\O0{��M���|+ک ~;�5��Q�c]��'={��I��yx��"++|�|��ԩg݄r`����3fgA)s�v��F�F&.ф��hHu�G������xg�R΀e$04�l���y����^�/V��\mpn�gX	xO�CG�#�w�R�[���4���0c"�Ԫ�$:�N7C�p	\`� ���-�j�����S�l%S��"U	� �7���%Fg�a��P�7@���V#A�����;���p'�PWjUX�F��:��gqa�+Fp�y�-�Ȫ��+]�.D(yWY}�����r3;�M�XN�bW��P���E�{��{��r��B\�����+�Ȏ��c��x��Z������@-�e��˴s>-��EP�J�LywG������!v*)�2Q���� 5V1����)�'F૸� ���W��W�t��y���4����Z���}�4>���f�֞=��Z�?c	1;���/�ǧw�c&���+D��n?~D`^G�s�줢3���g�U��<��N�0*7#���ځ�G�ش7ڗc�7:t<���oaJ�4�'Gg�&� �BG���E�}�G�����êˊՌ�t�U02k>�����a��wݒ݃Y!ќ��}S9N�V��(��:`�H�1t�Pe���H�^m���*��^6�}��1����%6beZ
�%w�M�t�%��^ɘ4�=�G�ղ�~���)p�\3�aכ	�?�챵�6�i]����G�е�/f�oD`�G�5����;r�S�|HB�K�s���K�[����0�4[0�%%ֲ� �CpyL���G��u�G+�b�f�H*Z���� �XI;k9<H�<��n�'����t�g$\鋕�O�i� KE>�u�V)���_�Xm��^`�j߾�8�/e�b��R�,�n��p��N�u��Q��O�2�U��eOt��w�.�U���\����\��I��ۣT`�� �H�S(����/���H*I�l�+���/r
܊^}d�l�>��L\M����~�yǁs����Q�9����e����s�i���k-�Ja�ā�q��q�<dP���P����{�,�W;�$�.� A��oXKW��A4��KfJl�7C�<K���o����-���(������xD� ��p��ps�~����%� �B	Zs��E��Tj$��,z�Z�v�[�̞�s,r{)�̯��Q?2��Ansg�#FM�Y�+b�(��6�
}����^+��4���p�˛N���j����2�C��-��6�,=���Y&�-��h�I.�ݯOL�/��/���W0��5�zф�}�[P�k^�A����@GH��"���w�������갠N�����_�e���P�f��I��6�lG���!6��t����z�)��~fU��gOo!媆����KVؾH$�@������Xv��Է^[����I��(ʃۡ��v��5�p�X[o6#�+����]e������~��[ �B�X�WJLOց���p���-�B�=�����s����)�?��:Nڭ�Upb&Z�~��"�Le�Dw�A*��"mcSn�`s�5qrU�HZ�����
�n��k��[�A��ݞ�sVk8���ҕ���lӲoOM�6d0!t}!J�]�� R5mH:�cɄԑ�(��kD����'���"�KI�\�1�h�aW�['|��(f�#"W���X��D�~�&~N�#��"V;=>���|�{�5��l��;����.8��,O��TKЊx$ұ(r��&����l�g ZN����7����c��_�d �_+��ڎ�|��DV*��'����>�ǅs�[v5c�q&���T�|S�qU�,x�� 9�Ɓ+#K�X��a5ٟ�%�Y�=���7<m�|֏{�����ɡ��*q�c
��x��3ȋ��ڼx�����"s�4��N7)��^,s��U�l��"�K0�+�1�R�eۈހ2��p/(����I~�e�&����� IF��� _�O�"9�'��U�&X��Ac�š���j8�l����}�;�����9RCv���p�	e^g�x�,���C�q��]t���n�9�f���	r������ʂ����^x��p{O ?���]`LSr5"4Ե����@(��w�Ĥ�ֻ�BY���
�
�m?,+�ì��V��F�&`Y|�*�ɉ- �l���{�Y�7$8�U���bV�95���u���S�����SLf޷坮NS��"�(��gA���i���	���+x�YH��=l[~K����/�T�{�5�m=�J:�=$�(�K�2�.�����/L�T�ơ*1�r9ڥh��B�G�n�"�(Iz�ܞ~�'����"_$k.�{ �+�	��7�̕���0��P;��"hc6�y}�Xri��B�9l�"kl(�d{4W��T1B��!��$�96�
F��a��%cL�|\��U).�ߥ��)�I�烹��^r�����K�A���	�Su���ˊ/���U����/�.��u)�����9+D��R�(M��~)����<T�`N�{�u��"��tE�@M�L""���~�T���V��p���O%M}'�M}ҐezDX��2�t�2tZY�0�=��Ւ�.[%��tu�d�
�s͟�Mp��I��OW"�C����8�^i��*nQ�-i]�%!�򴭪��/aS��������'׾�F'C6�b� ���[�dB�?n�3Y�O:�[`,#��򐋮|ސ��O{����V��%�~.`K	������AhT�
�/eJx@
�������,���sʱ���*D���k s	?��U��j���T+Q�%d١ݛ\�ߎ��^�v��%�F_Z���4}�\f�=@�X���o:n6$�
m��.�r��'�4�z_�T��p�@]�@pt���1��ʂ��i�,!�23��.��V:M��4�F�@�n�O���m����1T P�K�5:�ba�"��y��o�/���͡��+dBc"����4��m�Ֆ������z��V�9����W_V�/C�KĄ��6�3E��B�W>eJ�*}�M�ι���|�����i�x���O�s�!��/\;+&�*Z�	�=���q?VUI*n9�}(|��g,�����-@T붤D'-v�,� =��h��w�������q�~�wct�aj�I�m1��תT��D���lQE�����
6��n���d�e&��F��8�2G��p���5�9���#�}��t�E"��U3��3V�����1�]_�ݖE���ѭl_��{9	-)�-L�~���󆨪�:j�����?S�����:=!�<�D4r�J{ }^�U	�(�;����8�fÞ��"a�H�_2Z�������F�.A��_�{eU�·�e�#5����S�϶^�Y��ls(YM�4,~hYX;�K�=�����E���t��JwaZDUL�S��2�˔9��z�#,[�w��=0�I#N��vS�{��rn�%-^��c��/�FH�\��xf������r<\Pʪ�+3���L
[i�7�ܚ�]�;���A��r�%J6t�y�� �?yf`O������%���r\y+n���t��<K����ף�7��8n�(���)�$���;X���6@n���bsi��s)�JO�r�km�*f��!!E�U����S�ںitc�K�&�e5!��N�.C�Z		�X�C	�՚=7R��9�U��j��X��F�m��e�.H��N��J�[��<8�5��"�.�<�?H�F&�ۘj���=z���Io1B�>_B%�hF��XSS�H���s)�c����>�g�ԉ�Y�$Ap��iי��U�]I����vq���veO��P�#���B9��4��5�c3YYڞ�eZ,	p:Yjj!���jsE�Z�w၁��Π������(�5�n�Ek��`^wv�3�@�K�M��>�AAG1W1{Հ�Q`ch��	�����sˌF\�E��ia�`Ō�>��]���p��}��a߁��[
�˫��˷�tˉ���5� �l���4��m�c�]�-���'�8��<�7�gR޹6����-���]*�tE�����I�j7\S)��i�x��0s�#n��;C�4 �/�y�C��wl(�U�ϋ.B������D:x�l���W%�ڍte`7��(Rɳ�O�:G¾��1%	��I��2;��&�%�v4��{P���-Qg��A���2 ��]p�Q�v��DQA���)�$m�9�.��!�����W4n�7c2���©�0��80���+=�(u�L��ʌ޼��Px�R(5^E���D�y\�Cطf�/��o�̽U���/�p��w����3�^@���Qc{��vw`�!]���	� k��ATڸ���9��k�����E���~�����{��p�i�h7Ԉ(��K��K�Bn��3�ۑ������y�%fpy��U���~�V|{�G�d09�1M���\�]�/��y����8��.R	Qz���B�WY
�:���&�����-��~�}!WT�$ =녫��ÍC�+T�& �J0Xn
���-ױM�^p�v�)�ݑQ+�!:�����z<R�q���_)�r�~�Y�f�������?tD<�f|�g /f���T�r��7�l��R7]��I������&2'��涯ˎ�Qs�Zb�ʫe�n���|�vPgɖ�
P�m��
񜜞���^���>�F�s�9��05U[�@h9!�� Պ���$�@�ysu(p�6��=�Ű�>�?�5C����@ϩ�.��2�@�_F��N~�8��Q�9��Ǧ���u� �3I��
�"��#G����7BH��a�0L+o����
�˜���
�>e��m��-X�W�,^�5�l���d�.Ǎs���;D��5�:6nL*�Hj6k�	�=���!��d"��7w������b`�
�ܛ�F�i$ �٤^o�nb���):���	��4�lW�1���f4P��w������G�3(p�
hH~(�Ms ���s����f�M(� ��������C��ݯ}�vmfdG/��[����4�k{�m�\���8����G��Uk|��o��/h������8 p2����S��&��Z'BPl	�g�@nsA$se� �i|�llc�?W��q'��S	��]8�
����N���<��[�j=�C]�o�ׅFd���'/���n)cR_Q�k1�aB@���RG��~Ld��{�iz�Fq��{{���۞�#�2����VM�o��d=���@W��Q���fU6���<���D�&�Ԋ`H�s<#K�[CL�5�4�ԋ����?5ba�����ɋ �xs">��kx�{v�"�Y��][��șz�����s
�w�w1bؠ�O��.��O���q�|����g=/qM6���,9>?.��z� ��y�m1���}r�F��ӱ��N�I6��ņ2i�Kv�Bm�B��L51xۑ�\aW�LK����ړmx���^�
��c��?�e��#��C;�:��m�Hͺ�9��_t�$U�`���ʗ��9�>�;��=�w#_q�c
*`�P����$���g�!��W5L��[�q�"�� ������!2��d4������H��%6}%�.,!o�ja���I����6��mK%<��"I؉�[y�����ؼ��@L���!��s��S���>��\��P5��V�W�Jz*���������)�}��-g���fe�m��3+�D��Dv;��ў7O��,�
	RI*����)$>��r��	l]���0���V�MRk|T�EY�k�P�Z8Kl����;�[B�I�(p��"&,Ẏюg.����ױ��0y7$�Hʃ#�y��'^�Pi�#�m����L)�-��	�N����ެ�p�+��]��P{O��_�]��\2�31dS<�lƋ���8��������h���2���";Q��^��X��r)g���~�V��]��~���j� J,��s'R�"�8X�­�>az��אKe�UB��N��s+j_�	���r*Y�����A���F�e�jl����/%����M;����u��7|e7�aȞj4�*�3��V0+Է���J	��[����TxM#K=���gJ�[!.|h�%�� ����,$����:����tP>�iD�U�F�`hd'z^��w.9ruD'b�����S��%���^ꆻ=��iԦ?��T�9�h�Y�e��#����{F����ܺ�7�,���\��Mj۱옲�k鳒	0p�����B�*��?��eHE�!P��SZ���"����//!��;��|g�,a�+�f� $��wI���.xk���2M'q��+;��TD*w2"��P��X_�Q~e����ۢ���+�~����85��I�=+An���;�A�G������"
�h�a�٢"Ⴎ?�y��K��iH!��L�u�?���y	�j˜�i��M/X�-��M �%--
��O����-)�]���l��ذ~�MS<d����M�rFH��(yI|7�]y��e��.��$!?z�D͞L�#)KXDm�<N���.�����G3x\�[�H�n�s� �ҥ7W��289�Py��ƃ�G�����#�����j�m��1�)W�3�h��[�D�7����65_VH�G������ެڒd���&�J��l��jG#OS��1�n�R
��/
�n0_ĉ�ҿb#�բض�T��� |��
8�í�L���v�QX�� *1�!ş2� ���Cu�k�(?| �O�p�HG���Oxg_"���p���g�Պv r���љ��V�|�y��t��J���3���{�Vsu�碄�$J#��w+��1}0ϼ���;��x������55 !Q�eLR�C�^˗�Է�j�+�Mo�	���$�����}�%"R�K�_!m5!��R���گ_a!��d��v���}��F��L4ȫG��_z1�)�lR��?�ZTF�[\W�of��$�.����5���"�$,���$q۪bW�۽#Hp.���:e UvJM���� ]��|4��c�')2}��*�P>�z�<�F{�2�x����y�߄^��eӚ^�⤺�厶�@=N��j���Y1���4��#Ng���SIK_��D��z/ّ�2_��R�8������RM$7�R�6�p�27��7���5��Tb���䑫r+��s���x���AJh�	*���Mv�������0�5�X���n�۵68��wb5FwRi�dg�G#x�wͯz�"�k�k�-��>�8���+z�3�����br3_נ֣���2�����62o���%84��������	����%������Wf���,	�8^OG�u�R�u��z�W"+�7A�bM�V��z[ɼ�	�Q�!�ކ� K./���;����QĢ��N�1���}+/�y[!�t�vӰ�?��ZY^�Ɏ ZW�#�-�m��a�X`�m�Rd�Ȯ�*�L)��W+^JOF�A�\ ��2��|��L���=P���6���!^�e�v�4G� *����G��8XIk�;I��J_��=����x�[�j-�F��[9#J���񉡮������qH>�6���E�ř�)�Z[|\]5y�5{�	x�'�'��]D/�<�E��ꏄ")/��(M��c���paFJBãH
k;�`��	�Č�	�M�ǒ*��	�	撾���W �pH�2	c7��c�gٝ�
���
�R�|�<���"-����}�`��MVK޲�*�^�y���"y�g�/�q_$�{k��E3�đ�I=�y���4w��i����� 6 ̈��ؓW�t�o(F睋X�����be*Z�ʮ�I��m�{'zy�o ���������{�}��3�ӗ���N�a�*ԙt!�� 	��{�M�jd��ut?Q��"z��g����N��MM������4K���	d��U��$��� ���N~�A���(;	g~a2j��De����x�rQc6)?聛���#���:�e�cd�ݤ���Y��Ӏ��ێ:<��e49ע����ݪ�TG�&����i���I��� �G*�?��Z�5�o @� lS)C/�:�H�$;�1�_I~K��ܹɘl; d@��>���Z�:-����4�i9�32xo�-s
Y�*�!����Vv����\`\Ȯ�<֙�&��_N��`���ef_�1���?�Z3)���6{|��vL�Pt���0�F�I3��c�A�e��k�͠�"�V�WR��=��q��j�}�/�V�_��z�����r(��e~�e5f�#t�sl����'�F�~��� (׎�y�.�	��]���nAꗦ�g¢��
 3̟��'��/#!d�d�~w9�.)=���$A����������$py�Hۛ�=��g?	-�kl�%�]��n4,�"~
�'tv���f�D��=t5v�n�`�n1����R�^��)�q�<�ӆ�@S�L&������%���?ϟe�k��?��Ъ�;��7=��`U��a����Z�v��܅U"������w&����*O~v�L��
�2@[a�hsGt��������'�F������@Y��'D�	��O�'���?T��|!��v�1��Zs��.�_��(�|^N�3@&�8Yb������5��6��D�5�������1��S�"X�R�2(���/Ł�@υ,�zǧ�[A����9�WW�*p�Ѵ��1*���aS���y�J�L���Q�}=�Ѕ$8�����i�Z��Ѣ�o�g�3�{�q��QSv|�����fDh!���n�8��'jb�3 	O�\�=��-\a3��1�h����F��KH�ڽ����Aj�r,�T)����q^�V�Fˈ����t��;�h��G�%�cD	
�9��b`��8�������0(��9'd�KS-��q�'�*��5�\��,,EF�������}y&I���Z4���ϑ.!��Չ��7�3��k���i������p���&�H��L,qk�FU���˲�s���ѥT����Y���Q��WN%.M�8x8�t����00���/�zG����L�"*׋iD>�U�1m�0��^!9��1�D[!��Z+hݫ�"�)G���Y�ĭ.T�&	%���ѐ�/�V��%��m'#.^N$�_˯� ��f��;@KK~���-ѲA��,��}����@
�ž�v���)��'��b<��.y�J� B��ډ^3#Z���x̘��6y�[炄~h-mа���&�B�"����)�y�`t#{^����/wp�Jx�Q�ʙ7h���#���`#7�P<�t�aFX���_������rs�,Η���t��@A�2��e���U��1U/6�����tZW��W^��D��s �[�HίË́���BF��Ÿ�ѝ���k5���ĔE^@��L�F}`�:�t�سs?#��?T�HÝ��i.BT�9��Y�L��~�J"<c����M0[��Ndsb����[�]!@Y��J��k��OEU�R8��3��k�f������;,�m����c������g�n9��> ������ރ�<�ҽ�H��9}C����j��)��d��QtH���vG�ʲ�n�B�L	:}<V�MP|'1%݆"1I�XX��D���`hͺ8WM/�ǥ�$
����^�^�8��A�+�{T����AF��	9߃�	�2UK��A���:�r��w	���o�N4L��P��9�xt5�'	y{k,ц��;�4V���*v��a��WC2ύ�f��_e�P��+�#��q�~.�]�r��z2��S|l���O�>(��1���»���і+7��Ӝo�E  z�zņ:��\.����R�`O�P�m����Nhp%?L/�z��2�b�p�3�/�9S�,P����#�K��e�6n�ԍ��7\���S��A��|g��S�̄��,��Zx �c^\9�	�dL�j3������������:��&\`�e:��Ha��
��*Z)�ܚ� :[�����
nO�V�7�Q�ӽ��P5�K�{|���Y��䭍vmWX'�l��p�Q���P�vl�}��k;$��ɜ!yl��B�*0$/]�_���L�N���H)�ubRI�h���|�mV�v�i�DE�}�y��B����͠�%�n������.ĝ�e���T�������p����F�N)dYL0ܮ�Q)�qK�J�ފ3WSR����o;0�Sۆ�sQ���"�f��zi�����/�QF�����������m�[3"|u�Ƹ+M�@�2|+�CO*_�&���z���R��c�`f"n"�L��*�� �p��؍�҈�J/ăP2w1}T��,�/����ۏw)���@fW�����<���WN�7lP�m� ����i`��s�r�*6n�V�1b�E^�0-<����_���3\�k�YI�XBw�n�+�;eh���tM�1�$cv�OK$C���z�?��-yj7�t�9��R��0(�/���8���A�NT��w�@�0�œ��~�� ��躺y*��B���p�[�$0%�e�V����כ�7�Tk��I���˰{�:(�Ϗ
�Γ��G
��t�L��.�:jkW�9��A%%�fֶW��q�~�j�"��;�>.t�������(���K:��[z������듿�K>����c8���f_��qɻ~�e�7���s��YS�̑tcJq`\_qH? �a�T��j#��N@mK ��Uu�5e�P��=_4./�j]�3��a���d�֊ԇ(�H��� y��S���S��/�g��M@_�-�}&����T~7���(������*��DHb@��$��F��CE�y�Av�T��}� ,������Pn̳��$SV>8.	�7Itp6&6��˦�#_ E!j�Ȁ�aT��[��Eg7���|�7Sp6
Mf��g�h�q� ���Y'�����F����'��.�`� ���(ʺa��'��/P���Y��25F	X憓�ћu4q�9n[ƕ@��~��A���M�o
W�d{��lH����%uq^��� �P����� ˱9�H��X��ۍ��o�1����;	0��j��^
S{H�<�$Y��%z�jڒ�t���У�mޠ��m��hp�x!A�HY��u$vhvVgBv���hw�$[eb��,[�,,;2A4��C�v�h�]}9
+i�D9Lr9������d �b�*n#js'0��wb��_R�[�]��խ�[~�ai��հ��i˅8p\N�D��F�7	+���o��T/�Lw�$�E<��U>L6^^��ɢ/�z�WTV���J��`{�����d�#�Q��99!�5��7�B�(1���u�@�mB��5���Ԫ�Բ\#��t��ӕ87�Z�	JWK/�f�L?�e	~c�4�1	tUn��x|�P)a�齌��U�=��I�~�d� ��]� x��o��d�v��
�@�
����Dr �v<�Łb:�l #�v+�t����PI
��̈����Pr�{-�qx�k,Qk7�)rs�i2�E�{̦��ϙ�>��vlO	j	�K��v�H*�y?s� ����b|�C�����{Z���%�E�!�s��
x� ����^GvN���,~K`q]�1����w'p˥�f��ɱ}��T]����î��w�4Px��Ŏ�~���iZ�o�����z���'#�{��z$�3��o.���}y��)�g�}W��zR~���ݻco�Wʃ_�3o$�������gEP^��K�xOX��^\�z�V)�B4�$�����!�=�Q7���Uu ���@�t&od�I�:��i����@�и��ii�C��BNV�&	�)����ֱ���g�E,@��i��O�*��W4������nB�NBT��Ƹ.�o�H$��ٶ.|���"�:�%�H���B��4o8ho`DJ�ܛ�F���L� @�����L�D��7�X4������ftx����������y�y)$\�8vKJڄ���Z�¼��Q�\�!&g�z�zY�x^���d�ZK��h�yd�RQ[��0g�.A"���,#��ۍ�M��ǩ9�!Z�x�$���:�B��Z7+�9�{�bOB.>���<�8__/MXs���
Y��T�-9�O+�1_�>���z����
���j<���3�tP��n�)���;:����P`�7���>ZΤ��*��0ovn��9�'���.�Ud��M��Wߠ5��3�{�{�qp���-�P�9��aӀ`���r����j��9����a\k�pB�9��/�\T��=}�0���`ʿF2�@��Tj�U�+���cO��]�w�|n/iim��vR�by �����;����>(�b��^W����Ŗ�ʦ{9�So��%�b ��n��^��������4[.�,*�͵l:xʶ���D�|�@�I�q�)��p� ��v��@;$㠁J���b�����Q�9�0I č�D$zE�1,͹ȢL{O}'�bo�uo��Z�q[��9=&�S4��6���Il�\�u�[U���O&�Lnw��jH��^ؽ
0�����i�8B`�u��\�^vS}p�4����(
��xr�%�BA�J	�L��:��Lv|�����Ȧf�V�%K&R��!XÜ6==63�48���z��H'wP���6rq�Y��G������})�L�7N��Om.	�s��<�d�A�U�~�j�4CN�����ˋk����|(6��a-}KG�Uh�;{��Y>Z�N�EN�SU�~�1������^Bd]@E*�J N�D� �C��$'Pn/�ս��W3}����8b�Y�#�+"~X��<���*|X5��TC��T��4=���BJ�j�u738t:.���uُ�q�u�V����QߜT����.�$�Q1$QV�}�?rd1[��Jp�G;-��C�Z׊�F��?-t|_I� AF�/���_j^�͔(JP���9{M���&�����.ty�ū@��?��@Al�����}e,ľu�`��Fq��c��ؓu���� Y��ji� zb�����d�̳�;�%oz.@L�B��܆��.�^&�H���_�l�������X���!�cGUyv�ߢ�g�S�j��(���ɘ�����²C�U�TVIy������>h�=��{5��%O���0,�MΥ��ތ��3-I9z�o�[�;�"�G�ݘ�	poP�iv�:8u��g���3�/��f#���y�b��e��go��V���謯�l;6���3yݤ�cL���6[m�ܿ�3  �GxTQ�M3���-ΡK�u
D���f1� Ķ�C�Mކ����@�����������FptG��2&���p���`K�ַ�wˈ/����P^8Tr���!�lv9�},c����m�آ�C
�

��<_1�"C�Q*h�`L(�_[�a���{�rg�?_
�)u��$~��~�;7C>?B&�+�/�z맳:7x�zdN/��[�uis`ŭ�,4=\����j�� ���_�n����
�$�����w�eL$��!�U�ɶjR��b��d����˙OC������h�`�͓�b����m�)�����g��qtd9̳� *�HF����	�ʺ	S��Xg^�I��ĸ!(�,�����&W���__	%�B��ף��� ߾[�X�'�
Qz�񠌐\�f�O|�w��aCR�0/��n`|�߾L}Cz/��5{��M�`K������Jl��qᰰa�՞���e݀B%㡉�Gs5�m?����T4%�T�[������Հ���t��Y� �˶V'���0��57NN�I<�]��e_��[�JsA�|�������H$�4� �4�}�� ձ�vi�L؂M�6Y���i����yBO6x����>T�OsYx
-A���8Be<���; ]��R7E�[�7݄3ѷ�x�4�ht���tю��ܜ��"s@W�u`$�վK�0�;�@��~tx�v�����������Feh��ym
*ĿG��I�K���M��\��c΁fg4�㊕g%��rĹZu�㢘|����� F&Ë�:��"��#� O�CuwW@�W*t`��a0�4(�'b�r��QZlh��skzF*�Vb�q�]ߦW��{f��dw��܄�^N�����x�#���4���`��#)��WSZ�Wbg���C���xx�H����==#�~�>��q���`���Z���I0/1eQ25we��.��^7Æ�w��/-�����dt)�X1�h�Tbه�im(��6#<l��E�.h�!�*�?Y�_$N'\I+����}�t�Y
�=�r���'�+$��?�P��bW�n>����E���]l3�9OJ�ah&u��C�J�/�.dRj��}�����\�IjW;���J�m[���2T �����Ʈ8�u:�>٬C5�}zB e'>�̷�U@��@F�;��鞋�q��ӕ-v���b�Y��A�V�F|C;�X��)^�~�S2Ŏ�P��j9��$�:��fM>
�B�e�����:=���[��판S��f�u�X��������]�Ha(�5ܦK@f� � ��~}c��S���f�Ȕ�
�+�軣D#�/GK;�#��	���2�ޙ-�8�1A*st*�K�r���ό2gF!���wf�I��rs>�;,�q����{ʁ����"s��p����af.�X�g �_��<O/#���ch�3͜5�O�Ylǒ?���ǹ9#��}��C���3 �2iI�b�ZOi&1iηA�%3q����x�n�1��'���W8�B �Z����z�5Vml�wn�7��G&�ܬR9����oN{6��bg~�{+ɑI�0ӣ�2�bܢ��
��}؛d����Ax�4)T0��3̄b�}ϴ�-"����J���Є���n�CW;.B#/�|`�N����G��C鈖��O�MMd�ͨ����vn�G&t�0X���V_*L��fOީu#��!M� T������i�RQy�����ߡ���ؤ׬:<��]��6��g���ܳ���]�����a�
�$8�(�ጐ?��-�<]��J=Q>ʿ�4�I�V�5T�	?~�̫��GA޼��KF��@	)-��'Fډo�P�",5S�b�jz� F���I�i��"����T�W�FG(٫���:����4gV1v�i�f�:���	.��ߕ`0������Q�� |��!jx���<w8�aT�����П��7>��~<��!�Z��cj"�FG����j���^5t��}C�n|`{!����ɐ.����tTYʪ�nf����ː��]��Z��cZ�VH���"Qm�5]e7�����T�Ǎ�Y^�L��
����D:�q�O!G�T���1Q'G��%&p�f*�u!���>�Q3t�(�k�_N	��%X�*��.GBԿ�Q)��{&�������3�;f\ �a$%�QH:p��2�ʎ\�KN�Wи[����-��{�I�u��}����==y���ҷ#�%2��pc�~��o�Ӛ�~��?ʌw�����ɧ�I
 �"q�!���z�=_��H"v���D�q���u�G�����{���ȉ�D�bv��[C?��ѻܴ]X���D�Bv]�(���r���'�ft9��)Ő�5��FK����x��+&�I��6�[bŀ��y^o�0a���8�%��Eb�����ؑPw+"4,�����2'��5+�KX�\_<ƍ��+0b�0��Ȝe��:���P
���	��O�0�´��7�A�4qcCR1�JL[�m�0��.����:N.06J=��}d�,極��g��q�N�l�%�|z��(�U�h�����5˕BZ��޽�F\
����C����Ǥ�Z���i3�NfD��Ti�BғE��Y��j�j��
H	%!�
���u-p��&��_�
�(�G�p�2�G�s]�{��L7�
+_��q�%�dd?���K0�髎��Pir��,v����!&��r��������k�������Ꮱ�����A�EhO�!���7���N��^W�����(�7}�,�#�����;$�Z�^�7^��Ґc
D|���p�Lf����|��Wt���X�|�VRa�j�϶��g%vk�����+���7i"��TS쁽� O9ϔ	�����+K��ت�X�+��Q"��7oy�Vi;�l`�nY���d�n&���"̹(�������3/��6��!���߱$}���G����fo�C��b��r:�X_��>kKUc����\�G���^uN�
��P:^�������`�j��.$������D�QB�,	~C��g��z�V���[v��!Vܧ'n�������+�5���	qH*�������"�C���"z�~��N�0����S�.�4t%D�Ӏ�/�ڛf%��q�=�8��u�k?��2��A[ަ8��!��c�=۞HbK�F]�5�y�K)I&�
�z�&� g���`k��=!����(�3��36����b�Id/��Rl�ľ���N�����F����#�ر�$َ%T��)��m��rպ�{�@N�Rf�A��A�x����fJ
��X�{�Ĺi�?6�2�w'1Ox��f���!��`A[�*z�I�eQ�D�ѷf#�H���֏�@�G�g��"�xpq蒁�@|��SEVn_����.�<����ǒ�M�~���A�?e�
�U;S���_��i�j�T[�����D���X�DM|i"�x-��@B9�\JV��"	(�8�ǲy[�'�z=D�Yh}bg�I7Ӧ�]���ۻ3J�Ni�@
����{R_i��F~e������vs�PH�N�Mal����AGg�׸��!�\]�NCo�}�)���l�Q=����$.m����/'wH?H^�Z����q��1e
��s�t�]�f�<��uv�5Ѫf�&�D���{>��[����� 9��Ō��&��~wgd�?`ĐB2�Q��%P_�T��j���f��/62R��-��!c��H�!�����pYƶ��QR��q������W�<0E��ʀ=�U�,�^l��6&jB%Mm{soP�Ķpo2�}��e+�:��09k����:,l�	���:�)��r������W|:��TI��� ���tm�3Z"�;Gt����?����K4
�Y
�Vd>� �㐨�)@!aj.��CQ���բ!���'�X�:j�JQ�N�<A5�`�{?�<=o�=S�j+��c�yj~x�A���^I.���lp�QK<�E�.Xc��AL�ȉG���(�֒d5V�b�t���U�H�b(>L*I,�*K�9�D�^��+��;c	ѭ�n�e�&=�3�N���6��2����Sc�2��z����T��8I��X:	=�����	��'B�Ĕ{���v��蓛���\��`4�+4=W��ɱ��]^������� U��!����GаXNo��N�8u���L�����Jk�*�e�D�A�6CWS7˪mg�U��\�{T��U쮸��p�Gj���:�K��<g{��e���Wb��C_�E��Z0�� �}�B�(�5��QN%�K���g�K��d ��8>��+�8��Vx���G����G�ʳ���{�N<������Ӧ���,�N$3η��!	v�j$����{/����pʧ�X����.CaH��T�X��b3Q��#V3%�\"�q�������X�ɹ�U��	����m�8��CK�j3�#�������Ŕ�+����M'8�����,��f;d7�[~A�Ҁҝ������
m�W)���l����^5َ5+Bo��+c�6�A���AF0�p� �/��QRR��ǖ�3"�����V/d˩�]j�>s*�Sve1Xޙ]k9�"�bg%�5�ΖioߴAJy�/�Ԫ��*���
�U����W�A"�J� �q7��+f9�s���u�3�]ׯ��iU�n��E/,H��a�N��z�e��<jkc���4�H1p?j[�n�W�"1`�����'8i\ԱD��a�@ȞCb��גXXώ�VÄ����������F�����c9�G�.A	�:<9����!����&�i`g��V,g`%�o��B&���<��`�6�{��s��r����q؆��̵nP�e=�*�����~f�,"��D+^8�䝵�;��h�)@@)L<����,�t~�Ɲ��M�&2�C_�^�tC����t�Jfn�Kgf�˅�ut��<��U*���K{#�W�hTml��/eh���5��ѝ�B`2Ŧ��ו!c+L�������H�yj-J��tKg&��O���QFv|�R���j�w'���F0��J�2$�PJ�S4���Ⱦ9R�h�2���J梄)wOm��Wq�y�!b�<M�7B���Ǭr6�:�R�T�Ԗ�ÛuE�d���!��.c���9�Ô�-�� ,��T��B �Cֈ�>Y��c6,:�GO���e����$!!�/����"��D��3����u��O��M|�;<4y�C����Ԝ7�3'�5Lw����b�ZRHۛ�T�\��X!_�D�d�U
�^i���ާ����T�]nl�k�#�$m
B
�aD��������_�V6Oet�N�* ';��ǵ8�� �Ʊ���e��3���o�� �o�s�S�W��g�[��^���g�!�F�7��O���G�f�WQx4�!b���S؋��ʬ߶�N��~��tEZ��9��?6��g��C��Cv�|�T/s�@�?0w��>�h�1���C�g�BH���׌����ZIw�d�a��l�bp�W�5 :@{C�]��>=4��d2��ƴ���0/r^kRR�V�,��X����F���
��=���R0�U��	��XTWO[�gM�ˋ���,@W�@���7��Ӵ(��{��c�_G�&O��jٽ���!5z=Yc��6�g��R����޻�H�@��Py`���ͳ�@y]����7�vV�E���X�w�QaÏ:o4xE&!�
XD��o�pS(>��D��3E�Q�N	�����@h��|m����@�����P�}��'����,<�s��m�"Du��d���,%���J��٫T��K�����o�a�x��t�ο%[H��_�}��C�#�;�����\�*^�#E�����6
/ʂ~�F����$�
��GXqR�t�e��(��¡u�>+K� �a0c�h8��wE&s�X�1�-)��U���Vލ�	o~og�:�ɯ�{��79�Np#����?�sPr���D�N���-�%6��7Y9��߾.�C>Lb�����r*^�ݎ���;���Q��,j�K�g�>0�eD�P��o��g	&;�$.a��<l�W��l`2��f�o�5�["\@BCp�|�jI�X��^n%�?JH��;hTc9��5�E��(#8h�-�GnΉ�n��Yx;=RߠMo�����e����o@�bq��Z���6� ZT,�{�ڐe�t�nԺ���`�an����m�i���뵣�^w	2����qw�_[�~t?�hOD7~�.j�W�59G�a��?�K���>���
��)�_��{(L�^%#�^K�;Sa�#����5R!�b�8�<��	"�Bea#�Kt��������W53 {H�H�PA�À���U��0��f&m115o���70���"]c��e�.B9�P��R��&��%�Y��c�·֨Dg��K�g�BH�K�	��9�n�������2�e���f�Lvew���q¢�,Ai��?A�hj&%>�����O��:����l8����q+6�O��&.�v������9B��}�@O����k���mw�kO�u��@�F8��kF�ڐ^��	箺��3 C�N��y��=E0'Z;���?
K���K4O �F;�G�?��4�5��[7�o|e��) ����6���3��;�Yfz����"-q�l,.��8��1�$<����z�>j�d��v�:�ف(~�|Ξ�h���{K�W��2�{Z7��<8�0A'Sw�ps��*�����ĭ���$-k�}R�%��"g������rSDk�k���E�ۚ�4r4�Zs��7P
\B��O��ߚ��R>�12�2܋�B��[Ω@:]T`JN��;�~����LQP;�4�W=+ەg�rP�D��%���\�[F����5�ڞ�fҔZ�5�t/<�[+ǣ�c���V1�~�C���f2����T<.B��|�b���ɷ�>�utR��5�_�
��p�eh��n��;RHq��A�Y�+���p��O�2\g�_�#N���o�+���W���$��؏C��8��)gu$Jc��
O���K-�S��P{;�9L�2y�/rTq��WB�r�B�f IOA�m����k����UF��H:!�6��m�/�l��Σv�*�XGjo!�x޳�6KD��E���9�� �S���[���vL"��D<}��;2B*V%��T��aP�e;��Hh#\�`"�@���W���p	ީ��w65rX:�-W���7m�K�w{)%����Ҝ("�^̌�KY��j�_��m�������QNa��U�(�	�q�*�D^r�˦sh��84"?�p3��Ց��NHG�_$���JYܶ(㔁}����~~�d�Jp8.k���f��4����.B�nw��ݢ��M�iY�N^ǠY�#@z�:d)�|�X�pϐ�D_җ8��p�hU��lg����o��!�tN�.�y)��c�mN����Kz�c�]*Ԝ�W��lĪg R��xZ��ċ���(1N=/+�%�熴t&m���g�+J.Q�"�0����8�{�'Î_�2o)cϿ���}�3�1Z�K�7�xi� ��7"���sl��7��MzkF\�t���r`��0�EUj[UH�����W�-�5�ϣ�ʆ(z�ΖL�fA���<��1���f�8䏣G�z)�,O�[C��4�W3�r)s�֡a���qQ��	6$�d�f�g�Ы'�/�O���T�L׋���s�c4 P�j����1�s�A��ԣ�E�{Dl�\頪}�4�K����u�E� J&��7͵�0���y1��I�ר�~�<�<��7���3���g�f�R�Z�H�Ll[��r�ҕ�>�
!���қ�6��HtB�U��k������K���6K`5R@�$n�Do���
>�a3��>��D?d�꓾e�\,u���N�����Fu�&�l�XT9��J����C�gpc�C�(�)@�L2àc|��,��#s����qYm#Î�z5$f5q��I=�`ȻE��p��Mp��}�w�^�|%��3���5�Cۊ�����
�" q�_�ԯB�On�!��u�T�tk(�Vr(#N�PIz���wD��j^� &{R�#m��T{vn��4wץ��
���g��2� '�,����ԓ���W����5]1q)�8+eu��Q\��~�)�`� �'8�/�hԹ
��ܻ�����N'�RA�l��j�#/:�9�:eE$s��Z�YihM�.w�OO��yw��*y ^����Ƈ�Pݑ`ge�9��_��_���S�9�x��F4p<7+��.���o�<g�H<+�ؒ	R�h��0��s�I�����s\��8�Z�i򺀰�^A[&M���R��:��Y�lc�hDl�* ��R'%a6$[�W��񄥊ic)����8_Q�:��X��U�A=�c��"�H'�%g��%���7��ǍWL�f�b�׆�,|f �V>��RK����;����D��H�"b�`D���ڕb����H�z�t�8��vI�p�O��s%�-�@/���c����A9�Ń����ml�: غtR+"�R��lضO`v�ܨ<�&�V����~@��-�X�8�� 6|��{dԝ2�-�/���x΁7O6���VI��_�,s��v�5c"A�I�����������9Y�.���D��2%W�I�hS��M1���{�����x��F��}��8�ݘm���I6����޺���?�U�$�񓷻�6�ׯ}�r�%�p>9�z�ͪVg
���N�k���b��)�Yf�e���E�C�$\��?���q;9�qlqf�R5��՚1n+w��V��(C�bǴS�X�;K[;7Q*<�8�=&�ed������?yx#�K��*�d
��XA����is�ﵵ~,�iAM8:�5�,�90��7���G��3ր�M.LB�`��2�Q&�E�rT�ř�nӶ�y�ea:�V��Z�R���[KY�JZ��'i�5��~�~��=D!$����08k�an>Y	���/y�����W:׻�.��)tSL�՜L�6k)}ψ)Iz��g=��#�zCh�"/Z�Y���Z�{����?����
�/���\�L�`pޖC}E��\fv�m� �V$�d�&|�	B�!��~��)E���\:R�FU�(ڥ�>{ J��3W@�Ӏ�n�O�2�A(�~b��̄q/q�LC&��\��ΜJZ2i�Fn�c�d�g�1S/�(e>k��9��6vz{?��!a�����)ni����sX��>�'2]6�9��&!iP�0�ۏqp����7������2�r$
ɾ�l���o�veb�K��mu��L&��B�ȵ��ƆVۖAE_lv��Gjt~4-;aX�O���C,��������F3�J��$H'{�)��1�t�a�Z�l!�v-UlH?V���N?��
�^�������_�vqKz�SxE��v!o���̨���Xg�a�R�c+P��<�5+A�zF�Y�|�h6�o��>�HXM���fw���&o>�z��)�y9�j2�s�:�=���ʱ��&�uz�/��߅3F��K6�L�>T���?Z,U ^��4��Z����ܢ��U��� FJ�/iVd�@y�J�oH�PoD�'���.� ��6Oh5
r\��R6��q��{�<oGBlԳW�dSx�(�vI�(��)��%�U�D��l�;����4��m�d?�ke����ή����<�(����@j�J�9T���H| 8Cg�7��=92����˙���?y+�0ɐ �p-~��F�{�*N�M��
�%@������
���U4�_*['Ɏ�W��
7�~Ivgo��׳�0��T��04���`�>ި ��1L���Du%z���dx�Kd��h�EC�����a ���.mxom��ʹ}��C*��C�d�!����U�p��e�Q}��2&���͠��C itd�u"�b���7Ct�3`�+�$�ئ\Q��-\_�E���CZy�e`�d.�9����ۋ��C�O���^i7҄Nf&C���w��Xk��6�N�����z%z����c�/�0Y�-�V���b8���.n�C�I���ܭwM��iL����l���y��F[.8����Fv�O ݎt�qs��b���W�XN�6�gv�؝z��G��+t�̌�ar"7��+"�	����e>�ރ�q���
���K�����T�����`����d�4��2Z����6�p�'�Kyn(��>��6 ����>��� 6�Q/��%���l�z	VV�T��.�.��^]�(�RWE$F���e�B_�߽q��
R3P0�>�����Hvx��­�;=Q�J�%�etժ�î<�o��[��?�f4}Z?��uU�C��UM�Y���r3�9���J�^��8�_�Y�i�N��Um��ET��>�{B�9'�۩��:���N��|P��s~QVi��2�5͋���,>�_<\ȩ.>���䃷"�|l�i\���_��'M��ܤ0IH]�v �����@䥐1�Z&^���A�P�y�_�Sp
�����"J�C�b��s��9����6�~1Aa�Q�䁭X.��4&���L��֍��H���{z�xMt� t��\���m(�^�́����bŤ�H�]Myp5����#A��&���H@��$~E��%Π���)A-4��ծr�4K;�� >�z��I��LCz3�*��#ݚ|-XL�,J֋RO`�c��_ȀW��8�l��:G#�t����Y�}�Cl��R��ah����sl��~#��[�SCg���o�W~Wn�{ǂ����#9)���2X��wn��B�����ef����ؐ��6���]��g�y��L���b�v����oF��ԇj�kf_fڜF��E�Ǭ@C���B�Ȗ>��@m��7ζ�8�*���o9���M�פ�JP�2�W��R�8� 8e�J&$`v����.��=q�V����@)�<e\4��O�y�C2�G�e�	���ȼ�Uq�]!�U��=7B��47'�WאVa��ȣ(D����}G����,׆�r-��)i�������3c��2}�نP9 ��\�ٜƁy���x���.ꋎ7d�2�����	O�B��>��U��� ���fcT��o���ܸN0�ݱ�	�zZw�����I�ɷ��a��F"���%�]�Z�}`�?8d�/aIi��͞�&�����d�������m'i��r��m��-h��a̿��g�8 ����g�l1u�S4���;_�	`�$�|�A�`�0ȶ��\��E�@��e(��Q_�٬�e0�aN] �D79��`M�EFTN�����ʳ+�|���-W{�]�G�`WhV�R�ӦA/-[w�LPW���4m�^�!,3��ۮqZX��٥_�\9%�KK��������V���ϣ����RD���P�ҿ���UcK����۲γJ͟�f"�F��m�.�V�n���׍g|�����=���P=���
��_2X��B~=.������ѱ����^4B=iĉ��Z��xs�y$�����K,?���}����Y�[�XA�q'>�$-��4�����t;&�+��Dt˫���`yu�R�ҷc!��/�2Ut������nFKz���C�iY&������M��m�7-FʋH�N�y�V'E�Q�wU7b�e"�r���S]�vqn`�n�������d�ی\[np��6@L�Ya9����
NYtJ����u�rG2h;W7RbJ�S���^�g�	i^$�@��:�ȥ*��q�ᝆ��sL��.BZ-�L����Ń�q�M �
U�҃iۥ��/N�A}j>���s3�|�4�CǷ�����NSգ�f8V��I�B@���N�b�E��)�sP�?���P�h �-�R��`���x������	�Wļ����=�_��GV��l�'6�'�h)==�a��p�ۄXh^�W0h�g<�ߖ��/�߆#�u����j94�ڥ���0!���Yh���_��!��ʲ�H9��9����3YL�!��H�=�ԙ�Ze����z!����+|`ꀉ�?ǆ��%aށ�7m����I��C#��c�a�����F���r��"`��*��JS]�o��)V{�1x� }�7���a��c��澛�4��jʥ4C�p�����H�v#�^�~�Y�f�5�a'����~3�*i����Z� S��������<I�YYahؘp2*�F����9b�e����$l�R��ι��T6r��E�Q	+Q}3�b'OJ������5+1�ʢ�����Do�Ц�+TsF���W�b���䩰���M��X�2���b�(�z����&�+�=���Me0��� d�OW]�.��ET0`Kf����c��è$,B_v��U杻s\\N�a?��kAn�An�qD
͂�Ny�Y���E��SagJ�8 ��9Z�@)76����-���l��+���V�[v�9�����8�/�5�8��o�Ȭ(�zF��%�X��4���$J+f����B�����e�����.��"�����SL�#+����A���i��[�~�L�����(g��
�Y�O?'����J +ZN�:����4i� B��&ni�OC��8�?���vqI�i=��u%�eMo��6����K58f't`~/���3��~I�����
dɐ�q�7��v��3[چH�7��T�ţ�܃Su�o
 ��0;t@H��v.�,��@T��0�ʯM"ߔc���`Ú�Om�u��579�0Ŕ�Ѯ�l�.���7�e[Ob&R_��˹k�*`~I���l/�_�`�)FX�㷜tzC�D���8�J������̕�0�8�k}>��~{���`�(��H�k����dŢ�UTƀ�/t���,F3�r �(���F�J/�"'���ʿ��e���|�)�"�"�l:�7�ۗ�,hf�_��#?v_B#���랄�1ϓ�"�(<���T�����f)
��3mqY�J����4�~;�%3g��#.�yks�\N/�8��=�!S  ��.n4]�]�P=�z=�}��u�ۧBkL��)�M�����ь17Y(���]�i��Nh���ڄ<)��X�"���ɸ��2H��yQp!OFn��
��|j�H��@Ƈ]��ķ�e7�?���VB)9x��ע�c����� G	b�O�/�,o���� �����iNo�5ĕ���}�����S 9�P�uf�V����I݀��I��S��qQҒ�*A8��뾣���5�4�0��	�ɉFcI�NZ���� aw��B5ۘ�L�V����!�{ E��vvI����y�leS	������N?_�q���	{��7�A��x�e�V/�S�, hL�i��y
�����
ϊe�ͨ�у��c��ͩp�=� cD�}��{�MuL5s�|�������'�dK�|�5��šN���ePqk6��=y	�`ש��Zb'n�}.x3YL�d���#�X灆��厠l�d����\�<��j+����u**6�P�ͩ�~�!��	$lz΍K�a�%��&w���P��s�<����#�E8�X�'E}A���_�{ |V)��2^R�����OI|�J�$?U��Z�q��r�S�W4��M�0�����#�`h@`W�SϱI=^���#(q@e_?������S)�N��-��]]�����l�3�mz�:0o�I���'#R�-����[�6�w��H޽?�f8ƶ������䐋"�9Pa��l�$�˦�Y2�Md�yUu�-�6�]�o;�$�GF�e��D���ޟ�t6��&�+�ma����!%Fp-h����`=6/p;k��6�й$����d�P�o������?|�l>q�6/�H���<f��]a���]�x<�+$��"��bNd1�9h�9��g�$A����D{Am�z��i#��Y��*�,���,)/��
�Ӟ��6R�	!�(Oq�uL�	�M<H�,�.�ښ[@\��=�1���>`��B��G��a��wp�\��O:��3�-b��.>�>Y�`tY�!sn:��3�N=�<E��X���Q��(!�5;�揥����d�m	T*�C�-A����K�M���q��i@̉�]�n����5�I�C�8��+>�8�k.����l��Q��C� �5�*Z�B⑻x��zQk%��d�����a�ܡ��k$�G�ET?���|@iYȂ�]YV ��X(H�sOu�f#�ml��4s25H�R�9!���X_$�p,t�,��f�ˋ�j+����|���'�6��<Oa2�=��8���.e�R�	+{/3��a�t���C11
�շ���F�+pԃܻ[#��3sПw;0����<�w�{�\�_�.�a��lĲ�`�C��C@�
���rۥ��h��/��f��_��/�*�h���M,Dи���;Q4�j=���܌��&�f?N��-�u2U	����yS��P{��~��T���M��/�;����rg���F�YM�����%t,����xՠnB���(�p{��xJ�4��,��s�Ќ"�Sɀ��簠5BT���>B��
����.L���bDv�� ���Q@�� ��z��d��{��5�m)�ȟ�.�򻭡�@��	��+�
�8Oz�K�$���*j�S��	p�&�(�v��3� ^�)�YS[����	Ɛ�5�O��5f��!��Z����'�$'�ha|Mxz�0|�s�H�.�|�2S����Hb�ƚ���s�V��h�g?��i�6*�\*˻�)*�ل�m�S��Dh�Q�_v*�l"�֑���?,�	:��Y	y*��^����FYh�����џ��q�o뙾u=�.9�*�Z1�Bq1֔��q'�Y7�HCwL����i^��t���E+A�q�;.�{z�%�}���20)��h&�{���y���ω)�У*���/���>Me�f]�	I��s��BJ|r���{�Iф{q�R .WUR��1nc�Ra�Ό����9.I���eB��OJ��Ew 4g���ڵ3E?��O�ڼ�p�q����;���c��f ���W��9����3}K��Dw�X�4=w)���
g�ꊳh���� ���Lz��C�����R�Usu��J,mŷ��v�3��n�ή�y�fT�LQ���鞮���K�Ȍ�eUqO#���M���227�ρ@n"�Rȸoͪvb���l�C��6\������*)x��z�޴o���u��O�4`kv��*�H7�E]�+	��YYlYgCU�[�L����6g��Af���b�����x��v�'�dbC���0GA?�.W1��z#g�y��M�-�-y�"�����ɞ�u��`n�����o�	��,���6��l�Ow��!�~�`����/B�� �!���1���\� Џ���zw�S�÷�Z#k� nll��y���gP,���E ��u���~����Ȭ��$񽚟`���g�ỽ}'w�/����K!ev�A�,.����eﵬ[{�bV"�$�@��絓�%�(C�Α��0����^U��-�f���Ӧ?*�
[����ޚr�M��?��j��xc^9��6�
�}�q��8����z=t��O^=�J�ł�Ff?�Qk�c�1X����m�X4}�Fk�)6��*)�_	ǎU�5��`!�����yE�Q�F�3K�
�9}���.���q�ʀN��N"�8��J0N���^������	��Ȩ�����GQ� "1M�������=U�-И�|������w-ύӱԽ�ɧ��k}l�St2l���OT̫�,~�j&X:�P�S5���*��9��}1���I%m:�{������,KR���H�U�^u��,mΎ9=�_����	xN�vWG"���;h[N8X#w��cm$�E�Beg���֖���פ�|�D�-�)cb�?
��TE� �^D�ȫ>�x��~�Dqϭ2��q.���W�#����Y\/:Y�{�'�`��_� .L�f��?��f���j��l�[��7����e��m)K���||�2�;Hp��&"�E����\m���%�E9��t@53Ո��X�T�:G3L@���y�&�~��~�S�}�i�[��?�Y}m"R�8"ePn�1�3��Gy`R��g�*�-�L2^S*� x����/�^�<A�ՐfEȉ�Ú��,�9�����d_������s�k�j�~	+>��+:(�p�[��e��
�K �����`�Kd8S��Y�$��j���1:B1"#n6��-݈���=�Eڽ]���ٺ6rn��~yd����W�$M����*�9ت�G���߆R'U^�
�F��G��b����^�֎��6���@�lQO��WJ$_^Ħ��G��k�K<�;����\<����p1������;K��{������ޞ��$��K1X�mq^n����[d�	ʈ只�3K]&('�����z�b������V�BC���8S����Vӗ��k�ok�dֈ�%J�xj�H��A�F�8̍Qu��w�|��������$K��L~{�c�EO@i)���oq�;!9��[�x3Sw�8y.���ש�d�����-��V��5u���'m	�]�z��E��!4�݃|}�x�K{Q`��啛զ� v��ͯ��_9"�x�Jv<���°�79�c��ij ����?���U!��m�7�9;ٱE�ra4����6�������1�4�k�_�*���O��1'T�K\-g�`0ߞ�[�z�W���P�vI:u��n��%���cE�����R��S]�%"q��g��i���x�h)ơMmC���ba�jj16�!���o�l�dJ[�VlOS���Z�I�
�n[Iv$�_�HӮ�'h�nc�^4�-��\d��#���b{�:���������k�<�W)�=W*NB�.x9����S��YƋ�=���/���F���oiY�Si��W�3'��H܈_B�~XE[���W�
2ᲟC,i?�Oi�^����"	Ѓ��"5��1��u�ꧥRk�[�G�p��k�)��FWˬV1���1qN�k4����8V�t[��cT��ĥ���;d �z<���������>�F2�8���
}t�z��6��0e�:s����f{)���$�{^(|No��/�/m����i4���#5c<rHx��T���ϙr�����W�LCJ:;M�[�'H>�bA%��/2��CjվJ���{�����&A�>���a0؞K\yp�q���-�@>��D��a�p����sS=/��eRl�4<�#&C��`���c|�N1�o`�˩W�\�(���/|M�c-J��w�U/�P�
BQ����*`ju��i=_o�i������ 
��8H7-�H�s��B-ঀ����꿅v�G���Hf?Bɉ������HjNLՂ������D}��~�g=AC����+O ���F�;���
��L��p
�����=��ĵ���ȀKH̀243#� f-��w+�sI�~]M�X`�$r�)�g{q^���G�n[��{�Sa��Ta�s�柁0n��ה�p� ���4��y�@!h�Q Jcf�؂�ɳPu���~����T�IV������.���Nɖ���$��3��KF/�ڂݩ>㏭aO�XJ��QR�dcu�똗�J�=�'"i��U'ÊMM`R��>3Aޔ���]Ћa�g��t�A�U�&�[�\�֐B7�J��-i�e�,��_g٧���,���F�9��96@F�o\[䦱);�%��n  G��(p=}�f_١�	�S�ĩ��:Hm%�x��m	Hn\��#�,C��/j5%ww8r!��/�ˣ��h�twv��T.�Z)�ȟ
8u�)ܓq���ۑ�~v�fj/���y�j!.{���RD	��=�+ �L�6W<[K�vI:H2��/���?�܊h}w�^k쵸ߨ�H����m���d�5���Z>�ǋ�j����?�i��[9�s{�9F>��H�%)P��JW�Sμw��ÑG�W�"#�p���P��AwP<��/�[ŝ��[�Wz�C��d&��:NJ���;�jZ�g��!�b��(X:o�8@�3??����&�b1�Rm�b�ʤ*>��CJ}���?`ϑ���E�����S�,��fD�Ԟ��gnj�B��P@ދ��<R����eZf�Sn�`	K��75c�tq�;k1���S������'���dH)�m�#�#���?��X�;�D�X8�t6@9m���$�� m����^Tj��sAR.�$���E	���Ie�ʾGN�(� )��ֆ����oԧ�آ2�Z#Q�2�M-���:�Ų��h~���NVͺ��ՈpD]�z�@7C ȁ��3dIc�U�L���(��x���?w��z&�%掕:֣��K�e���a��:?@���$�g��du�X,I+�)��$-D@-}j�ڄ��M�^�dwxb��|�ޡ��#��JK,�z�!��πT ���4zY�{�<s�4Ȣx}���2�B's[�P8���zC�	����_D�,鹹q��Ct�*4[�(�.�r	�z486{ͅ��= ���ݘ{�d�o8�l�W��l_/1���q5���!�t�t��k��/M-n�Y�^��jraA_*�k�K�x�XG�?C�R,���C��9�^���P�.YJ��;z��<]@:�N'��]F�\<�iP�q#M/�dw~����)��>b��]`�4C��D0�^���G�u��ev�G
-��<-G�Kf2-�A\�*�,ezS��hv�b�r�|��(��lp�Q��#����@d�$|�4�k�z;����S�#�!7���̉�EwU�s�}�K ���U�M�Q�߼�T��q��7:�.��pC3R�B�O�Ѱ~��h����{-�#iH>��}�:�-L���\��u���}T|Oy�˶K�Dl��R���j��댂6]`����P��G G����jά���{Ș�x�Ѽ��щ�#fU�18�5.�?��ڙ'��T&Ӎ��H���Q�b��{౳,��)�F�C����=d]�}�n�W���}�<`k�rxH��0}���o����<?�`wf0���^��,�K�{���+���q�S���ejO�^���go��TR/S?�#�"�_�t��\t�kD����܅�l�I*G�Ê���^>ö�`~R.���Z�uK�O!�ZbӴ	-C�#���3�Cya��/J�g�):)ϒ#����Pg�);�E���/0��+5+�g`����k'Ǯւ,�{�_���#�}
�Oʥ����A�<e(�
0���� �m�����J�<�9�㙕�7��5s���A�ƻ���-���RX�B�Z�PCv�wwn�,��(�'�'���U�vv��3� Hr_�bBY��`�����$T(�\�L�jI��'A5Q��G�����e`h�V�Ndk(����1+��w��1)WB��1�jӀƝlX���m�_�]V_�N����3��w-.d��p�a�>���!t���I ��<~:Ê:����m����[`/���޳��E5e��aF6	&�X�i�k@N2�`b�%Nߤ<�OW�C�����������;��O�Vp6Zx�c�E20�r��W����}�߹����>QXP�Q=�.�Epz]{�w����3!|�q����fU5�5G|������up�c�J�%(l;4��%��p��}|-_����Py��̾�ٓ�9���Y�G��֐\f�5
e;��R�T6] �H 7D�O�+��7�IS��n�������Y�<7����	?	�g=��*9
ۜ�;�j��ݎ�6$~��4Z2��e�,}�T�&sa���*{�N2�il5j,�P)�м} D0�l`��T4���[^���P!�G�G�?���=�;���$+%Q<�P#?h���5�熒I�x�=��:<r���P���<et?��R�ti�m��=�ZF��{cE���'-���l7��K�BB~R����P�I,���	щ .m���S-�f��a����ʎ4�i/�`#4�H�l�����u���	U���i
�C��'zq{p��}kCZ�+x��l�.`��w���e�7��z��\����@ێ���H�!��&���I`�˲���0/��)�rldA�*�����c�ʳ���Q�Y=��+>��.� ��@�EJ9�xN
�a�ib;͍A�0ċ��>�NP����/zM���@�����Һ��o�v=u�ﯸZ��v�y��)�D|�W-�I�'�`g�=��H�(����`�������۞7�>��tVÍ��M�.[�	M�_�XـG;0g�AY�δ���UL��5+��_9 C��9B�"����)Xp�	R��B�D!���c��y6�S��剏<&����q�O��3`��j>�����|��cf�YΛ�މ���������^ז� ������H���]�U��m)��g�r�<�H�t�x-S+4a�T�ܶ�1��PGo@Z�M �j�#�|X���B���Sx]��J�$"�prS�u�KG٠���ܡ�n����M�GZ�@*tn+����k;z�O)����B�v��C>�a[>�-A���ү�(�N�)Y�������̮X��+D���KR�j�&�򏘻 �ܰ�bE�tJ�Eߘo�{��T�TȦ��T�'�1�����}g�m��<�C)̿I����J�<��ثۯ��3^��B��=s�E��*x+{��
H��>��.[Ŭ���S�O�hS~>��It����xM���|�<��'_������X�4�ފ�0������>ī���������S��{{0Ͽ��s3�}W�.j�4�d�Q�UY"URQ���ƀ� G:�^(Mv\E��>�pqd6]�h�@�����L$���?
�8�����&,�[��� �i�{0O�TXF�w9k�/{�t���=YI��`j��G�� ���FZHN��~�hȧZ��"
�n�f�����4�S����U5�S�ˠ��o���F/pϪ��Ĳ2:<�*�;=p+GM'qnY��"O���UK�o^l4>�,��O��z�Y���u�����8�o��WO�=G/C*��MIo�mժ�E���J������Txv� "ڛ|y��;��>�i�^�G+O]�c�@פx��ס��܂���ʿ��b��ej��|��wN�jd9�4f?;Z�036�!�lP�PF�Xf�{���-��t�D�)��.�;�h���+h����}?6K�3��z�J��_��j>O��u"�cn��(F��Aٶ�h���?H���T�门[.�픙[�9I�wI��)E�L`M
�_�a�OH�L�$,'���� N�R��N�Q����{�h�?�mfB�\9$���85�ѡsF�#�p��鼉�T�F��'���g˩ �i�Q?�q��alt��$��j�IӮ% A����l 1�ja �\�u�Y,O�����gG͚�$g*�j�p=>Ȳ�W<h�����R���z�c���{ ��4V��)x�
vYG�Il6	�`V2^����S:���5�%~N��Tf�]~&�;��K��?ت�)�'N p?R2��I��~�捙߱�<� ��g��k�6�������6bDI��\"G��PQ�L��WG��E���υ��'〉}���$��f�^���t/�8`T���k�a�M^HVQ[\v�ۖ��HU;���}��ML�)V��-7�Un�)�և��>�Qۡ���%%��ٞ:#Ȕ�A�|��د,�2�U̦�I��0��Z#ZH�<y?H]F{�-ב�wU�/�ٜ�O��þ|q�Tж΀o�2�x�k��M%�r�hM���H��+�3�]�e~9U����W�?�z���Z���08����t��HG
���
aٲ�.��ذɡR���c�j��.'���Nu���ֿ�rT�'c���
�OVi�}��T�i�-Z�r� c���,'�h�?��MKɂf���"��/� �fr���%�%���?��c:7�YR`( ڍ�hS�ԊSz1�⍮��J�Z5�ʻ����+�����^6��IX,�E0 �w�Zɴ��̨�Nc����hz�lMs�����ȤO�mD=�����4������/*`q�&A�γ)6�8M��ڊ'uVL���xM>��a��̓��?��d�1��)p.�Q�� ���<��J���r'%Ge�|�)\�j��|c�`M�[�b�}����Y+"�P��q^O;�?��gO��+qB�A�?�~>��(0e/�I����ކ����6c�T��sr��m��Ӟ]*v2�OKY$`�d�$���pUo�~K�ޙ�g�����>gCX�����-PO�~��A�F��]�٢LBf�`#"��$ol�,~GV]����,à�Z~z�)��<r�ʿΓo�'ËbХ ޟ�ģ-N��b%X�G��(�E�48$|��a�] ��EAB���],�;f
:�(i��2r�t�|�̚9����{��UjM�>���l��:,����+�����=�f��D�G�����Ln�)��n���N�|	����ג�e�ӏ���O���%z�C��3bb��e;Z0n;�tJ�w�Ǎ'�k��	�2��ȫÈ�'���KA�C��ކ�wێC��R]����V�\ڔ�]��ޖ�9ttH+��찔۶h%T���o�8;� �S���;������|��4	�����j1t9G�e����	�s'��`�H�FG�V��.�L�`��qY˰�FB�P����M�����L�A��%�XC�/F�t���*��8�-'�����v��&��QN�>=�]e1Y�o��4�����TT/��?�$�D臺Oj��մN���(:�ym ��e��a�wh9<�{�ʋ�9�3/��փ��昮V�m����prɶ�-?Om�B�Z��\)k
�����@��IN��`�mIqa�h{ɰ5+��#і��Dm6>2L��쵛�떇$ʕ�-|.��L��Tf9z�(K�!���/s��|q=��1�znu�M_ֵ��\��l5�Y���������R�I��8����QĵJ�y9�T�O�: ?���ޯG�`t�&,������ �[l�C|V�"tP/�xdS��A����-M�t�-!yReD�wY@j�w[hdދ�F�T�pEq�eg��/ j���W4�CϨ��Ϝ��k�ʹ}�����A��u�U���m�w�ңӾ�;`������KbbAD�%nኄ1� ̧"����jwA��J�i��+�������D5ҷ��f�Y}F�.�֜�}�Nm���3�l9����m����P�z7���$� �ʨC�����ndMթ���R\�n7%����AT�[��ʱR�;����(q���$��Y%N�pj������_m����	�c�<	C�.��%qt�q]�"�9�qb4~�岙ț��l� �.����
�v�,�a����Wx�Xԛ��6�.�`��A��sԒ�QU��:��]�6i�!Gy7+2Q��F��!������ �"��jD�J��hj9��ԧ�x��<;�Ogj�(I_�A����"	�Z�N��v�;�22[�,���Ȼ�� ��,���ا��Tr$^�<���t���c�[�X4Y�l�Ҽ/w��������ۢ<�FB-ZbZ�3�t71en��"%h�X?y��OW{U傘6TE�F$����BY�	C��)��_1�ݫY��3�r�Q�\hx�� �!u��|�W��,ǚ�dFЁM�|j^ҙ�|Eb��/o�ѿ5I��Q�l�G�6���=%X}�杛�4)�29	�́GT0^��9�Wũ�l��b8��<�K���J���\���\
����;`s���6��_}����Z�3��곻�?�t��5[���
�o̢��q�m����Q�Zv����p���_��d�%��l���I����mYW܉Q�v[�:�8�X2��QN?u�O�"?��Y֜J)����Q����'B����O����)"�Qo�Jt";�&?K�JŠ�8L�A/�'t�s�܀@4b�-�a�s谸\���vь0�#�R�4�b�D�8�q~DN'���d <����
e��>�vZ!g�����2�9g;@A� �&qy��X�a~�fY��0��b��7E�=_�C�j�U>���e{��HX��p!p���U����+���	ѱ=�_��˩��$?^^c�U��3F��kq$�{.���p�Цx�qC$��P9������&��N`�=�)��o�U��w	k���ȫMԮ4��&�R�!y���Z<��r�Ƞ�w5F�� ��u�;>�t�/�w�ނEv@Ksr�݈�����s��_�̈́��FL��&���b~� �=�8�Q�+�����|���JV�X�κV��96����E�e����g{�h>u[�/��@��ԫ�=]��S=L��F{y�k3�L���ے �t��v��+�=?!gWѸȏ�X�=�����x��� ra�p�Z��j��Qw�&͗�U �1!�c~io�p��/mÚlJF�M��VT��x�O;d��C2�\���̿�>�� Y��XpJ��̾�c�'-���b�����|Mc���ۍ�c�O���{l�'?�ۙֈ��΄W�3�I��Ӣ� yc	kr@D�I &%����R���pL���d����fg�mu4�܌��o1J�m���{~%��̓��,D�"D.��ꉑ
��TKi�!�kZ�y��z3懴w��Ov�Cs#o׆�p��JK�Q����}S�O�h͞蒲ύqz���{�qU5��/SW�F���0�¡�dEp��f��w�'����3�(���f	����v��!;�����J�Z-�9T��8_C!\�Ӭ��[h�%���)�d��i}RIg�?���I+��|2Yq420����n�d#��~#Ѿ�[��|C��o`T��S�Ӝ��Y��o��g6��jP�H��Ŋ�2%&i�\��G�j��Q[��ɜ��7���&޹����3��)P�up��#�f"�s۸�;��8-�d
s�Z��'�/g�9^����?ԧa��2���9֨�\+	A��V��U���0�=��׊[Z�����d�n2k`��l_BLB��Y�3��j�C�8o�l+�aW�<�(mkk��}ퟫ��
�����r��qr1���˳�+7�apR4
 �;!���d�y5Xq`��7Keʰ���t���d�O��P~�����rX	�n�|b�La�J�UV�/��~���p�XzW���<ɞ���w����I\��ž���\�3�`��)ӣ��G顭^&CP�.4���j
|�T�qC�����آ�ˮ�cG�ҙC�>)`vЪ�r��M���E���V��2�;�]̅�X"U�F#.7WWU�YQ�l!�%�!̕�z�*�"ݖ����CW<-�'�r�r�7s���t��`��4!m���(�Y&�/1�	���:Ώ����1�c�[�6	B:�a{X��!�p��^L
;{�?�'� � �vN�KljWULK`9$�v3�G������x�l~�w��[y�J���>'�B������բ�m�R� (��%d��I�~���8̰�.��-W�W�^�O�k�zѺ�0�JO#i�e�b���[x�!���@�X��2L��Z�f|]�5�:a�܌�(ycu�p#���2p�$����1�n-Οk��_|����;x����Y�m����_,�-"�S~�z�\5�R��r)�^��9`��MtƤ����(�_�ȅ�tA�~�K��׎�GpN��PCfu_��F�`�zd��ʮ����W��Q3	�t�h;�f��Vͩ�}a�1G��j�=(jDP����� �������ߎ����B�#=��w���ʈ���;�=�E^��<���Qw⸈L�y	��o�!E&��dt2T|N*�J�<4���}Ȳq'���$~��-B��к�&����-X���(�a\��T�)K@$�Lȏ7?E���Z��p�T�fZ؏�6=������;~��z97k/鞢γs�¤j�SGI��N�����&/���@���M^"y}}F��~�>��![2�}��[�� ��W��t��=�}7P�#��t��wDc��
�a*�K#�7�MB��Z�������"n���B��-�r��$.mw�.�Π�5�]�|��(��zk�45z��0��G���X�=+{�!CN��l����(Vlo@4x�"a����uVC���e��k`��@�J�0�[{��X�`XK�P'�����hS�:4����*�t�m��4�Fqe)O�8�݂6>D��9;M>ԶD�ڀ�	�OQg�l��r,%�
����:��d���X��p�;�h�ڿ�Rw�Af,�`�@sޣ��� >�򄛰��5W&:����;�щ�C��}0��1�ނ�~*��q��a����5D��0�(C�"�%���Ab�O������=�иCO:PŨ_%�6|Ө0x���Z���O	£	A�
�R� �w�O|�P5�L�C�_�G������U��V+4�9є��P�Y�^�X�<�K�^���E�4�ƐY��c@kY%��aGC�T�����s]G�Zx;mbp^�e�a� ��o%\a��ѡ��R,�.[Ls)#hp��;Q7�5;�r�}����~��k�D�g�q�3��
$W)[�M5�yŧ@����7l���bb�	U�#�t$Z�ı�)�@t`7�yz�|�+�Ԃ��rϨE0��/��ڋ׳OH�M�J{�ࣩ*����"'B�#Ra����c7!/7MT�"�$#��E����' �E�m�w(�#6*C	�l���Z����~̪I\���.4k% iTYGK��P_��	��4�b]�=,9Y�̘��f"|2s��&�\�-h�9Y��"�3�6��$�1O1ê�9Q���wԏ95��	�WG��?Ek+�X*8*s�-�1S��2�m8ZB��V��k-9R��I"�3�V�*il����g��7��o5s��P @e�^JL�t���̟8m��C?dd�ۡ�-;�M%{�݄�Z/�#�9.pPc��^n�.#��"��GQ�(֍�kMeX��LZ����m�d9���Ɓp�E��y��NB������ou%�&}]h�o����B(��Q���t��E��q~ �yԐ�7�&���3x���0��������+- Vo	|������ܯ�3t��q���/�����53��tz�\n��T.����4�a[ZO@�D���)X@e����
�i���c��*��!�4W�$aM�hzGe<� ���k,��>��	�"�[�虛2Ea��z��NmBi���)�il��$��ռqK�� ��^����8��@v2�mG )G���X*��S�Cn��W��X�iE#��8�9T 㸳�����HKN�u��$z����]<lu�P�V,ʜ��u�RI�,�]��`ܢ��T�������!Og���}4�����	bٛ�6��p�?zj<����|�g��;ϖ`�+a�޲l����a�ӰGg-¿J}�c�O1ɍ�w<��d���҆ե)�ĸI��W#=�ƱJ��&�O�9�\�Z���>I�Fi��ٌ�@sd���jAN����j.Tp��`+��z���������F!:jB�2�i��C(X�jI�ƕ���%2ө� ^�:�^��$X_bjm���-)W�+�ݖB�'�!.�{�����A)��7 ��e����m�Q�w.���G��@f��&�{��
;��z^�0�X�]�56�a�&�پw���>=z7;�[D;z�^S�
x�dGJ��x�)��h�0���
��R�R���UQ����w+S0�]�N��9�P�zTu��<Yi��è
[�U��ժ��_M@��"@Bo�>^�t�"��5�̂�_J��>Ka���r�86�TO�R�����*'����'�R��E��Ḧ́��STf�*�]&B�U�u�Tz�=��<
��w�Q ��pm&�Q�����Y���T)�o�mJ�|�.* V��%f� �_��}E������<�!���z�C(�;F��D{�=�\|�����$�bV�k�\��֌��fR%�~�EE_�������k���/h}���,N)��yC�)�s��=F,��"JRr�@�aho�D՞�Gû�y�������fy�����������m�:�;c�D�^Nk��]D����!���oSI�3����꺫��j�$;��S�+a�2*��ĩ�	������E��~�i?������Y�����~̏�y�:�3O�wdKKz����i�k����m�~��~����i��L�
��y���ۚ��q�K0}�j�y�3
�;�ɏ*m�1�q	ƴ�!>�Nf:��'湰ݻ�	�aW5�х��p��p�xij�\�n�L�tf(�1��L�7�ʒD��>ve�p4xX��5	[��7�;�ƕ%b?]��7J�^f�	��}�u�ɭ*,U\���i�����y|!B������E�Xg.�ڦ�
�#Ӆ�>�U��Dt���	B���e6�%}����� ���N�=A����`o����WzZg�� "�!��C�ı��7���D�1�4�:]�֑��Je�_�M0eL���X��ծ�@guO&��ܒG�j����e�f�׹�'~�7�xuJ�b3��.�[5�l�R&S�`���Y�U)�s����Gr8�ڜY�U\��^�H�.쭊������ ƣ\���Z��d&��*���Q��LX��X�
�V;�ޣ��y������ }8�?
 ��[�X�\+n�Gp c�+�"3�s�h���	�����^V��P�}r"*ԡ�K�tB�̍o�'�vDs��a�6�՚gށV��%k��K]�F��<�z��g�L�Ҹ=���ZS��j�j�� �/C��'���f�g����:�N���C��K~;�+��GO��T��$��ʀwW��8.�m��vO���&k�<о-G�U�ji��H���8� )�0*�c>�?ry�"7��yύ�8�ɕ�I(0�J�5�`v� 3�H4|��9ܬ���nA����؜ڝ���a�.J���#J�3q�Nt�Δ����.��j�����`�w��,b�����%@fN}Z��^t��~������'�?�ܪQ�N�A����A�{���^�D97�3-7s��q&�fGV%��Z��w��wF�DK��z�����ϳ�z(V��,-��38��՘����xt�d*�E���`n� c*��j�ydeN��de����[$�f�D���j�X�P�4��l�jP'{˻�8ΊI��M[B`H_��5q�$~�0������blBw@R���9��Hʋ��e��g�_��k���_����^�<Zz�x�n�x�y\䭓/13�2�X7��8�I �Ӊt��aI�����n��$\'��%�v��� ?le��&w��6��� �v</���=�Ƥ�wͺD�b�]J��Ov�t�D���M�o��@TBv�y8<�?p�W#���ʐ�XY��t����7���W�o��\���\���?���{H�=�`�@%/+�%��hJZH�Ż=>�O�u�re��*��w���T$��6�}K��\Jแ��!��m�J)�-��f�K�2�Տð�����e"�P;��1�$#.Q������ �&���fF�W0)�w���U�-㈌��m 8���(F:��y�d4J	��8�I=�(*|'Ƭ�ӟ:��L��L 7�M�8p�N2c룪�{�	��!���GG��l�X���nx6�G�N���FVm  z��!`jx^����������������GY�S�1O�F�7H��wJgvw�z���-�8ڦ�\mS|-�Ҙ>�*��č��K�٨�L�a2����M�E@� �\#�6�Ծ��B˦H�&}Յ�� T���Xk!����6��I�=�m��ca�^v5��3u���6�2�e��_�$襻���h�A�J��l�ј�6κ]푿��h��Zt�@���)���e4�LO�l�
Y�n2+��+��&�?h1x�C�CmJ���Ȧ
����<��G��*�����53�!���n�e:p^�˝�4[S$-��R�a�1"���kt�J�=�;�X�ڵ��
�6��|���?ho�&���φ'�PE�Xq�e�*uмG!%����'22;���,e����B�,W�@	�#Id�+}�K.��R�)��pv3=�7
÷�x=5�������H�uP_���w���#��g�>&/�����'��d2nou�W3�(����s�Uk�Y���%�S�~f���� ���h���Q���ukE�)��P�A�4g:L�oJ4�:��;��W��%s\ٜ���6)�H�b�
��/b.���
d��- �9�J&^��[ Π������(��A���G^����q�?�F�B,��}�ˇ|R?�:�q�	N*�ٽ�xq��$z�V�
���ԝ��:���^��x2��P7=���qS.���`����VFD�Յ�#׳˥������;��HΗ��(���S�<�7�O[�%���R_<[�}_�=�t���6�LӰ�'��	�H�ir�k
���H�4��;'���<�bl��$6��ĭ�d�q̣5n�8�J�`@�O��;J4�b�aSJ��bs���*��ӱg�q�;`�냠��^?��0��ZR��M�x9Xy��q�Z��� ��f��>�G��ᰅ�׈���a�t�gι˩���o���n��=Z*1�F���}��J���&��U}�ݲc�A$]}�h��@|_{+����4�J�m��m�;L�+�6�:-%Bj�ӡ&�4MAP)l�(�E�A�a��T���U
������S�X������%m���]oHzh���"ѽG�I�PQ��I}�r���'�/����l�z7!٢a��fM��_^w7z�p�v{�,TGϧ��;-9����$(�_������G<�c���Kt�>\i�v�,O��<u��}�wT�;�S1���Jm����Tt�=^�9R�Hkc
�a���+j��m͚���s�CB�У�n���y޽�;R��0��������G�5�k�����D�;z��hC�dJ�U�T�K7{��@i�{�O:P����hϚ��6�m4�'1���e��x��C�6il�C0EL���B�q���#���b�^k
�~���Zp��vbA�y?��٢�1S�61&p�����џNA��l;k�n�:�n(����ĵ='*�1�?��^VFU�\R���p�訌��D�ze� w���Ϝ��$[�W��X8��hv���7;J]q�YR:���5E�x�4mn����@O.d{�*�_�5ڑ2w�q-s��7��n����j^���o�ũ�=AI����8�kr�핃>�JA!_P�X<�����K��\�Xp��0d�	�T���I\��\ѻ�'�6���^>���K:������Ch*;h�ہZj!׷Ӓ�)3��5��*�I�M;)��xU�""@r�f⺥�5vb��S���1���]f�X.�v����jR�N##�"�}5_n�\�At���>�4��ͻu�+���e��XkQ[5M��8���?  � N+��b�_�]%Z@>��o���fZ��o�0��S2����I���t�c���F�bp�N���:��A���X��"�z����v��!v�������N�{�/³�m��FT]������:Bk̐��=t^-]��~?�$�S(������]�r��'�*�t�����5���j-��؇�ݏ���d�8�JՆ�{�<"ƅ�Q��'S���O֫#�%�D�n�L��ŽSr[�c�����:u��K��T���"R�a,�����^^Rzp��W��e)��8Q��&@���ۀ1o�
C�`��h�����3�O�u������+ړ
�91F"ήޭ�i�������-/^�S�;�s�Y��h������ p�׻�#�G��@��d9�.^H��N�*o2��庤���J�}������3fL�j��H,������J���G�ys
�f���n��������R�1���)�v#=�WZ���55�D�czڝNw�7�����u�����p���~U�/�o�-���=V������E���H�����ڽ8�G��كg�Q���g���B���(���~P-�n|��=�ڣ	��V��#��|�� U�h�Nĺ�dGCлl�Z2Ght9��o�c�Ꮪ��bV:��8[#��%Lrpx�Ei��X�V�,���p�o�$β�`��@��O~��u{*�)#�}R�n`Q��M�K��SO2��k�}6p�_�w�1���r��)!�;�6��9ʅ�#��G��#����>��n��Vv�ٯI�#�{���Ja�d(���v9k��C��8P�p��6��Ҵ���r�Xğ����Zh���9��	�e��<0�t���l�ls�Ρ�H6ة&�#oj>҂��p3�O��smJ�6��bR�-,���l~\�=(�j�t#�:��X��Py�4��y���|H��*ԨR�NI�6��/�8
훨��)�
��I�t���
sKE�%�S�%"@&����Б��2ֱjY�%��}1I��&�)5'�<����&�@SF(�F�2��뗨)/0~l�9a�Y�{����W�)�ّ�و��*��$R84r�b�W��7���Y�R5�o���H#/V}�;AH��3�ÿ�P��K��L��"�!R��gѺN1rd��C�ĶyL��O��\��$�-[��81k�;IM��Ȁ_瞙��$����Z���v��׉�L�l����"���EX�cgY���,��b������`A�pG�#�fI��?T0���F�+,�А��o,��U^o0q՜KD"8��k*��s1j'�8r�Ǣ��,�QzС�->L�%�I#��2/�uonţ��Vp@t�XG�k�"j��#�����<�+�6�6�Vr�q�Q����N7X�"���=G�Tk��������V�����篾���x��d@M�ȁO�k��9��KE�<�ɼۆ9�.�~M�49�7�"�<���u�%)A+h���;������J��þI�8��ը�� -��4���8��~�:��
YFn�Wa���mK�t��<���=VI���D�����NY�P�s�o��,c��$з��8j��t>��e)�Jr�,���1ọ�}}K�Sfлg���ғ���TS�:st@� �k�>�	8�C�&��a�[�Wc���Q��f��4�*�J��3[Ra>�4�QA��%�	�L��謸v����u���i��7��(o���@\s�̣�d�kS-��GV������)�@�UBej�Sx�m��y�( �O����u��1$�ݒ��}�\uo�K��C-�+6��E�$bs�-|�f��|� 2$!'1zY��	%{ �;����x�u����_��x��X�M�n��:�.���͌-�� ���ŃR6�3hQ��h=�>)�Cd����G�l��;�$s��{���ܐ�hZ��g�F;��8�O��]��xnPt���j���v�r��0v�
�#����^���P�����%���.@ڀl�Tȯ�`(A��9����VE�!ڢ��#��Tz��1(l���V�밤	��P��֮F*���hU�]�jj���ub�(.L���)�VfYV�� O��F
nx�Mۮ�� �3����'M��&�Pᛞ�'�4���&�Kqj]�b����3.�E�{L݈�0o�s��5
T��癧=~�Z����*T��2gQv��
�uyġvb�eϡ���ꁐւ]Vq��=�;%<�Cq;����⻉���F��q�"Ԗlx�5~�S%��j l�k��`�2q�1�z��od���
���U�ȴ�A ?=��������.y]=���H�7tȣ'�ji�Q4i���<=`�N��77�߼>����J쥨�w�F� ��,-`%)�BU�?��=��}��ԗ^ci���7�6G�\o]���v����^�b)������@y�¤8��g�~��$V~k'愇z���ev�ꧾ�S�@8���œ���K���y�Ы���ø�p���4'����%�d�P�m<���� �*Z����=^��Ro�g{CŇִ{��㔃9������c��C~ԁ%wc�t^dj���y���j!��l�@+7W�:Պ7���t�f�$��9 15���i(L�~������A�r� _'	H֗���U%ah��O$�y��o�A0�;ܞ�<.�,$��U*�.U�q|�Щ�h$���P���UA~�j����GPY�4��9/���XJ!�B�U�PRb0[��\oxb�G�DP�Jue
�U&t��r�>`w$���i�"���Z�&=^�o���cF��=����B�W@��#�?L+���-��_��`�<�% �/�]��Ğ�r���'=SmR㰆
s̭����:�*�~Q=� �J����_�]�:{c�����:9�Z�5-��qxjmqd��G�
�kv\�gמ�Kz~�Y2��.ƙ"�_��H�ds�����1k��%�������n����G�SP�q���#Qr�2���,x/��!kA���cdk+���?*���Np��} ƀ��F:qWᩗε�L27����϶�P=b���,��:��.�R-O�1�y��.?�Dn�$��D��i�ؔ�Ӵ�ͻ�;п�٭$V᪗�u�o0j���vvj^�Y<���|5�C3�}W�;�We�|���T-´c��g]7D���M-B�J|����]�]DB�e�O�UۂQ�2�;�xmY�M��%�- �~��N%H�-)2u�������Q��ծ���������<u�Ёo�DM�'3��.�g�ֹ������Qǟ���JQ�HO��9�]���r��'�8�Қ��9�퓊�n� �a8�${��!���A	�*@q�S�T���Ն�ߗ�2ĺ[� گ:u�G�+�hA���y��mJ��xI�Q�s��>!U�)�œ��c�H��.�P6dK��°F��	�]�Ų��%;���9@~�SA�R�WPRQ�DS��٤���{���eD[��X�Br�Ćq�f��l�f��}��|}?%�^��8�E�~HK�v���S�Ʌ��N+�`2�d��rP�m?���F)D�SX�n�(�6�N���5�)5 r����-R�i�"4��͢FЊ|̫}qt��������+��C+ z����a�ǗΊ�(�� `���̋�2�Z�ep}s�FM��1ox$ņ�m��^������N�;��vU]�Q^6�9؟�vq�<�ߤ��PP��?~�1O�ur�*���x	�|x2L'["�%P|��K\\��.�-|���՟����lu$��Ui���a�W�KpL��)!A���La8aE�B�0I�so��铰I��G6��/s�ی"�ޟ�h�=g!�sl3����5u Ԭuky�3d��1���� ��T;�7���p��x0.Asܒ�v��[�fn�\�l=�J���.�˗� ���;A7.k�x��M�0�W�lV]T�O'~
�vͽ����/�;\b��O-w�rV�Y��4P.?����T�	r� �X���_�����$�G��f����Y���Ã���3u"@e����)hE�|D�᣺#�9��!*��X�H�s�3��ۀUE��g]���/�䦵������e��1m"o'���a���J;��G��7 ��:�Pd`����I��|��v�5p�a��p�Я
���u��i��I�P�H�]<:���n_>/����\Y00x�l>/�I��$Ċ���[��Cc�0%�q���z�gfb.m=_�L�R�kVo
�xs^�%,�&{{i"{j��6����_�{�Uu̚+z?�/;	�?;uX��F@��Iu �5~E-C������碀볬,sl埔�^_�x1���O�5��3�()tS���>I��j�w��$Ws���l��aq�n��I]|_]��Oqd�"���z��Ľ�RT���I�.؆%*q�9a߳m��@�l�C<s�/G��C��$"��r��o���-���h�DژMZ��t�͠����o���V�h����:�@c`۸�a2�(�D=ʡ�Ԓ.�&!�ᚰLS�ҰV�PN�칱Җ��u�%�'l���=Zf0@�PJ���̡�	�\Q@��*MsO�i�4v��K��q(�ȸ-�Y	��m@ɴ�R�*�#S����z#�Vm�=/��de�Fn~cu|�58o�NǠj�M��w*WeE�%��$�b��(�S�鋊�o��7����L2G�"�
�k��h���V�ՠ�gXf��e�G�Y�Ӄþc$����ܠ���HX��ٵiֆ���-����l!�f�Z����9_I�3�2��,��V�ͥn��6�HNsA�-������_V�#©}=jlvBy�i�v����S*�%[��&��\?���N��[vv�gp��m�(v���Жc{-���o��J�D��v͹�e�����'�
<�үt�l;�@�������m*U�y"���ye��H�]+P&�O%`�~��Cw����_��Hg���_q<�`2�I/)j���=d�����&�z�Pb��j���ȱp�D�V���a-�	\��c��фĮ������;"�H������mOP;����6a����t��k�T�cc�Jj�$�����a�hR���:��<��(G���������8YLw�m0ŏ������ K�j���O��=����ve�V8##���o`��#C���m�R�߸�@Q�h{�7��������V�|* ۬ ���=,ƘB@�����V˻�&Ɏ�a��zlJ�v����;�p��B3Ń�Ω������ܨ�
���%+�jD1�>��+��V�������݁�a$���1�}F��BΥR"�^�	�^p��D��-�/�3IZ�)vbz�$Iݓ!����zOTǋXMN���"�0,��-��v@,�M_K�c��t�Pa>��P��m:���<+�^~<K�}�`��r�J�ŭ��zsWF�С���S�Ċʘ��s|�1�v��9�ڼܕ0����gSL�L�#@Z,
ů��
��*�
�X���D@�㔛m6��p�6�WI|��4���ϑ�]CD#�a����͗����\��Oɭ�N�%�����fX���
 CIl#�n$�jf;�;&�h�k�	d2f��L��W@��/Y�_3!AV9��v��Y%D��?4����Y6�����w�F�6u�J����ś}�5�2ݏ/u7N+8���ԯn��w�/m����t�ų�QNLѷ���z��হ�Oq�æ�eN/ �jW0�"�=Po��#3�*7=����݋�Be�ދX���W��0�����Z���
Wz�	H��U;�aɩ'����z)S�y��fN�@û��B{��ǧo��K�?k��K��������i�;����H0�=��jܲ7�\h�^D��%s9����Wlwm͹�{�^Zu�qT����nmX�;L3��ߜ�9|��o���,J`5Y�8�həG�њt��?������t�^k�;L"�y��a]E���eT|�:I�0Ο�ѽJ�x ��2-��	 E kf�-{���,̷&g��9��ׯQΈ"�9,����AY ��w ִ����%�y�����R�����ZgWE�C3 �Y}��*R�_�"�s�\8)`d]1�(����A�]��Ⱦb��0p���(%�1�Pm9� �n�-z���;?w���g���[L#1ɣ!�輊f� ��3����DO�j.����x���޶ҏE=t:�����gY �Z�KVsP���.�z�J^���M���x��U�����>C��T+�E�:C��s�zj�,�U��	��4d��Y��R:F} ���"�i�8�Ds�m�L}�p�3�4ǟ%���׷�p�?a8�jz_��_���[u4-��.N9 ���G7�$�=�"0n�)C��b������ZA#�Fy�>��P���}���!���\a�� �[~�J��Y�.��K�|�3��y�����Pb�?����})y� d3�0^S���w���eQy�8������r������S`��Q��:�3貜�,b�1Uu֘�f�� �xl����?X�\��VW�nr�\us�+3V%������6a[؝��Z|�����/���oPL��鿋�BUO���s����-��t��H��hqʒ�����9!�M��e��H9cT�i�lC(��_�k���x��5���y��e��N��e���r�b��y�̨���Р��7P�<�C1\�̭Z�w�%X�)Xoa&���sw]2V�K�����A�/Z�/�E��[y�9T)��
����}�Z���d�ʼ�5��$�9������ۙ����mƥr	��Ef�_�1q1�IC�;�+�c��3��R�R|�)�s��MB{t �tMota�>/�b.�lz �
��	V��X�?g����19�"XD�����
�����Θ�U7�.�x���s�H�w�_���5��%G�Bw���j�;���XhK߭R�l��T*�{� �Z��Z���R˔������"y�x,Ea��7Y��[�_�'�p�<�����.ȉ��35m�&%�,��w?o2<�;<3*����"U81���t��ߥ|k�B�g�����F2�p�����>�uU�qW�8�GM�H�՗oD!=.Q�U�0��e� ��Э�uh��vDp)�W4�R�#��E|�oe�9*.V7����K�,��fV�5d_P��	"���1'){}�GI;�Z�2��|Z�������Ԭ�]���I���#�K�S�@�����iom�I$�6�?�-Bŵ,%�a$�ȿYڜǢܔ�ڃ�L\F� Դ{�9qK�?\7v�o�6��OqѺ_���C���H*�u�\�+s.������EQa.����د黚�,�*Ich ��tE%Im c�k� ���8���'h<{�`���)�s�l-��z���-�iS�'d��닦ꁧ�T�4�#�g7���ܢ^57]� �J���A���/�x(J�lL��P�D��HC:_jM���M^b��!/�H��_'!�}��q�mF�ORn+�S"�}�5�*Y4o�c
�k5呪�K;���w �1�X����["�'1��K�>ܟ튔풄��1�"��L����kٺ亮�D�XnMP;�>�2�yϼ(g�:i.��	�����7a;��[2�2��Z_M�~�>���q?O$�|0�xvo}b����&z����ESH,]�u��=�~�m��<���� ����~�9�G��EUT��ak0|����.ԊI����X�3j�9q¸$^T��u��ff�Ds��Lۭ���g�}����h���K���E���,�K�g�sN�uQl6����d5�֯�<٩�)\�ˑ0K�������p��bE Tg��[N>��nM��E]?�Y*e_ko��%D��Հ�Z`|��g_�:���q����`�p��v��
�����m�	�qK�f=��=��g�68�Sj��v�ck�R�V'0�jU�ؤ;7ۮ��o���cc��`JT�n$�Tft���d�@d�ՄK�6D�>�8�E
�{2��/��z�3���S]g��nS�޽��t7ė7��Q�fvh�X�݉�Z@����"���u|o�9 ^6C�a'�ps�5�t��C�O��(J�F?���ib�VPu��f�8�S���_��H�fF\0��y���e�F�2��~��R$ٮ�8�x\��US�wX�op�v^���8� Op?�|��p���)���-_g?Ϛ����Ǌm�;dw��=]��zuSp�=8F*��k�~	�7�r��ﹳ'�$�O��JAQ�dV�<�y�A��_��\�p	n4��M��	�4�γ�����:D~�cn�Z��H�Zk�\�LhӖW�b2�$�[͛;��v"�FoOgvZC��v�Igy�"wFZ�׌�.1o��n ]�3��4�1���K��ꅡ$2W��-`�����G"+=��0�vg��>Èmod����[�,A���!��#Q��}HcJ{5�wMv7ѳ@���Һ�|��yEx�鷢V,ѯZj��:cW�b�.V}7C���>7a�5$�ŗ�Z��c1!�H7��)�R�?��m�u�=�	sA%�C��!J�=�w�'uE8��x�O�b������$�E�����1�& ��`F ����{T���z1���D4�M(�o��x���$�A݉����6��/� ��­��%n4d6ٱn~"MӅ�Shz�7���I^�2fTU��g�9������@�ྶ�@]��¯{�_?aq��V��"Q%GI�ߞ7e�+!��eۧ�O:�g)�1�������R�7��U������-�����fo1��|�������,Ȃ��Н�s����E��ˀ(����]]|ͺ��]�������]���-�Ld�:�'���w�	0�H۪�IÙ���%_b��?�J!�g��X�{=�U����r铫Gn𻉂]���WM�}C����,*+�<����\�G��h3ٕ��|�`j��E�_��~��F�^њ��%#]eH�
X=C�n�?�~$�*,ā�RJ�Q��M땓#E󥙁��v�!mA��0���K����B�D�&�J����ջ'�ۙ�%�9����}iY%[JʄT�*�,$s�U]���̘�����h�����"�9�d��8�2�c�C����uo��:@n �!� f���z���٫��_i����r]i�Ne����bA8>I�Rߏ���t���O]����H�(�c=�c+Ȩ��� w`�ax�w/X�#f5%n��"�)u��&6�b{G�w�ʎMhAB�P�䀕� [���|�4�g�]��|�I_`I-�3$OT������I�z�4XQ��)w��g<DL�:!/�Cڔ�����.C�� �6��(9���Go}�#UB+!Hݴ��:��v��[d[�����ȳ�a噽��S;��}�h����?L�aԾ��[���]��uc7k�JC�8Q�dý�0���z���)��l�l�zU����E����Pk�,&E�`A5\��r��-����q��)(�@;͖��X�Ƚ��l��C�,OYcn�	��.9��(�И���ʇxl��nS+��UF�X�S��,��g�H��������{o���:��>�9�զ����4i@f��!ij�̔�h18S8���՝��7�(dh�$�`gH}.�F�gG��1ȱ�Z-��<��El�]�����uw��� v[.������K.0o����-%�I)����&D�}����Z��4P��ʮ2ȬT�a�{x���5cL����z�h�Ϳ�#������JH�#�:)��ܶ����O�M�!���6�t��mV�l��-z+��X[� An����� Ӓ����!D���>��B�&�/��oZ���l�wVQ}?��F��k(y��k�DԈ(_}!�.4xe#��z��q0<o��l���֩�ѹJ,��o'��o�'E���	������}Y��6�5��)�b�]�?��F�N�P|�9�Ԏ��jS�.	��8�(م�ÿzg�M�bk�U䞿�ې��{�]���l������d��M��Y�$����T_� 2fAd�3e@�J�c<�L⌯��2�Xmy�9I6ǻ����%g�}-[�AE(צ��b?������$W������ݟ��#<�LOt�>�����A&��t�!Ôm��ӳ��b��Lh��+��q�d���]F�
���s�YLr�+A��;��K��T{�Y1�����ק���P7�Hw1�|�Z,X����*<:D�� �d�P˙�,M�G֋�{�;��^���	e��,�`����z7ƪ%#�&��~����r��(�_�σ�E��O����w��%�c!rk�ԉ��j�ހ=�����/�.��Χ�ǔ��ѮF�L[�������D��l�`�ռK؞}���p���HOiN�&��0�� �Lju�lӶQ��%H ��R=�%��H��\\-s��q�5/��}\�J�
h�g]uSf����C�S�!	0�̳7��Xo8�g������,���_������!���87�������m�&��ӫ\��c�N9�o��MӇQSڇZ�8J���?,���;u��|��"��d�����h�=�ё��(BdM6����)X��C�ei��1E
{�/e�EK'#��.�s���YN���^բ��p�_�W�RO2 nk��o����+��n��?�K�o)�ƘT���R�̕� �+>T�Hr���uX�2�7���B�Q������&Z�w~D.#(> �8U��!�|=� ��O1���m��2�M�y��m'�#�ߎBC�t�d	ZD�/���D�H��w���hm�6�}�v|G���0[7��/��#W�bD�(X�����:Ge�W�_RZvq7��㖝����QMe/�Dx���w�~�cww'��P/K���2
���7S�PA�_(���-�IɠN��T�	�Om��1�K}TK��ݯ�z�m��V��E"��KH�g�8Z���%c2�B2nȎ��R�J�D���<���v�{8�`�2���fY�􀺰hg`��Q-Γ|�2�J�{����0\��ªדkg��ت<�g�"@F~x#_�4<�1{���/e9����j(`��1����|��鋉X����� P����@ПL�e� �·ɱϜ1p����عS����_ደ"l��q��ˈ���{hR��@/f��.��ʔi�֞ǟ����aD����Pd��Eg�;��e^��3R"v��� ]j�4�|9������	k��L+2K��Z:T�6џ�l(��8L0ݚX1sKQ�E�ǟ���������2�v�A�:�J�J��	Ƀ��(����eGR��(��BG��G�Դ��f�˹o�}ڄw���3(o\7c�`lr!�m�{mQ��0�N�	؇�P���� *t�N�`wX@��nc��K�)�O�&�[q�v0��'�7.�T۵������]�q�n���&h�V��d�U��	>O�9N��O<����u�����kӦ�.�z�~&�O%Fs�T(ڜ��h�j�	'I�ZT6���U��_TD�85����s���ϑ�<'���E�$�q���8MyK���>H,G3���ފ2̢0�j��IJ����6�2
:-�a��섯�������P�h��w',�^9FD-��z��~"��9�c��}}+"�:py[,4�߮ڱ���|#�K��������C�c�rV˱��E6}�����y�&�!�r"n��o�'T�jwZ>�b�p��ӭ��5����-(����ݺ`*�L4��B�0^M��F�}t,kfZ�^��KYv�t�SGH� ��Զ�sd�1���nE����s1�v�?!<ڕP�u�r�T� ��xJ�68U�B�M��T4�*� ��K���I��L"s��	ڙ�*yH$�q���/���EN�3	�~�_b"�c@^��8��S
>���LgQ��/��8��<%�d\ԛPJ�'2��Q���o�K���A�f#!]���^@HY�ӝB���X��Ͼ�h� �\�qW/ �(��,����F.C�hV��2�,'vZO����L=��鋸�  �4�B�Ss�J�8��)�PP+���	��&������1�흶��S�l�SB�?��!����B*Ѩ@���"o��;@��E#�sm�� ��u#�r���4�c���yX�-�S[���d�]h���M|��aTd8�2S'�名�m������D��y�$���%�&'y��sz����ײΫf�E��y��j���rCr��7�3C����w��e���L���CaU�&�,}�N�����s�u�(��Ņ@���'G:F��Jz	vn�ZpX��Tߓ��1�^�,y`#5� �U�)6�Gф��3�lG�o9?��^2��wm'��JGBnoP
T&��{���q�C�"Vz��ތ\�[�>/��Z������_��'K���ώ�Z�F���դL�ݺ�K��*�A^l������ ��=�m�ڪ"�Q�&/cQt���W~�����7l�eǲr�>�B^J �����"{�����/����Bn*`B������1�O����V��	��\��/�)̝��x�XI�'N�XZ�p���ٔ���M�y��0�W��|�\����ڽֹ+h�.�K�Z�QlhU��� ҆��1.A{W)|\J�����5>� ��^�<�l6��z�pVT���-Ȫ�S��� ��1扢z����Hs��ԩ[3�TռZ����2_P0m�Cr؍閦[�MV���;����5�wv���l[7�.1xH���u+���!��i��� ƭ��+��j��p���(�>�E7����1���Y�{E�_*��'a#|'���`
�7Z�K�L��i��ks�����z1���erԒ��(H2�,�@�t?ƌVG+	���|�G�uqP�G�����h}Y�1S<vk�`�*��]�p�&a��F����[����&흻������O/ey�i0_y<��,�o�K�0F�����g�@l�5�hMG�����zd�+�21�o�G	��)��88)��l(��y74�}����<�X;�?���ȃC]���-N!ӘF�x�(Kb<2v�W&��1X�m�6�"�b7)>Z���X���*���	B#����h��)F?� [���iǳjcw�J2_G�V�͚Xw؞���:�;.î�������;Ga�3�=ͳ���k�ѨA=b�(�j^ͳǋ��3Ҙ�����c
�j?Y�/�GZ�o�2�e�{�L��\��K?�S�?�`��D^��%L��l??��,nz�������������;2!8#ov�Ϻ�W3Ö�A���B ���߼�y��Sb����Y�B�9��)S x�2mV%m;8A�?�5�ٰkm��+HB�K�W�ُ]��(t	´�9��G�gh�$��:�U��{"O��YGp�n�6~>3п%��JН�.o�eyH4��4�W�%D��!��I���>
�v�?�!��F9Y}g�D��gk&Op!3��r U=m<ck6�-��#J��r�5kT�cSwu�V9؇�'wGI��E�bg�?e�!O�g���WBb�����ٹ���|�ѓ1�r�ф�h�7�+~�S�5��@�ۤd�q�o����ّ&y�=J��K��u�I����b�Vv��\���&�X�(X�������R P��#���܇z�_g�S��{�1��;������ӏ{k���w�o(h0���ޘ����<n	^����p�!]�[w��m ���3S}���ӣ��
�U���3Z�i/�-�w]�$�0�#A��pwP'���O��EJ$J���ء�8�����y���7��@�2�p�Ƃ�,b�By=��;<��rϧ�_�ǿ�k=aB^}؊ދ�1�5�7�m�V|R��K^q��8�O��K7����ЌW���+t�k�.���BUǹ
�A�t9e�� �[o�җt�h�_�Jk��:Z��B�r/N�c\�:���L_5.�� �d��~�Jit����#�5v��Pԣ{��'���t`�@[װ����n�:���q��h���� �Q��,M	�1���u�'�0J�:�����".X�)?��A:��Z�Z^:/�X-��KN3	��<�[;����s�"6�ʱQf��>�!�/%���
X�����waZ����g�C��}s��I��~�i����y}��7��z��߽�����J�2��a��=B��[��x8fg�g�h�ؐM/��.��^���b�>�k����ִ�d�>�j��A!�Ý�f��d2p���gò?&�V���2,c,_]���U�$5E�J��H�ҡ0-���q	"�wgv]o]"�:�w:hZ�96_��Fe��B�2��l�x?���U�gj�?��w���w���� �X����M��\e4ۙ}���?@VM7\b�������ˌ`�x<�U�XF8�͜& ���w멃�^;�5�
m ���!0+���&/u�:8�������)Ge��Tp����k"��F�A ��Eu7�бUF�[,��o1V�r'\�K�-�D`,]���3U��$Vtp��z�e�2#�,ݴ1���r,�{��{�+oǸ�+7;a���R�ҁZ籫  �J���<N�|�j]ff��A��=�9��7;c�ٞ�s	�ʾ��w���?�}�1�	С���;������y�?t��4���
Qa�bD/��ۇ8��/Sa��'2�m�H �^�+u����� fs�������/ZPE1U ��)ʣ��T��UT:d`N��<@cV9ǫ�&�2^X�ԙ�&+M*t�ٮ7�|����:n�D������Z$�J>��'5��o]���
D�E���A>�����Oe��V�*S�>��A}?MJ��p�A��L.�v ˂+EI��.�1��%���i�:�FJ�.#��p}vY�vll^�p�|��3憅D�����C9D@�0��U8�zWO����,�OY0t��.��ֵ��j���%�I�J�04#��mz�>�'_��g����[���f��AZ.��(�{],���*�܏LD�@Rz�9j���<tݻ�xh�,d�w�Y��G��B�	:V[��ihB�I�N��"��ɩS"�6�o����F
H=j͍NՍwO���dq�#U���Yd����S�֗�����$�.<�FO�L�^�7���5�%ք�(zڸ�?�ݝ	�mrֿ��<i���;��7�i2�h�-W��I!빈� 	�Ν�R��[}�1.�q0]~�<�����lS|awܙ�皱�>��P�|m���~$׾`x��WFjL�r��e�_{�N}�k�ON!�h�t(��Q�
�(pRt�Z�Ҟ�T�$:T�s��R {Yl��`�Q�B���0k�x"P��W�׬:�'�H�
� 5a��8�:i����N���j|U�=��?òbAR��~��f�F��e�M�A�����7�?WBl����R��ݘmW �G�żD�����C0,��ʢ��ϷZ��W�$�c��3���.F�5�K�ݥ� �����fݩ��� ( p֎� �Q=�����U!UU��h�BAk��DM���N9�{T
5z��N����wj�tϣ��n
��T<q+Ym-��8[�h�s�ӓy�$%�b×�W��%�"����=O��,K��>N����b�J!=�M�!�����M�S�g���c Km`�^�j'���}%�Bv	pY��~�w�]j�@�X=�9�?ł��b�o��uP��$ۦ�c������yH�.C�'u0:�q� 1�by���
�1�P��U�f)����Ӧh��[��U�R���u(��~M�@��ص��"�X�<ba�T�,���g'Ӿ��ʹ��<�_����X-���l��#��l%�+�jAe�n�_�|���@}����>���w!T��9���Ίb8�ߍ# pqs���Za���'%�(��Ń��)�����v�_z;Қɖ<�9ʴ-�U�av�Z��Ap�p���� b.0����E޸�@)�.nS�6�r�ed]�T���Q��9"^�� F+7T�8.ځgs���⢜ئ=�����;-���c��<��π�))sU��!gM��T�Gڗ����N$��{E��]v*Ȉf�DVͭ�\�Il��x	XSd[���@Uͼ�*�`cz]<��pP�wv��e�ٍ�!�]W��]��7�ݜ+HO�1�x�)�_s�#c�z-yM�L,a��ÿn �|��r��EXN��bD�Y�d"�h�(���B*�O#�FԨ�2D1��:��Y�q�z��A��ي&�C�YW�u�c���
�^~�G�_.�u_g��
w�k���E�셹`=�A@�\�%�F̿E>�Xb��Ж�/������U���<��9u��D��B�B��o��2��C&I���3I�h�L8�R�7As���WwIw2z�<TF�{��<��-2�<*�W��b\�N#���8,@�Q�䂙,���X�͋��ܪ��O�9Nl��R��_��x���cKɱ��Q|��eu�����Z#��^�SSE	R���>�q���	�W� �.sF=���0����q�r��H�JQ�|�7�dg�::��^�ES5�vP	��G��{���_VY��=�����ylV��zBP�0Ue��7���9(�D�˼�����'�揘Qz�qܙ@�W�?�G:���Y���H蓇[���7�k7C[��J����q�x����s0~xu�^� �EY��q�L�3���*d�@���E��07zp?[�=OD>���˓hA:�IҸ�	���#�tM�Xq���n�2�7B%)��-FAA����H�,��>E�7ߡ��En�s�\�ᑋ��� ���zH~�����F��p�üI��O�[�"��B,�~wr�3�6�$|t�Z&�ұ:Y	����d��@��L�����i������x���\��Y��D{a��ыm6���g@�`1��~k4�7/�&��rl[�ihUS�����P��erCjl����P�~�<��/%�̭��$O] �[c`3��*i2�	Vh8�!/�<m��ļ���Ӻ&�V�E�C����m��(s� �*,3�b!_�����q�v�	�7�c��#�QS}���Vm���~�F���+�;�ݸ�&�b� U�?��ɿ2�Pho>���u���ײ��K�p�����s�������k��\���O��E9>��8�(W��S �DP�r4J�@X�� �}��2rТx��G�)��4��:�r��s�{��6?�����PI�VGo�.I�*����UAT4��]�+��ڈ�yE�᪡)F�������:�w1<1��V-F�-r��>�9Qq��q���J�i�閨�[s]���]`0E��-m�Q���!��T~%�7�-E}<���E����f�\��<ϰ��j�4Ly��ǌ�ਪ�����Q̛�o�q'��ڹs�ב�.�o���SҸ����T�Y�|����C.YL��Љ4��.��XJ���bO���y0����;���_��o�C��r�m�;�I͂]�]Wsb0���PB�־�2�2�Ñ�#�צEA=�}z���s'����D�f�#��>�W����P)��s� �� �n���Y�4(K��@�cKwͶ�r�ύDJ�<��j��Pڑ�[ou5
G�Qg�8�̌·?󿼝�pD���&�G ��o�x<@�,6�KDq��}�*OGq�������%�"iU�yG\}����^g>�&$�.�K7Ƙ-�l�-�r�~ծ�� .�<U�$^;�D6�81z�c[�k�y�Y4��-�q��B}jE��8��9f�� ��<d���A���q,XoLR�?E���!���(���2��d�Q��\�6�i��j@�85��L�oK Qҭ�k�B"�^�_.tF?�;epp�L�D�Ʃw}�}9'_f$v�P�q��v	)��d[� V�����eSS���\��Iw�ź�H5��p���"##��Z(v�������/���k@��S/�6u4�#�p�L���o�����S��hMm�A�y!�btLwi��%�Y��ҡ�s)8þ�^���-C� �1����@��b�d^%x�>�)ֳ�d&���p:�6�O����R��;.���b�
�t����]�c����{�$�?!�S�����%����JST�D��YOLGϙ��m�uKg��O���h�1
�:��]���=HM�K����H^XSɉң-'(��锃M"㇇�����-2��,*MC�L��ފ�_����^H��J
��z�м<�·�?}L�1�ES� #iug�K��u����V�9�\'AF����5�%W%m�&�<�h�H����x'!�Yq�˯��SOI&4��gP�n<G���V��cL2ob�����-׫��wS�,FB#���� Y�Wvi[@�q�LjlJ;��e�8Y��j-�J<����;��!�qR5�b┲������-�_�4�bg�Ğ���4�_ۯ(�1�f�6��oQ2mq0���|��"c��U��3ŭ�����6��Cހ�.���eU��Jz��1C���/���B�?E�#�7��]2\lD+��mk�5P�j�(�,e�ӫ�+��3'~ɞ|�'3�b�����IXE,������+���
z�+�4�+��
8�5x{-g���1��0H�f̥����{�짰��V�)��!�i����D��A@�_쾄��X�H1�(_2����v����sm����ٜ����'���~�Lo}�Qp-�s�้T�䫙�6�Gkw/܏~c���Y�H��'
G]��H����U�OC$MkfȸLb�+���
	�AYD���X_�62�[���Җ/�?0E3.JtN��y�_A�qX���� ��[e��hj���>������2��5wcCŭ�)G�F������W��z�׋ץN�e*�&^ ��C����o�l@=9?���������
uOb�R���?O4�J�g�)��]�4�!H����@{�#���J2}KZw�W�-�H��E�3a4:Ô�a͖.����|�W£���.�ǎ�׵���S��*�f'x�͖IK�ˠ��>�&�I�����2gzo��Z��"�wV'�-m"�����`�d��}�F`�i�=ie¥G9&����dK=�*�@�v�A�rM��b�#,ٸ�̬Х��ý~m�oY銮${)?��.�R������i��c@d�Qj�N���$��m���$2��6��5Ֆ�4�e����`����#�;��/�� 	;i�A��lF�x�\
#��`���#�2�gj[��o^x�=�^��k����[��d+����W+r�������˥U1 Jk?s�x�$�t5�_�gl�4:1�M���1꟯F��;�<��%{净�':��h3:g*4|D��y����  ��S*���`�.�K�Wy�CI�;������h��f�W�YP��.S�G�V�|>
4�M`.%�T:��W��0�Of�x��.��s?���s�s;��]�#������|$4|�=?��P@�#=������@���:
�����_�v |%1��G��c,0({ߢI!�0�^J��CL���0sk�W����̅��B�f��h�ZKuf!�嘮h��VD�p�ǽ�IǤ��(��(E�$�
�-S�!�)�'+�ɒ����>H۪���('B5��]���]�-�!T�,�ĨV3����Y�mN��/#�JD��R�;���"��Ӄ���֟e����i�&�����E��')��v��=�Qu��_S{�Eg�4ė��@u^��;���x����c�w"��I��*����B\���dYIw�#Й���`�y���Kd�Y���"w�{��f(=so���0&�KʒsЩ�=��/���eF�e�Xg�
��P6J����#� ����M�>0?��.2���mr���x+���F���݅k~�Վ��Y!
��3]Z~�yd��y�,{%�Uwϩw�$�s������"�_qy��ݤ�Y%�LY�p3����c&���&����hi��u_!+����֧;Qe��G��s@P���;<������")��& 1����it��4�Z���I� ~��VT�,qeS�x&Պ��hL��&�{��$�X
?svV��� ��J�Qu�d���5�2�-<�⤓�^�p�ԛA�.�34F�T��v懂�ؕ� �4:��f�Wh�`��hG��Z%��"һ��A��vg/l:���V����k]OÅ�N@�[���y�� ���
 �Y��,��z&��,��N�&�����(֘���<Kzf��+�ZC8�Z�`t�
�x�`9� �y�����m��膎/�U��Aw1G��7;�@�Y	Wy��b�+��"����y{.\�Z��ܟ���S���Y6m���6$��Ђ�c�z
�E:�&#a��
&��C;v7l��]�C����#L3irz��?B.?<��Ϣ:�=)�N(�%74!�/����*;	��ye�YiF-{d����y�`�4���[3O�k���gq�;�x�i��\��x=g<pP��b�8�K��a���ָ�]��Z��!d���^��l'o5L��1����e��O7����>pl���t>�{v;l
�#(^�"Ɨ{Ǜ��������~����DHO�^�_��-o��m:�/��c/�7OZ�5l1S�&�y��p�vCgJ��D$����6SR����cn�N��Y<��O�WZ�J�1�Gc�g?2^�p�v���&r�J�z��8j�sG,�+0�����3�N���;
���W?�]T.dm�u�i.l�"�4��n���zGK��`z���n��ึ,bQ��y�|*I�|��5����y�4篅��(�c?���|�{��b١;��ڒ�p���W�H�hY\�����H�B�/=�Ӎ��t]��CӢg�X�����,}�:�Z�
�7�>��'���ȸ�zxeq6'v;�ƨ����q;���l6	�%��,-���i�!"��֯��&�c}�ȁ?,Jq3h�����T^�ѩ��M8H�Dla{��Dv��;K<�cp���qx�ƍO�E���a�&	|n1"EI���Ak �z�[�0Kס�����'�_�{�l<9����~�[t�@�<<3wxЉ2�r�x��o�ٹ�&�$j�q,�A`OP�q݁�6#:,N�U�������b0!�5�3����@�Ό_���N�N ��~�b�����D��I��#�}��]4��!dE�1��6���2��x�N��U����� �LL|�bɬ ��Ϊ��������~�%��RX$���K*�{%���	2�N�
�,�%r��A�k�
�7��ԯP���G��_�q�J9��7��]���IZ�h'"�^��ܜ�d��]#���%n�8|z��]�����~<��>�%�3�3��o&��#�U/�~H4���z��$�F�-`�.l��6e9Ͽ(C�.�Q
9�Y�=nI�p������Ӱp@9E�R[I9��i����ޣ���ᜅ�ȗ��yST�d����^`�A�.$��f�P��=�Ǳ:��L9̇��l��;��x�>'��*h5�A�E,�M���y�Vu�Z?G��.'Mnc��j-JqB���H������/�����ԚVVv�y8Bd�xM�{��:?�
�����h(X���dP)�|��v_�:�տW>����
Ӽ���gbÒ��Qˤ��.^~�`BM��k�EY4	�ۗϘ�><��w����2�3m�r>��X[�~�p���U�I/%�[� Y0�[a���^��ɵ�A�� �n�BFFB�������a=kz��x,YL�|�����*/+Ys~h��ʂ	*5-�N}�#��3�[�^�6J:^(���-D��Ș���O��]×;9do���� ���me~�b�s����@���G�bky�7�&9[���I��aV����YmC��{�=�y>C���Q�y��qS+�P���XW�W���u��ب��Fl-�a`t]{��Z*��YL��$My��l�������"�n�����n�����-6�$�s@�h(d�XW�E�)�J��.X���fy�p6�e~@��>�C�vSv�m�W�|[m�#Z�_���^\�!_�#2�^�u�`Z����],,M{( �G��:���?��ǲ9�4{'�!ʩ�A��V/L�og�%��	��V)�?�s�~e@I=�i����'���d�d��'E��x�92���d��1�T��g>u�U����`�_�e�҉%B�q�#�N;%r2uV�ᝒH�{2�:N�ބ_��<��3��dƒ�v&L�ǡ�.+���\}y�����eYx����]�ʊ&��~�of�~�$)r3Ƭ�� ��@�l��Qu{��w�����~"-��)�ẽ Mk��cWTf���ʩ��o<�T$�+��q��>�N3� *��U��T*��h�Z,E��С�3Q������sR.����l@�*�Lӑ���ĕ�8�@,�sNL0d��'��3B�h}�.N�n��}�fT��	@�b��l���;y��-w��π,JSǕ6�X��y�X�������R�l��䴉g԰H>2��w��r�Ű_yҋ�6��� ������
�6��C&��6����73����ID�|/�N�XW6#��&�.�t����ԟn/=�rAO��U�y鼱�VKFl�1H:%[V����O���;<G�#���D��C��g�o~K~�iX�Zf��U����L-ld�ohDYiwDʥn �	#�rv�~���ޓ+�2����i��|�� 
%'M���>�~^�lZ{;Eך��j���g��
���K-�&����C7�[&��D� \Ҭ���5,^7ǣVk�W
آC��8A��1x^���'�:�� �S�UXD�gBP<�P�i?���T1!����۹�>;w��տ>`;)";������wL���d�p�`}������B�mԞ{�h�W��4�R����g��02��,���h'����X6��@	D�S�8�l"�aOx���T��n|�p���w�=���ێiS���;���X*-1Z�'?N�ꮧ6��/Uz_�ү/�K<�/g}�f�a>�A��<��LE͌���~/O��/w�ho'��*��H��'��.��b�z���(�=����4��T�g��}��O5�BJ\��d��rr��}�9��"C��.i���U�|߾N���� 7��o}����5�����)��ֺɕ7z+�w���IX�;��x{u�'�jģ^C�/Y���T��t�a��C6��A*+��s�{"[2�ǘ��`��$ӳ<�bޱd|ĉ�cLj_���Z�prIh@�7�T3-D,D��o\̅�CI	����:-�m�h9'���"�|C��U���g�>��̠��^L֥V]�7�A!q�}�7D�{��,ȑ��[� k�M4����$"�	9���y!��?�T=���q坅[��}���gt���Ymv���/�sG�,�ͮ��!t�b9R��M��/�L#N�d]yΤ�����uR����A��C�U�SQ䉾z9��VA@�9	B���h����YYR��6B�Ø]�J�$�)<x2,���nu���R	!��M֌�"k,4T�6���[��N,�]�6�7�P��q��v��?`�$�̂w��(Q��;�<�N��V�����펓�v�	;T�t��:�x������6�R����!U�%������5�_��,`�~����x���5�S{�bzj�>���+�"���k�ʹ�A�?�G�v�*�TMM=�|�GǞ�C�������B�ZTiV���ܷ�zr��2��E��Tϑm_jdbX�ܕ�G[}�HA������]6�Jip��n�8��A�JO;ϚFPm	�"�ď
��f9�]-*��>���P��&��w-0�}�P�H�Y����R��r4W��:�9�h�o�-���	��"�LL
��z�����uDl��u��5ɗ&Kp���������[�_~����^��m}2ݝ�+�Z�i�s��Y�ύ�a|��g�{ݤPxEA����I�u8����f~&ü�.F�f�Y�L�G��pTc��q1�@Zr*m s޶v��!�d����#�c}Y"wǬbkg'�5,Q��p::}*��x�Y�%񻖩�����fF����^&%�/��
�e:93�_����Gf��("���ڱ,N,@���
�����o�(�P�B�K��k�Eڥ��p���D� }��x��^sm�V$��h`�w3䖜��k�����#.
?ܢ�f����-��gxD��nO`�ƚ��JH�D�CTԆ��P�^RS�����J���x�,���s��������)]^&�j�ex���íe�d��E��R�œQD^�-GT$������v�麐hFY��t�{�G'�7�#�^���~o��&�<L}�N�oa-ԯ�����(��/�p/ɠ� �G�y4��6�i�z��_:�δ�!s9�[��뽢P�+8�}z+g+�Җ5J��j��X��M�
F@I?%[��-}'��2�8`��>cA8��iS�O���l��N�Y��´i�<��� �7�ҙ�	�����)�"�r��=�����"O [Riq;3��D�B����n�=ߔjq�|+��0 �\N��'h3
��Kf�O��p`?3�Fl�?�l* 8���.�*��]���ΐ֨)�uhc�p�o�)ى����m!�}������ �w,"]Z��Q�	��vvARfg���"�t������ԟ?����?�I�+�^��VDz��(�kݛ5��@��@��~��b1��N�uw��Y@�*u�ޘ�>�sժ��,П�KR�-��T��l�tA���ː�H,�ST��Okh֓���DT�@ò�q�bWZ�E��sD�ڰ�n�?�����q���K��צ�Q>�ߙI�+̱���R�[�k�4�x���~n�|��z�l_��m��h��;i73��ֽ����`g@�ރ0lm¦HKF���{FQ"l�+f;��7::rXi�U ���`��{�����2������Zj�t��~�®V>�C������C@M���l�fZ��`Y�ƴ�"fsb|���R�N�6��A|`�:Am*�Un����oS�6�|�)܋�Gk ^ZF���<�z�lH��7���@�c�E�ӿ&�$)�<u(�)ߪ)��9^�	�E���n�y��'�
��#;v�L%�ͧ��OQ���[����V���"��{Ԉ?�YĤ��NL"��5�7՛�vȚl�P�K3�����B#v�[���|ɥ��p9�!���o�9N��;�=�&�ͽ��H����q�[���
ٵ�W��`�G������&uv93��'! �qF���k�f]��������x׀Θv��Ĵ�w�v]�\<����F����ȾNB�����w�A�~������7�Z�,�SP�囏�.@��d����E�r�v�ݨ�#{m��G���\��Nj����D�e��1�OSbFJDFx���r���Re���C~{�9HR�@��ycVŕr(���K��B;a��F�^Q����Odz�:�,��<@!	��.�͛��<�������(�JTi.�TAE&;����� ��,��nz���=:M�ؗ�|�������{ܝk����4�uV��2�˔��"�Gv��P�����i?`trS�#�?�عk���?&u�ӯWΤ�L���sy�n�e���}��Kc� �Τܞ��o'�S��y_)�^WN���X��b'��٫��;���ӽrFխ�R��DCL2��>iK���s���2�/ۈtʸd�����ޫA���VE�#o�\�@���/�G�Y�b+!���k�X(�|1Mrh�<m)+	�i��ɕ=|:����w6-��H��mZ=k-���cx��ꁭ��ɔ&�BQz��/��R�J�e>ցq�������aӏ�O�4�#����&�,��ɨ��1�����Kg��j�V��k�I'
d=� .��i&I�Rֱ9��K�U�S�
5���TZL� =4� �nF���+�����t�-��`OC�	�s�"*�80�4\��b�hm�8�
����=���W�Q`O�!�X7�H��omv���_��� �=�X�2&,�9���{�:|�X�أ���9Q	�Պ}��WYnme~��_E�!�7?ӌN�[Q�fq¶�s������ �@��2�E;=n�$A�o���u��鼁�݄.j]��8���+�=[P_�*dc Qd ��~����y�ݿO�^���u��qj�5e��Ntz�����ȵ��]�iCap||@�w~�u	�7a���x����>��7ߢ�Ă�.F1���0�֟G�����u���[�gC{S�V�#���(�D���A��XT=Γߤ�TKŠ��@����#|A��R7�D0����uN�t1������e��U(�~d�G���Dc�����O�>��dF�rUwB�b\_� v���~hZ�IHǅ���e\ 7t�+��N9#�A���ך,�x��������#��a\�=�t<����D��	�WB\�ήQ���=%�b��~U\n�9�Ͻ	r�j�ۙ(��D��~�'ǚPW}_�������-�T(��e����e4�>Հ��3$۶��L�qẃFΏ�Ax�H�Ac�M~r�S���xsPF��+�e(�e�ׂ&�{�q栟%v
�������x\أ�Ոa�����|2"�SC�+���LX��O?����V�CI��feJ9�[&�Y�f��|����q��eӪ�e��� H(�G�vw9�Ɍ�5�^Z䲨���q����j�ˆĵ�+0�2�w�bR㈇��Z���ǟ.�wD�O9��9� �o�D��໷��}�F��������[>��j$F=*���#ᇅ�������D��g�T'X'��I�#��ކĞ�˄���Xj�����(ڥ�v;�'���^_G'���-��uj4ZrSi�h��4�R �r]���n#�2pSS�w�
gL�G��ݾ� �j�F<����U�l�+� �$\������p����B��ϥ�AHw=�Xa��{��D��^XxZ���V�]	M�"���A�f
T���p�YM?Gg�'z%s�r����7:"�&�����5߽_P��k�&��	����a#�};:M�� T,R׸�����{j��y8M\�+1���JE=���&���G%����<��s]��!{�"\'�9����ݯ~���(8�6�Z�I6��/v}z+��V�$�"��C�*P�ϨjBs	��BF�T���γ�t��o�������1�ms�g����w�O=�Fx���7D�@�I�Vm����ҥSY:4ٳ�H���o0���E�W����H��$%���|�Ԝz{s��?���'{Q�t��q�Ff�F���ڕW=C�y��h�]6���z�w�P�����#�^wh�����ƮJ��3��#����8a��t�"N���r��G��7���|!f��#|�E��z3�����IFk(�nNr��'����Z��ܸ�ճ).����P��	�]]M�d���Py�|� ��Kd�z��P$�Zb�����tz+��OQE�:�-�C�"��m��)�5����2e�=���p��[D�rx��q��4�p2bu���y*3/+KJ̜�2���C\���=_��	r- �h������*��v��Q�D�Fс��vT�D���@?[|�@Ґ����1�"��A��od�?wT�Cve��/�U�ɫ���6��mL�C?Z�|@/d�ŵ�2)z�3m�p��=3f�7!e�5�ަq��@s
���s�6��*�צ(벥A�Jc��~�at�4Q�[���U�����n��=_��{����yd]�N�h�3�w0����"m=y������ŊJė;lel-��5�9B��
��&dX,0��ٰ�T�p��i�6g���NiJ'����Hc5�:+�)k�>�mN9n��������s����9J��U�������t���|��gY����X֜|�z�M!��G�����'vu��1/��o��m�F�]&��:��F�~<�Ê�ѕ�@����B��<f�Bū�t1���-�⸂��b�^�f:��$hy�g����H�>]�$y�'*�sx@���'.j�}U��A�"��K4~S�6���D���N0ߴñn��f+m�Y}݁�Ӎ@��?٭C�*,�Ӡ��4h�_�c��I�i_����A�Y���z@}�<@D��V���JҔ-�>����Y}�|n0;�QT�W,޼�d(���-�6���H�gϣK+7�O���$��_�K9���𬧷V�WE>�6��k�T	�Dbf���^�����?�.kW��cBo�_K!|ɹ��?��G�Wy^]�-��mM/)R���ء�cA��36w�ӵ�,�T˳�R'��{Q�c�	�	�ɓ﵇VH��?SE���D*X�#�_��y��A�.�dh���.+�#	���{�M���N��,����c�A8�*gJ���7x��#cZǚX�&�Ik��x_�L�����kԜ��}�i��x��]9��t���+�rPb|=�<F���|w�S�%�9U�����)��I���%0B�>�k��~�咢���xy��61<��[ݣ�:�V<���DN�w�,�~��������q��j�H_�z�l����o�3��>=����rB�H�����#�7SV)�������+��^0�An�|�@V�o��ՋY�͆�U63:g�����E1�л�ԝ���穀%�3	`�P.���	��GS�ŕ;V	�����7+{�q�.uz��w�U�{p�-���{��j^ؠ�?ޭ�]��)�u�0�����Z��55ˢ�t5W�dK�lp�/՘+v6���f���S�20��!fU96�!���&��j�j�9?\m�I?��[�i�.u�ѽ���|&<���D�
�878NǴVv"a���!]םH}��e1G1)��ۚܤ���ٶT<�)K!�Ĭ�h���xRE�e�s6���4�X���\i�����=�lVBX�7����|��K#�>��I�T�t̗��B�Zf�����'�0yyXnc" yA��Ӈ�n���W�:uLuub��TP��½�'_R4��Hn��v%�)P�[�*��_�/g��������5�FKdq���L�$�RȻ`!�
gf7��X�&��ٚh���#$�����������g3��G�E_�Y�j�m���+#ӝ�LJ0����/%�b���ut<ǅ z�1�q`����C(��g��-�_�����n����V�@*�8J;fc�m6�|�`�9�&o�(��?p��!wU�15p�EJ�/^��R[���I�
����������?�
;�6ig�������wz��ٕ� ��E����R�l�x���L P��"��폺���	����Vty����r0['���4c1NDx`^��
�δO
N��C�Dd��4JM��'.�pz��teo�F��=0��oߒ_p��$;��n�O�V?C�-�G,�Ȏ`���#�Ve\7:�1��IE�E#�|q.�\�����Q�Ԯ�Փ�]�����u�7�y�$B�p��qN`譹#������j��AD�1w����C������C�ɲ��e���d��2�ރd��t�"zWvJ��u�������.\�ea�g���@;}��� �N�p<|ebF�'�@&�G<��Z�
���7�\����|b�I��/Q�Γ(����3�a]6کU�(jY����MG�Mi��}<�'�T���s�e��ք69��G����}��o%i�q���ɡ�]��v�LX�h���o�5~��O}�����	p��Ό���l3�~:H�X�f*U>X��M���R�ul,�d7m��ATr��<i��f��%�\��d����[���7��<�����Y\
�},Q�b>4z��KGB�N��i��6ӂr��p��g���!�'�R0��{J�3�%Ӵ4��v��ٕ�eR� ^ec\�]ꥴ���$ƬI葍�y�7C�#�M톒(�<KNs��捸�� q��qu��`�X7�-��Z#��#���A�цR���Hf���U�&vǎ�Jff4������&�����F]��
�o�Ekn-��8���'פ�hz���A���.�_�N��;�<_T�$B��a��.Z��r��yi�IS`�1i����e���5���*W�(�?><)��M�x��^Ў����t�	U��B{�X��y�M6b��/�D�
����M����I~®h�6ෛ����V������X|nT��E��M%
6&l���J�����:J��U������Nu�uY6������П��*��wDJ�;�����U�������s/7X��a8O�̍���N���G��:�R��J�8�1iZڇ�
@/�����U� ��`t����^ve��^�K�T=���O�>�1Dq�8���؅��&���j�kax�]�<�(��m˖�vǆaz-�,36�� YY��q��.۬��Ѣ��"l�"$ ���&�@�;0���*EN�'0˸Ӏ�qΚShj�mh��_��<0���2y����b����_�-m��^��$z#Y���:[G�;W�/C���C���fX��B᝵`'*�H�U4���G�d	e�YX�'��i������y0�M�7d@*�ȱ�U* ͏2а�u��e���nJ_�/�	����x���L#sy�=�� Z�J.�XV�Q�5H�Ҙ6k�D���3��y�WH�C�?3
�Oݔ/��P����WP�|�������(⪦��
����I�@V�����Uv��:��m�MWH �.c��홞��jQ�3�[���>�!u޸(U*��b�7��d��yY���J�hNm49y�Ir
� E�������
�W�q5��}�c�-%z�-���C>�Z9s��b@�e հ�P����������&�8q-��^���$i��� �[�p;�O�G��o�ͪVq�K���e;f�3*��Qę]��#��<�eT�p�Y�I�V�^L�T����=�0���g%52$��ڸx��",�#e�6�gFHQH�E��Ƀ�EC�8����u�!�_J%qͷ#�E8���R3��Tl�BYG�M=��'2Ա�RS<7�!��q�+�$�4���G�\�~����e�Ƭ<<'���%͌�Bp�OM[ƺ*�^c��1��.e�2��4�𜏞h�q��-"�ꢎ��`4�|��\̐d|���Q���ܩd7�n�*��ox��_��c�b�pi��I�w������X��T���~p��g�v�H���j� �C��{�(�n2� ��-��B��i���J��[�.�w��� ���2&��]�{�N`�X���p�.�H��Ӕw����V�w�0A�c��;0��?���L+	D� ""2���h�:K0�鑸\��n���V(�'y���A���[��ߖ4�˴�F�{��~�$�Il���i��G�bd���Pyt�D�i��5Nb=���X{�.f�j��l�DΉR��Z�q��z��V�G��Q1����R�-꾵���e(H���˝�Ϊ�ԕC����n��T�[*b��Cq�~��d�,VV�������1(Ͼ:��^��/#�'��
7�����QiW�e�����7U��Oy���k�?��4=o ��]R���M�f|��
T�a�`F����#����$��������|��0}�.�vmK�%��%��kT�^�;��A!vsu�3eb�f(#�)#�kߢ;N�D��ޱ~� ^�����t�yST����1�T �P�vN�������y	�--'�A���,��p��ԧ�6莈U,�����;���/�����Y`�,����x�4%m�U��#;u�� )z�?>J4���M�_�Wۉ�0�W��GK�1h�[�Y��״-��x�S#O�����f@��@�*�ѹOQ�ݱ���W�����@��W'Ԣ��
,�s��kH;O��ʏd��&��H�L�>~��X�C'�&_Gl����z�ʒfI�Qx���D�Ecg5y;��8��cF��E�M�(�.����_����Ș�8�5 5��@8���8�3Ua��JdV_m��N3|�
W��z"�q����&�ap�����"s�O��U�.&���;����U�|��"���un�n��t;�l�g)&��뺩嚯�R]-��?��m�t7s!��0�
I^ϯ�{���D������$�>�D��o�Wg�����T��	٫��QqPP<�T:[�?C���ٓC
e����-�aC9>]?��n��K�	�6���:�MkB7v��+N%����M�i���Rjp�O�l5M��4=Q١�������,��5r l��o�Qxso�.nN1�֜tnm�s���-"e����研������H��R���ݕ�3�,��}GA�ș��0�&2.u}hx�긋�Z#�,@�9��eke��k�Nz�O��>4a\���ِf_ă9ǹ������>E�o���]��ˑ�:��1���ؕk�uv��*�pАr#G� X咡���c⠢$:�����R���d- w*}�y�<ϑ�,�
n��m���&f �:wB���S@g�5w���N`��T=�[����yb�����!������۵B+�d����h߉5%B�\� �������T5t�S��	���Ұ��%�b�{,�@���m_������[
<1�r-�%��ȮN�揬w�[S����ii SQO��W�x�"��}�6tT\�B>�X �8��/��g���C(-����B��nh��:'q�#�ڝ�E*.$��U��ޥ?0x�����(�±�8�+%2� �[�~�=�ئ�^r�Z~AYH���?2ci���BG�O_#��@y�7���+��
�M�	��38%\�_c��t�k ��y�n�]H��)g�)J��̐l�T]f���K�'�;�����$��ڷ-���إ�
.���d��,�����o�'�kd�	�?�~Ĥ���~�P)�F
,�Y�o���\��@��exץ�C �6���j�|�,�$ �*�-�����,���h�LK�2����F ��W_8'Sg�����������ؤР����b��$>ekOE�� !��[^l�i�x�3L?_n�$��uҸvȈ��8���_�A�#�g�i\�wH�r��\/��B�E��O*�F�3�D��/������Cv$�3���[����q:/����dKv�������v�,�3�Y�ރ
0#�M���ޢo�E�B]����I�n] #t���E�B���o���\���v�#f���$�~�͎;:%gr��X��*bMj�,�_P=���*�����0N"�(�e���aUO�p�ͱ\kL?��.��*�i����/�t�%�od:CM))#��=��Y���` ��Rq]����SenS�Ј��s�%��G9��V����}�B����M�22��=x�*�t�]�GL������{6�ho�r�8��tpt�8��υl$�Ž��!�;����	u��0����N%*���뾑�(��`���Ka*�,���K<��oW����|��L�C��JS�tVG���)-\B����9;�Y	_m'�r8��Gz���HY�V�,P�>͊(�q"�y�uH�\���&���F�pv7���5�qc]������}�b7m���H�l�w}�J���]�`+S6xU�J�@-�:�s�r.��t���6�z��I�$�p�jGW�h�ܪ-9C�Dw��ŋ�h��nps/������y��քdq7x�ɣ�R\��{7)�5��!>k�C� TM��JrՅ���쯲�Ί���/)85�*M��m���*�9*��U�޴v�,\�3bϺm��y������x�h��a�p/�wo�t�*��s��eY��eI�E��v��������g��{��������Lt�"Bʚ�����7@�����pŎ}��&n�ݻ	8K���%@1K\��ipW���A����tS��?ƿ/�;L��e��&#_��m8X~�^.Q�4C��Ri�� ��<Hxӛa��]fY���S�xN4�s�x�ʱ��6�=/��Z�H��UL�ԅ�>��#+�'ۑ�b�L����ԡ|=���	���T������ۈ����#��R�Ż�F�l&iL� �+�l�p&��%Ξ�q�<��g��1g3���_��/�v�_��~�m��Pe���ρ�����Ā��G�6Mw���biǡ�`�^u��	�]�O�>܀��!�J�1d����9��7���z�8�2���B��! �*�;��?;�@&�E�qb����F��FmH*��M���p<;�&���޽j&���6""\q�/��R�������c=a2uA�Phs��Ժ
����������$�s})v�5~��u#������B�E�|�=M,�=�#���E�.VZ����#w��H��㏐(�S���7m��c�hċ��d�W5f߿k@���:(E�������("6��@uC jaQ�z���i��G�|�W�Li�t_a*i�m� ���=��;E�X�����Ї��E����)~��͒RЮ�[C��P��r��7�� +��0R2���/�&gʟ�Vpa���Ĭ��E�I��[��uL�_�O��Rk.��"���5i}�^�����h��u�Z@)S��&ܽOw���V%ǻ]d0�����88�ߤ��Y�{�����3�]��] ����o��PZö|.��&f����ż�e��>��R��|ע���	�fy�'���D9���2&T?,�g�yt��7�:F��_;{�D�@�U��߳�8	'x�.��C��0f*�lMi{U!v\���3�z�٨ g ϩ��,؎�E�������F�f�y-$_��4����%����g��2A� �%ǹ��9�ff�U��Q�k2����5�-�!U0@��	'���ɚӕ�D��=tQ�ZE,�^���L�T�(y3�]�&��Єz�@��ѾS��wg��eB����{�p�:R �0�2���RCc��X�������4y`�G�-� �q�{�}�v���!ta���f�0寮B�O���}�S�-ҳ�9��{�!q)�T���M���5�����4��P{\&����ve8R����2Pk�R���L�`��ʷ@gl[���A	�e��P�(=0v!��?�%n�&��Ⰰ��)թ�ь?��+��x����d�&@�B{�")�%۶���1/`8�xX!E<�7�CG{ �H\���;LM~�x�b*�
|�5 �G�V(S�k7�}�ԣ���4���ov��%��'�1��aE���c�����I�Hح�s�tj(]������֍F����h����6e2k��@<P�JBKKM˘�l>��p�n���b"�0y}�eh��(��T��+C�׼�i.nb���Xx��|��5���;��	W��mʻ�:N�S���t�MWc)-�Bcd�&�eKdH�w�Gm��� �O%�J��{�ێ������𷵪�$�8�4�D�(�y�����ǩ���+J�>���F^:vk�M��E�4Ժ��ɣ�,���KiSX���,�l�����J�h����ld2�A�#���<}U�2�޷N���D��=�r��k�RgR�� �e�/���!� $X�_� O�ܺ�� o ��bēN^�wO�%�3�U<2񌗕v�?�M��&d����X�� �5���s!}��+�H����{{�$˘�ݠ5�FX����I��[O�����ݮ���N:�M�-���[C���A��w�H�ٝW��w�zEW�>��IA�G�B V���sW�ə�N骛���o�N|���r��Z�~:�,��1~�(Ư�Kz. "Ls-!��ɿ�OY�D6 �m�q�Ηx�tq$з�Ʋ�_��b��Z���������:�~�/�8�)4O��� ��ne����!9��I�sr�V�!Z\6�vr��?S&�����ݗ��	D���K����[����Q�ڰ*<�A�閹��=�i�����*�O��������¶�|"i(d��92��,`ͱ>)DU�/ь���|�����{ހVG�AI��d��Q���[L�L~%���I�Y�g�(0W�/�XׯN�G{����X6I�|M���	6��̆ؼ����K\� B�P���	��M���ݏI;N�>�
:�>��B�$EPzg�rD�ef���f�hy��V��ː��s�K�ϴ�#��#�&���$;�͇�tN��,XuK�V�TJ�D�&2Ŵxj���bu������es��T�s:sü��8������{r�z	��Z�n(��>H��U\�Z䡔8�!Nm"#Щ�E�k��)u���Sa�s;�R�_����vEB�_�[c���w������F�r^_B�S�=*I[ZX��\//龱�p܇:i�´�ݺ����G����}��%�&�^[�ʴ��#&Q����7`�f�����2�zu�c��.�u��ә�$���x2+Su$��vP���Yu�<(PPDl�[=B�p�X�AY�BR�_����k�k���:��@k漺?��b�G�3�rf�J4�~%6v���G�k�D�J��ELʍ
�'�#�M��/�LGզ	H�ɔ�ׄ9f�ד�@-x���P%�C6�ĄvU�!l"�b�v=�eV?�} �N�K� �D��_�J�ၜ���3YO�� XqM�3<�����Ux�t&��6;������Gm���з��a�H�_�G���5�V����U`�&:��<~�� ��g�ϠZ�QY�,!Q�ƒu��,z���Nt��n+�(I���+�4�(3���b2d�G�9 8�1�t;`Wt�����wq�0���s3֕�V�:��W�P�CV�c�^�ôPu��Y=+�6SN�TѩK�l7y97��I�����"Wݗy�IE[�>;S�&�$���ט�����*̚L�%BQ��B�wI�j8�)�<;�Z��7��/��#*���wG��_E�B��2p�^K� 2�bݕ-��K�����̭K�t��oZ�3��s�PB!���]��`7�Y�k�="��1X5}����o����ԬG¶�,�.E6J��Qz��(��ҷ��!����'�b�G��gsr�qM� :d	��R�;<�zJ]>pi���>Q�hǥ�0x8`8[L$fnɩ��Ik� J5���� wS�ぢ).��p�������z�I`2�%��d���T����q䲽
�� Q7�y6�P���h̳��O|wӬ�m�58�]�B�X⍛�z��_�������a?���:=����\���$��RG��h{{�hD$@��UΈ �iK�H�>�r��m��izD���b�-�6:��}Ib�������?bO�|��Q�����!�oĜf&w�no�<����F�Yg���� 6TC��l���n������:������:��H��b�j�Lf�)I�i/�������Cm`Bl���U�y��!�yw֥}�I��v��p�!|���a�omyVA4���-�M�N0ǎ�*֫�Q[�x[��m�!荎�H��"3��2ot&c���I��4ѳ��>j�S�]Y�zR����+���r��7Rz5���x��﨏��HWE@%䦛3n�}I�����	�T�� �N@�7(0���2�8�S�	����G�B�T6�Ǹ?Z�
l0��j��u{�2��pv|_�MϨN-� ���%�Odh0��?r�(�2T���M���=�K"�r&�ۜi��Ѿw�Y�����{9�Y�QpA�Ȕ��WqdO�s�+m6Q���ـ���`	Y��j�+m�tة��L���#mv ,�C7�Z�b�X>Ň�'�6�i�Q!���W��ʆu!�s��*���I���+h��j
���ghRF3�_F����]x���X�������;�z1�!#�K��g�߻	���z�ߊ�[������67�t�,h�=[e۞b�g�e.V�Ј�w����AN��_�\6���<S?��Z�k��!��C�p1l)>	U3�Iz�YSD�F6�T�0�ł�_�e�2�/u�]>��R\����P�������͌�|����ɺ���D�}l����5��?�ǗD�=Ԍ���A��ԅI���W2
��@��	jqSA� ��:�+�����Ή�p���?�]��j���F�I��I��.cT��kk�]�t�s��u��
d��#EV�!�l���o���I�ع#[���;���M�h��Nm9����M����J^Gz��Yr)�k�m���w*Hu9R��l}�ـ���Fё��F�>�B)�1��}VJr�fja�o	�0e���He��ݑ�:k��4$�b�`Dw�H��R�J�i��6Ȑ�n��-��խ���9K�@�1�����鵸h�  � ���ޭ�fĪ�1�����tUQ)4�no���y��X�`g1&�j��i@=3�|�F�����R2l�+�qLj"���k�������֩��'H~_L�J�����+�MUY�E{�'=hv.9��{۴9򪤫��� l��ޚ!�/쨲�C�J��|[�"����
�b�~:L1/T/�c�zK� �8;y�� �	�O�λG������6��\u3?�����F�P����(�;�o{��p&�ԝh�|׫<�m̅H�^U,�W��[��6���ZDt�bN���Tk�0g@_^#Id��ݒ���jC�[���l�B+�@��Mm9NVݑB~�o���*!���8�B��o�I쓏Jl��@�O)��3@�*�ͯ����Z.C3н!qt��[ ��@���:��g�tGK��.#��~�A&Ʀ���)2�$3Y�ρ �1��)yJG��$]8w;ڼv[�)��W���Iۿ37�S�g��Z#o;"��D۟�A*��6$,f��
��?!�  f+����Ұ��1�nj�4��#�vճT�ӣ��+1Q&�vN���:_iJ���5�������<���J7�̜��_)�ּ�=��'.�	[/hU!�������!x�����-����r�i��*����F��v���X<ܟ���э5'��A����y���Y�$]�\Z�G��JG?/�x�{JM��aN�Bxw*if#���}rȺ1�4��+�Y��.5ZQϞ� r`f�����Yyj��0p�W^Ţ�0HF/[�3+qŶ�����ꭇj&�����>�,Oްl��X�8:�f�`�푷g;�;}���)~��`g)��N9�U�{I=�ۖ�a�4h`�V��ٓ���+K���j�v6�n]�>���	�q �������j�+�!@�$`��V��SĲS����\Ii��~�xOe2�Oq���v�p�N&�DS:;I�	�!̿fٚ{N�yX�Ph�'���_oe�:��^<_Y�8�'��r�>\�!�� ܱ�jjO1,��w++L%u���dE���8�Mf#-��u��/�j�������a'��p������\�i7�E���K˝9�_v���kE]=ҪZ�����= ���D=��T ���ע��/����Y<�)B�<u9��ɣ�rb%�|z-���xI���f0JH5[������ �AF�l�X��G��i�l�	��/���ڣ�T���Fr1�.L>&�U,s��S�.��*g�+��b�wT2mz�� hTݦ} =nEV$�g�0�P�rQz`�9&x�i�������Mj]p���d��*���p>�c�GE�R�T��g�K���7�����/v[Hњ&%��Ҙ������Y��R�|�O�D����~���T��+X>h�?R�Y�D�Wp����0�wg�T�ϗ�K�i�{CpK��J�y�赨� �n��T���M���2X�I����p�܏q�v��'Ip�a�K�����`�p�'�(�jP~�Gx׷m�Cu4��(�
�@�~�	GV��PͶ�.�E���0����,A� ��Bc�\
B��CL�)��
�L�6�W�DW#vYD\��8X��Õ1/�f%R�䱭��r��luITH����m����׮�hK�jZ�O�N�i��(�������� �6�i��e�+gǹ����(��Ԝ�����"��,mnz#>�{eƭ��S��?��mY4��:uKB����.������np?�]�sGCU|�����/�1U�,�k;�qyǞb��9r�GDHd���"�0
����O�@I8�f���J�M5�ꪘ 	h��<a��Q���o�<<��r��J6�ޣzn5�+X�TҪ`$�O���0.�Q�t��x�re1��5bmW��D)K,���h�Zh��x���,�Sl����P�r�'���Ԥ��5�>�T@�|l�h%��~[�'E�n�2���GRt����U� /�A��$�#����F��aLg���j�q�q���YʦqO��,iĝik~mT��O�Z���������klR<ƪ|=%X�l�~r�;��
Oki�Y���0,�s��-R�K��c������gP�4���-�)S$Pe�D��C��3!�AX1�%)�i:YT��H%��������x�y��{˛!j�$=c�"���ȕ�I������]�y��0y�D�ր��5���Q�x��Y�\�� �l��=�S�ۄ�4���dj����5��%v��]��u� �����-&��6�F:/?��؊ u��ydxz�V��~��2x'�����n�+wq�e�-@?�G�����9D���'s''[�L��.Y���޽��T{�?�[(F��F��Z7��<eJP+�=������`�b���������)&�c��Bv4Q����2DY0;EL�뱇/�-A�0�V��dZ2��/R;�?��!������ 6��
MoT�,4l�_�-=��1h�(�!b*�*�e[`E�!Ti�<p��(�}�(8��.Bj��`�=��!�ٙ'��֋C�y%���\�O7�>��!�ik�������=��m~����� m39�؇	��9e�}�4�c�ʎ�u.E`	�	�l[� ���f�u�jg�_��S��wmO<�!� 1H�Ñ/���� 0<��X��OM���/��/�B._x\���n�B�,�9A�n�|5�3���a�Y���J��q�5�s��}|� ݡJ�c:fAY� 3�����^�R0O��]w��凁Tx]\g
ĉ�qc؎a@�(B��T���1u&�sqsN��Nw��*n��Ƣ���	?� �$�60��_#�GLD��^BT���˶����_={�;�[韻�Bi�(l�=��C��׹z�QC��~�*�w^�-�S��*�)t*h���O=H��h�D�g�!�t>�O}��
\^�EH����Ya��̫ |o�!�5�s��8=aZ߹w����ţ�I�̞�=O�w�^?:"B�Z�/�����N�җU܇�K�%\��_J�9�$��y�7A�V��P_���!�H�#�\�\���m�7�@wj��I|�g�K\��WnE&驂�����Rx��7����ef"ʝV�8���5�x)��9��h�Y'�DϞA	H2�E�6v��}���(�Q�	�x/��9��Ԍ(��6'��7��!�+�Sޤ��A��X>�.?Z*�\�7�<>������&C�0���N{RM�-�Z����:�L�$9�L�z�q±2��i�_U�1�5�:��b������~��W;��R����4��;�R���	,�k�b޽�W���(�Vi}#V�$�0�,�c6���9��C�g�E-Tn(qɧ؛���- �<�r�g�2�kИEd�%5߽�3)B�:
d�m	���R�����V�8#F"Qk�P�*݊���䄇�吂��=���KV�޹G���Z��T��tԧ��j��??J���6�Jނ�0�,m��xT>6P��&��6nF���&��t����>ŭ����h�V�c����ݘ�(5Z����̫�&�˻P�L�"V�h[Kj��õ��Biy+Y�`�*��@�`��>�o���\Oi�\�NZ�a�ҡ����t"o��3��#Ņ(	�w%��܍l��n�"��Ԋ��9�PG���o$�f�D\O.IJ�bG�h��T�
�"�0�+򯫣�
�)��-j��Tx����d���P��0�\VG-1�(�P	�{��ȏz-�/�ޘ�L��)���j'���bE
vdg�)s�o�&�]����Z��K3��� �󝍿+-)e�� e0W?�T�NOk�*��]ս}��wI^?a�q���Dz�I;x^����cgV�6�9�,K��8��*�������q�6q�=��������[�%�I�Ehu5f��z<v������Tb��"�G7��`&<��;���c�&u}̰	$PV*_���qK)Ԝ����a94��-�)5W��w���D��	Hu+�i
p]�U,��Pe�r�f���{���D�E�����Zy���ӎǞ�G��x?�7�Q?;��)���o@�M$�����^����X����u�̎��.� S��֒���_iLm�7#�E��C�����R�RC<jIN�������,m�`�S0���n��'��q��`}A�AP�JRK�<�Gj��v{Y�������-�U��]^S�w�]�ȶB'���x�7�~wlO�ǫhl�&:o;�9n�_���g���~)�!�Sz�5g�����.���FZ&v��S�����E�^̀����"�:��n����b��q~e�gΒf����w��_���"�!�V�����/h�*�v$ y#���Q�F�]���E��������{c�����7�r:9�&�zP����6w�K�@G���/g����M�R!N�����gH�m{G��/���u�Dz�v�sO�����f�"�q�w��6(H5I@g�����4� 0N�����2���
Y5��4��{�v䀧�l��/�Z���A��z�`��򛓫�=ufHS����S�
tE$b	��K�@O�:�0~�b��U�p����V�	�z��ͼ��ķ�eˈ�6���_���ӊI�zC%���P��X��["��:rK
d
���V��A=z�[L{��K|K11>�F)s��b�}�.:w�jqJ�d�8��\sZ\m���ti�7`�<��rl�u-�ITm����������R�uE�b��X͒N�Fڟ�������P?[������uO)�?�����eOT>�33�%�shv�7�]m����)�h�Zj��m��4(J��>r���K��+��P�[�2'>"��;<����ק^)����8�w�4z-b�K���� �1m��{�V�ޔ�~�-�w�yv��LF���Cm�'�O�b. �χ;���dx��L���Ov 㟹vt�ϙY#�:^����H+�ۉ[���1�G���a�j�%��^��s��5M��ƶ��uir<��T�Lrx�ț���M����F#�Mo�����Y�Di;���0�K�BC�E�+�0|��{$�҂c^Q~�mLBP/�7���)�1��̀6=D�&�%V�x�b�c{"�P��0�K��P�y�v%�ʘ=�9��*q�\�loXDD��?2�X�����x��4�6���%�L{��pp��A�EC�R���SY]:E{@�pf'(i*ً����ڸkLaj?1JQ�+�����AP��nL3'=��7���9��(��9�<�d���EJ��=沜��hz�5�BwzS�M����{��i?�1�	Wn�y��~���@&�h�]1i!�K1\yc�_�x�v[�p���+����~�`�L�g;|�g4�G���/�{A��js>��]˸ŉ����
�6�*���J
��{k��*�l� z�I\��CL�iAЗ�l��"D��x�v�lxDy��������ȵmT�)�|0g�Щ8KMLX�����W�b=�ޢ�P���w}�hֆ/��sx�2��q��b��^B=���0Zru΃��g OSx�m����� ��VN-@:�� ����C`�AdKN�td��S"���y@�+���[��+����	��ˠ�g������ot�;���f��2yV�<
F;d���ZLW1�5�>h4p/ۊ���D
7R���R-���:�,ԵEL���tμ�-�Z?18��_�X��_����3=/[ۦXyqz�4��^S=��Ip��_RrÌ@m�K�9)M�ž\�f�ٶ;r<0����T2��W��lĿi�Y� �-�_�DLxqk�������-$Eʥ��VC�l��u@��O�d�w�\̪��o���=�I͍����i�jw�~H�c�0�J�=�#p��H���(���M"�o�� 8Vn��1ʃ-�r�jD�/
�T	w�iTEJJ�_�f��$7�IJ'Ԃ��,+�x���H�0�m�<BV�?M/@�U^<g�����3.	�TqK��A�s�7����!�\��D������B�.Ջ/n�o����3�DE���Š
���/��r�32�h;�̡�����-k���/����w\�m�L��`oƔ$�T �6A�g�_?�a!�#�q��ӵZF
���͈9~i3�S ���I��%��I��Z+�ڼ�EUaډл�pA`��U�z�����7"������8r���ށ�<Ձ���W"��+Lu�ʞ�"�����Ez�J�M���A�2	A�xr+�B��p�rB
D4GPӿ1�eَ��r&��7Ƈ�-�E�wB8� (�_;���zg�ͯ5�wj,��e�G���ص���ս�J�kDB��Yld��s���e�3�`{�#Rd� ��dN�N�%�%{b�f�Ae�σqP��0��3��6YD,V��B,����bER�C=��^�[뽣�0>du�\��OG�<�\����N��.Moj#L�yt���,ݥ�b)[ޓ�K��P�.�(ȷ��d�*��*��땖*������5HS�\R8X9�;�^UPDuy�G��Q�5I��P4�B��"�C��r[4�C��Gc�f���-�D�W� ��sȮ9�xE®�~Ik��*h���J#�	�A�E�ܥ��빾Y�Ͼ3�Ӹ�(�q���G��;��Q�]D�5�[tK6�mc�y� ���Z�ŧ;�n�A��Q0�Q�N��n���yF����?�2�������.L!4��֗�D�g��&k:ך�i���=��ۺF�5!:k1[$J>�v��$���x�*0�=�hz�e ���D@T�L8�ls}�S�I�V��㽅�$ �딹1iG\PrF}u4�V�������.�Yc<e�}5�� ��L]�P.����X2c�%p�<�G����&<�:��:�wյޑ�M��_��� �q^eX��ֹK:�B��?��i�	�5��W
����L�99���kw\,��g���mQ���bh+?��R1v���
=�u��od|��G�&y;nq4V|���ϔ���	��GKcp̫p�*���gY*�͞ޱ]��z�v�ĕ@,lk�(]��́b	h���zjBV��OTb�b��6�H�kѤb���U�,��b���L�Sp�T�c˂!]b��J̈́pk�²�%H�:��Ɏt"<\���Tu#�W	W�T����s�ɑ1E
B���<.gt`�����k�Pkk�:<���P*
J\��������כg lD�L^�;�RN���"��A.���8q{�Q��-�3��Qe�-~*�z9"/΢�ה���bp�>��6荊�a ��=E�-�}�~�����B�4���M�ͻ,����U`��G{N�Ɉ�A��tg:^�螴ؕM��{��^YQ$R��I��Q��,xN�!�5�F����"AD��+��#N�Q>�<t�N�J1:��`����V�g�J�����A�֋/Y�����;�F�.����\��n�^v8��P	��m��vzg@`(��9�U��.�ji^�B�����RO�C��v��7��:Fn�0���S3�q'�m�K�ůS�VƉw9�����v�A�|��\B��쀨Z��v*���������j����1�?�3�}�����/����EeA�m�)�{|6�F�7��m�+�E�<@`�L���+���*���q�>'x@�����XZ�M�w(��7��I������Q'�YS��9�Ah���ɖ)��0}n�[�)�]���a���6�<�<� v��N�;W�7o7���^�.��{Dcf��"�{S¹L���	!�`?�����>��=?��*%��h)���
'N[z7��H�+S�k��T| �-R��{��X�D�R�%�!^eM���L�F���y@j&%1S���L!r	�NAh��]h��G�ġ������aϞ��%��56�A������&���$Ϧ�n$�
Kl�A�S��#�rZ:�^��f�g/��Q=0�poj�xV����Q;��d3��>�����b?a̦F�-���b�r)$�Sm0E��2\GT�$��*���0�r��}����1�3H�4��b���e�����T��68J�O�y�7	��(�)����c�Nͷ��T�
�G6��b��1�P�2곩j�tI~�(���銫�����~q"X]� x������7�@���j�P��~=ŸC��(���6��kkMӶ��G�a���Dg���X86�jW����U��C�pJy\>��ūG���I��r+��O�z�R����}�y�S���472Z��Q�fF�W��/�	����d��$� �+b�b{I�ldܭ�\�^E��bg�xZm������ޞЎ�N8�l7��2�����fZޏy��4F\<��BN5Ik��Uxׁ��F71x�Pq|���m��Bmģ~{ޞ�`i�I@A�&㲴G�L���� [������P��3>�
��J5�s��4�gay(^����t=�%�"����]�g�a���D��ͥ6��l;� �h������2�A.��#��[g4�v?Ӎ ?���{c��\ɵ
x�(,�.V�!�^�'#�"6 J=pGԲVTc?��1���hퟌX˫��o���Z��SK��[�yu�yc��n���������2�XZ�ɈtI�8·��P���'_���G~	R����H�)�U�[צ ����#e��?��_�# :��� ��t�����:�	7�ʻS&ze�dϔ+�pa�BP!bcc���$O�m��I������\�dm�~Im���G�5��]b�^\2�<sL���&iAE3dbhS��̜��@������OM���h�#w壒�I��$v��3d���F?�E��ev��e8�J�𡯲8F���⭑a�ƕ��E,#ji�]���z�F\�����	�f�j#�;6e���=��n�7:��\|!�������D-ދ30��
��[� r��4�m8] �)q=Ǵ������f�9��ҷ���;�@�Wg���*�X;��WW�����-:���A+�gF�jS�G���hai��4��]"a�ˁ�_H�A`��oi��rg����w�l-h}#o�y���#T�d0H��維	�@V'u�*(���yA�"����S*��9<-!�Bt�iؼ_ �]�0x��N�fm���w���X�^G6�&��N�d���Q'5T�3�ʇ�bjrh��8�4�2�n���~9���8"��Oe�����DHwTK���m	|���c�%�֭"��($i��hQ��-��m���t�Q����d���ߒo��{��.�dԪ�[9j�� g����EO!",S�WV��k��	k�5��ڦv��]l�R7�=*+a���J��#�KdrB(�"/���r�}j�rr:���9�CѨr��������D������N�q����tJDc��)���yu1k��a���e{l��C
BO��[jZp�#����ٗ��+��j������{a2b"�����\>�g���NY��au��!i�;�火^K�hI�^�/�E�u���&�_t`�р�;Մ^)�;��{m`9'�x�?7���-|>�q>ˉ`GR V2�4�W�Ǳ�R��9�m�����	��tk\
��>�Q��Q��"���AeP����������i�h�V6U}|H�9���V�egP��p�OqQ�k���	��~����u�q"��7����z��Q����ܠQ�5�@�L�����4��Ss2���qZ�������@t&�s({�w�K{Ol A���+\4�C)���	��/�'O쒧:�-v�#zǛ�H�7��
�"l��'=ZtO3mʂ�;g����5�W0���Ew6�K9�cM.����!}�?���H��W���hewЇ�hs/�k���j���`<4X(�W8{�4�C�u�Jx:j�d�89HQ��gۉ%�'��ϭ�n�Ja�s,b�b���/Ͻ�=M6N�I8m��޿?Z��`�ɻ���k���ޠ�I�"���J{���cǋ��Q�����p�t�����J[x���mnW�~b�g�J���TV�qP�w~��\Q�{�C��+�z�ֻH]���C�B�Bd��,������ӭ��<V�^ ��SQyЩXߚ��+��ئ�c�?�s��[7~�B$�u�P�u���䊯��śi��3?rdH\�Z̅ʪ����'�e�$?�:�W�H3�+L�Z������xf� �*���.�"�a��=5���{6��X�g��EV���%�y��N��'��]��ϱ��)r2�{�jr��{=��[��L���9�D�	����fG�UsϳWx�ť�Q�P_�F�CL$l���eD����ħ���f�;c#(QJT	0����hqL{�I�K;LvДe(W�1\%1��t�� B3�F���nn�b�F�|Q��E�/
�~�ҁ��/�c5��8��Z��z��ܫ:���_�Xg6���^p�Rqb�.*�f��9�������F8�-��ٟ7�#x�ւ���տ����e05o�G�\���/�2�h�A:yuU8xU��A<� I�i�S{ɸA	W�B�,��EP� 2�d���v�n+�o���j�T�p��l�Yf���!�u�N)*��B~�_��[������c?��5K̽+G��L���1���F� ����5)Ǵ�wc=i�i�����<|gD��B��Z��N�[/#���Յ3˴��W�����5��i��?[(�㾰�TL'F,���f$�.�SҏRCYj����/��Tr8�JL� k+ܨϼ���b�,���L^�|T�+nv�a L(�]ᶫ7F�4Cg�4#��'b9'6IL��n�H���{Bf�������6��Y،��"��W�Nx8~#u����8�NoI����1���M�;|V�v���\p�������҄yS-|x���F$Qd�XfL:~>�_#mħ���dM����ɶ�0��i��n��X<��{�p���)��f.5C�x6���3��8�>��aQDy���Q��Dg������P��F�� �%  ��<r/���Ù��Cn=�t\+ �����]?���
����;l�B]Z+QL� x�	g҅��O-p���������®�G�r�W�W��~���
˵Vm�kZF��+i��!�ի��K	�j��!�K�����\��s�	2(��t5ƞ��A�SU4a�dL��y��qa)ȩ��<��E^rJg�H�X}�����-� �v�B�DY�:�/+u2 �o���+��;_ɦ?K�ݱ����=V�17�3H5��;��2��>�'�m��M��kv�@�G�`-�<r��t���3s����rMy�����	,s :�^�k��xV� ��h��#�,k��sU��gL�ݿ�\�i�DE�2l�)*��1bc[�	XO��Wf�O��'I �^%ca�nsV�y�նU��6&�	5X�:'��D9������eoA�6�
W#�Gk���)�0�ULxW����d���׋7qnҨɫtd�?����;�8��sf�JO�]zp���Г,���I����H��{|_�o^!˨~���r��CUd\�w#���%,4������=��(u9� �L[�HbJ� 4��D��(_lF���;nQ�	ټơ��/�F�I�����P^��o�L�r��65$�eeN��nTO|��W[[S�:v+���r~s*3		٧�t�񍨷.����-��Vc-0��+�<˧�iQ��-�V(@qs�X�N m4VZJ���O~�#�k�Խi�4]��9G$�,���UkhQʿz��	�-}c;�Bj���4CӢ�"Ծ�LdGܣ��^>�A�q=��#7%aoXPv����4�l�8٧���5b8"W#L��i��b�>"b�G�b��0�*����Z�]�7yޚ�̈��cc�G��zw".��X��!!�����0\�A_��(�·������`ZҤ�F���c%N��#�����~�L�(i�m��	I�����&�*��UYn����R}6,��i��q�����ǉ�K��WbM��]7�ʈwy��}42��
-���фIy����+�:Ǘ ��NM�^X�ŗ%g�ⱋ\���b_,z|Bs7�d��D�C4��RBzlREJs[��D�F|��adp��m���$>1j�dv��j����v�H�ؔ�a��C��^`��f��|���1n�a��T�Y=��2��;?;�"�]�(5��{={F��*7^�X�|Q+�ī�|���?�ȑ����ϕ.M����`�+�Sz�?��7A�*�Iq�|c)'LR�uzgT켌���B�߻x7�Q�WR�<2C�xw�X�`�c;��ҝ`����.�i|���|��뻑��G�G*+(��gW�>��0��T@�i�{;%̬�1ཤJ/�L�P:('�*�!&���?l�ß�.����_h�|��� 0Zbq�(zhSz����v���aՠ�>����D��[�I���Ba��N��h\�+����#����P�ȹk_�!��h!���O�,6�|���<�Dʁ�锧�UYu���J-fn�d��*@�L���f��j5w���w��̦����5&�6� q�G���$L}��|��/%��s&��v�*��dNz�eU��,�������ucs������6����e�:�܊���s@TD��R4B��۝5ђ���iFhmc#S@�ϣ�$b'b��dv�b��@[8��·
��k{h�~�),��T|5�!`�.9�7��� 1�vSU�)������T�a`>	���N�&�wǬUQ��-TC7�p�W��`-N20y�axM;\����@!z:�o���%��[]at�����~F�����֑O���ɛHƼ�ɂ�3��A�k0
����T�w�1�բ���v
a�;��1�g	�9�����~C?S��a����܈�-�,�g���s�a���s���_X����R�ҿN��������..I�]k@ᨏ|I�$�K�!t�bO sCaS�C�JQ�� ����ہ��D=ӆ�H๦MV�ٲ� �I2�:���m^�yR]�)�y O�+T�*�d�?_��~!�9��	R�Sꆸ���%(��y�MC�>����F�h���j��>�Æ�p�^#LI8��`=�G���E����%�0��b[�RBD��d:?d[���S%�S�������@�*65��X���V�S7>P�8��o�K����"�7GS��w}�'B�K��<'�T��W�4�3������U���K
�I~����9��qU:�z�� !7�◡e��L��]�)M��t&�L[���	,0嬝َ.��� ������
9�-���=��Ě��u)Z(�&���.������?�Y�eo�(@�9*�VJ�h�6�h�`�9�o�M\fg˦73�߲ӚI�T;3D�X�9Jʔ�W�z{��zIS��~���3�q�+ꭌ��D�q��.X[2C;�:K��h�����89nX!ǒR-�ܒ��x�7 ���$�U��ZL�	Wʥݞ5���0$����T9H���4L��L�*9�I�e����,�"�̫:�sF��Ch���2AiEU�iQ3��l��\+K���T"�,���m������Ň�a�5�.���e����UGXԧ������j�,��)���X��-R�+�3���QW�� ���C�U�6����ja�� ��z�`"O��W���h��!��hwz0\�k�	�7���6j3/u�D64S�(/F�o㪸-�YЈ�f������✀�k��f�6�#��r��&֖��}m���'���Û{q �1��CSބ��ᜐ61�X X���ӿ�w�ǫ�@d��������c�k/�;+���~m9nI'n0��H���E��t�����]ZZ!�ug���WF�<�a&H�4L�}~�T ���z�P�Q�U��o�f��5BrF��Q@EcF=5�E����4f{���L58�O�I���<��O�e��/��d�����򑗬�͵g�Oκ��D������<(-5�� r�v9x0�E��F$9-�g0��S�t��:�B;��ջM��3b�	�,������d$ܬ�c?�Gx�O$
�l�*e\�(�^:K���0t�F�{�"�2{�O$��(��@�~�G�n	�?;/o^���)�YyɤiH|xn�
���:RZh�;��I���F��7�p�x̀�H�rZN$E�Ջkma_�-�QY�T�F�����{4���r�UD1��s,�sP`�_��Τ\��Z�}�n���-�ݐ����ٙ��Kp�v!�gS�z�u��c��㋰+,f�&�@�/��h�|�(�T��p���*L��������&Ĩ��\ez�&h�M�F��؁OwH�bQ�!!~�a�����}G���[���`+B����5˥C�oNͿ����U5��2�|}O��z�J�
U���Y����wg��X���儱@�#Jk�Aj�+M&���nL�-�L��x���t=��QF�����1�a�
��B�#�K#�#�7� $�o���P�6)|����m��P��h�,�x]��91w��LQ��7a@4V���Μ�mDQ�H샛�OY�D��a�]U�>],�T�i�U��,sv�'�C��yP��Б0�C�A����İ8n�v8��q<vAR��5�����d����^�P�������A�ֹ�9�$�&��h0��N���ʝ��I��� �Uv�0�CR/h�5�{�
#Et0�'��� ��pA�+/8�sg��HUk����G�5ݪ�X��a��K\�w�8�%�y$��O�ѓR�R����L�텽�$�ý\�#JU[�WH�w9-�^�ٌ}��O.�/�+�ؾ�]M�<ƊH�/:�{��1�s�ʞ�E�ue�$���t��&h)�?�x㐕�[�Ib�A�C����~�z���o�7��M�1�2��ڀ��?�ڐ����:q��Ѯ^p84:��C`�;�g/RYS�&�X�~�'͠��F8:A~]�HpW�ě��u�,�@��k�Z�裛�֒��=���p�S�\�Q^fz0� t�^S�����$���/l��(�Ր�ҍ�O��a������-�'޲_��b.z>�wY@+�M,u@��3�rT6�}�=ʍb�0����DF��ie�����΢�~F�*I/5�FM��g���ZN��Q6�35<��nan���5�v�C���]�A!i��1xx��	b����|{+	&=��˩KK~PO)*�Yj��(���^Z�ޭX/M7�6���&Rv�T���L�0���ΫwC�Qԓ��Mq��Ao�'%�TH�׭���$���t��2�j��q��,����O��@�F�1�}���4`酊5հjA�W�\��m�w�(٠G�Pb��m��*]n�I�c���"�|.����.����03����dC�0�`zI ������`���K9�˓���ġg�"kR2F_���AFD �V�M�$q&A��c@�֜u���4�e;!�n�����օ<7O*��#Ptvٕ�Z��9Vx�332%m�*�VBR��P0c���D��/� �c��JP��;&>��K��R^NRT�����5�)Ә(�vlX�����DȂ(Lt���&�3�q^�PƏ<|e�ݫSm��{i�*�ڿ��hU�e�"�L!&;Y�\û[��� ��#������DEՍ��#��l9�{.�.�B���_�<�d���Oʡ���hY�	���t�M�4U"�}�%q
%w"=4�hSq��ebܚ(I���~	��@��Z�����:�`@���OJ�`��N3Eԇ�lq25��[�����É�1�o����q23[���O�;Cz���ULU�4(�c�?zm~�M�NxA�h�2E����'����"�֍Mw�=��͝��O�����c�%�dr9�K
��<U�ly� �vly(f��n�@Yr�$8)�10{�H�i??xg�������1��1 %y8?�E>a� ��d ������u�F��{�2#a }5��L���s������jS��f����R#%���I������-Nmm�.�a��Z?���κȅ�0@�y�짔5o��W{�3 ��@����	�pu�!��whz=}9V��b�̮fC�$ �%�fa�߲�����S������֞6�G��ygJ�_:��=�4�M���lu/^r�R;��������,	F����%li�d��s�w�W�P�< �c���y�K��䭡|���Qq�0��<��:�y𮋲uRdx0B߈G�r̯���+��y'vQ`�������V<VL��:z�^�`�w-�	f|-�M�g|��)�6j
\�1�jf�בC��;Rb{t�m�����DK�CV6/-gz�N2�8�\��wK�SբR�@X���Px!�}�@_�y-�TB6'�
�nH��àP���9�?��	Yc2m2��E������V�Ւ�������ENB����#v>�!>V��x�����an�I���T���¢ C/�Ԥ��n�x����2dZi�릋�*��\}
��)��F%�o���'�il��Lz;	��k;����sg'O�xCpG�����~�|\ѫ��^^F�m:n�7�������)�9�F�Z�3}��8� �}����$�5#�����x���@�V�<�1�'�JQ<�GOۼ��~gz�r��1�k��"�ژFkTJ���}^΋-��7����@z�{x���u�f���Sm��N��!B{�ks��Ww)���P�_n��<C�IiZH`�9m����y<�m)�ٺ�J���y`�y���#�]k�h�,j�_�����'a<
K�c$,5�?��=���3{VW�v�I_��_�?T�4�� \��T��%}��� �I��^5���L�B��͏�	���K�.���D�M������^�X���O�I���* ~<��ۚ�@�^�Y����\fS��cR���� c���:��5����=���l����̸�<�5-Q����C�� ��Z�zM�M7�|��R�R�*tzS��Y������Ħ��4�ŘT�W  �y.᳟�֊�wL��3Q3�E����]��ug�5��A��k��S�i?���
}����Frd,�� K�x ����-c\��k���:��韋߸�a!_���dH@��R,(�B�^Rvi��[� ����6¿��I߹�G{�	ɖ��$��C-Q+���2��J#��UrC�Q��Den���(�`%������nZ�t�[��v.&�gQ�~D9jO'%�����o���v�����+��q�Q��3a�]:iv0q�V߾�O�2yG�W����0�� ��iq�
��\cd�/��.��Ҍ�H��`���~=S�<��Tjߝ{8Y�:4��D�����U���(�cEB���/���r�1��#��j�uY,gw�ZB�ُIe��6���䏋ҟF�>=��G�7걳&dǞ�	��jʂ+_�~}�&'��sN��&���x�ܱ���{��� + ���"��*�v���vo�N6	�As��io�b����^s����w4�� 7h����%]#�����.��g�GGĪe8I���R�L�WGv2�*C�]-sX�~�lWE�rs�'�Ww�˟�O�p���1��7�hx�3�hO�1�A�#�U%*Պ��ɠ}����\�^V`Ab��0��%��#��*)�X#�T������R�Ft	{�C���ڟ���1���8;<ǔ��	#<uf	�T��Bf�@�=N��lp���P�j�^@�˖���}m#bQ�
�2��7y��P��Z��Æ���X���SWʕTʡ�� �������B��sY	��!4���9�����ۦX;�t����c���#
���ӂG4/6�!۲�uD�����ūC,�Ir�j�ҵ�w�������-?�9���aˑynC�Ϲ\���:���
��#�v'�	�ʯ��5EI���O�H�ݡ�W���$[��Ƹ ׏�_�@�g��J82A�"#�����ҐSW�B5_�X�����K\�O���?�ZY��%�� �]��6(
_:ы�k��.�{S��?u|�G�!��6��è�(�[����C��������VW�-��9��%�xf�h�/t}�!1���nF��vo�O5����6�J���Y=߭/�='G��X�'��~����ݿ�|V�XsY�.���{k}��F-+ʀ0��9�;���D�ӷע�V12]�d5�U�A�së��TGSpG�@汊t$S�y�ȉ�I��� ڎ[�dX�Y0j��9s8A�dH��M�)m�Ӄ�hLd������R*�Q��s�e56��Դ�W���~rs6��A\�}���:s+QU3���pJ��� ��>��X�I7��
�~M�Ѧp�W�ߞ�6zo����R����+E?m�}d�n��X��\��[�\��2	E{$Z��>��<�e,�aM�_�S�$	�p#¥�YJV�0�����Њ���Ќe�*r�tQ:�d��Ɲ�h��_��]Xyc����We�"�
�� �6�:��5`T�?�Rc-��HO}E�5��~ӊ��7��D5��w�7M���A��F��Şx��+�6ɿ��#[�ʕ豟�����;>�6�1���VW��ֵ]��������#u�dv�
��4$�[L"Hs�z��l�Z�&g����0 �#��	ڗf'�^$�iz�z�˞�|%˟"�3�;�n#C��_$�6��%(���if��/��呹L�PܴJ�I�[���:��q�f���4c���Yu.�д�xl�U71k\�.� �Wy��������P)���x���������εn�}1�����+��=����x뢵1늇Tm�P���e�u���;��FNψ�x� T��7}d 3XU�z�0UJ�INs]w"��c�?(��\s`�x�v��!z �7O���7��Q����A���}̤���W������a"��D`Wa���*�����=ri��I�@���}"IZ���I�]uTu�~�;�R~�_���2	,�	{ikƾ=��G��\|�Ul���!��m�����^?��O�+���+�j}w��-d�y�p���TиVJaٹ�������ϐ)���4�u�c��Pz)��ݥk�R�L�����T��l�Tm�h��$��]�G��F���E���3��^ �Tp)��O�D��+�E�8 ���{.�}�5J�[+��З�H\�N�~�z�=r��A��HA!���Hdɿ�����? �Ps��_ � �3��S��[�7-_;��2
4ns�"�[��:�	sJ��8 �15�U�>�iףO������/�*@�x�;�[s����'ч��5���n7�5j��P�PR��'(��▪��B4�IGTOԙ�5�W��K2{�db��;�0�PAj���Z _"�~�ć�LBV�X^c_�1�{q�f��#d+?��|6��F�Y��n��s�:��zB��3��ry��{��(H�x�CDa��'�7xXkQ��Ac)#��C��ت�A��`��,C��_���C��^�l5w)����)��N���O=�Mo��
�[`ֹ����烉4&��= ���$$0�
k��`)�s��ؗ��x��t�gw�o邾�9����g��z��㒟��6*�椪�]:g�m��H�P�<�
r��QKc��{@�Ղ}�f�����gO4;?|i6�w- eqф0!�����	�"*���>5�P�TK��k�d��"$�t�T^�rt8�T,���;�O M�2�1F�S]�>�x�z-�6^}���@�/wb𣔋8�j%��,��&�b_BkMwC�igj�aΒv�z{#xp�:05�]��&���*�4��J��^\�#ǎ�8�8��#����۳��
C�|��� �+	�=����0��a^�����+��ʾy��8[�MC%�yi�9��n:(��*�B�Q~����	z��t��F�6 ��?v@�è)�QQ�q��`+��;1Â�td]��5�u���`�_��&k���Cv�4�rg�6��V��b J��@&��+�H��~8�5|��+�zZ�ܧb�q����0�^�����͜=�/UR�vK)>�_�������-L��x����[��:zA�>!f��=��R�)(z������@n����"pؓ۹PZ ��+�ppu�ol4~_)�8�R���**7��
YR>{�3E�W��}�K��QR��q2-��2���Ѝ����6�ؕ)aV�1�\_�\۲�T/������R�%O������y�aC|��c��@O��T�\<2;k�_���%=���񐓫�;�49�N�ĸ�'0}����G��2�yo�̾7�n{�A=e�%5����fF?J���	����X��y{W9�V`8r���ix
7Ea�:2�h���r-3��]�+�'U0�!��N����`Ye
�P���B�F�Y���ow@��5L7̷��~t0��H�A��i]�;2<�D�:�crj'DbP0�� �x�OG�!��.�[�pgm�{NPi
Z������3m���6��� &�mB`��m-ڵS]��²s`�}�`A%T�O�pi���;����x�=>���?p�	���?M��W��x|�������0�*�/π���	��T�Y���E�[�4�]6�"O�k�R�U�ٓ��R��?�M�|�y����� "��ڬ-r"5��|�Sk��BsMw+?
z�a��J1��[žz�5F�f½�4�J.-?��72{뼋�k �`�p�
����ՀC(�b��ʹ@�I��w~�3��C�:/HDj�
�o"C��t��P�ё�����#iyTF�$�.�i�̣K��3Y"�<�P����q��!Sc�&�kp�J ���e��1YO�s�~��B̈\б/�w����̺����8@͗M�XS����3)+�f\dh ¨�X�Wݣ�il���T�Y��+��l�]��Cߍ���jJ�C�&��0������54N�3��`*�T�]��a9NH�*@����1���R������MQ�c�����Þ������f�og�l�,@o�]8����^5��1&B834�gw2S35��U=rr��/0�q�g�\�aW�z8aO��#ۭh�-�X�C)��iVS���!Ԙ��f�i�M}���~����l��=�N�/����2��6� @���:�����b)�{�-sEwS�3~���n=v�d2�y�K� �.���Y����:άZ�ϫY|�����3��^�8�i2�m�/�9:Ű��^�ei�rV%�A�i$O��`u�8x螘��h�b��3Y�૞7�7kE+"�&%;T��C ���Z��C�����_�:>��h3��-ݱ�P�P� �g�o��[�'R����򆋅���D��sn5���r�dzг��t�������U�xZv��Ģ�bD2nQ'b����D��^�(�u�����j��aC�Ȳi�M!i���hP�0�O�� �d��f|����@黲���ķ�t�;ÜYk1�[A+�$<d�Y��#n�LQ�X辽CKA-2�%�3龋����=��ak0���m���vѻ*��I*��E@��Ż=e��i�r�J�ŝ�+� ���(z�|((�8����X?��������y&V���{@��v:��'�r�Z��1S���AG���$
V�����r�[F����5Ax�z�t��L3UJ��3�`��v^g85���;���تk#[f�*��)'�ƃ�� �h���ԑ�>��-7������X2�$�6PӉ�P�AwZ��`���\�MU*��ϴ ���X<$STKsK�ͧOwu��p��0TM�s!u�K(��ٚ���؍����vQ�vϳ�Q_R#DC����@�&�o`�:�F�1���.����x����0̞�R��1�)s�u���Wk����L�yTj�a(wP*\���4�G��DŨae�W���c24߻`�g����1Q.��Z��g=˙ �_����ɰ�)�f~`r���L��6��@#ApО���E&�lG��(Q� X��m'�gz�s�d�\5K��(#��x/hX��W�u�l�:AW�v�>�FY��@��^a�~�gJ�-p�G��3�`��5�������q��5Q��(�F�燐�q��O��
�t��YE�y͎�(S�\~�U�`��Zj���C���c�;���GXǝ�ֶ�K�^2T��&���f"��Ŷ�hcMcM/y�%&4;���R��l�'�38Ew�DnWU��l�7�u_��<��;y���Օ�Z~��o����ݪT>��I�ƛk�sq�:??�͢�Rއ���[ԛ�7L��D�6����\��Q��|,�Q���U��gF�Yh��L*�R%p��ÇxTQ�ه�s.c=�D���>
�2&�.rE�a��_y���ø\7?���:��������}랾����`��R� ͎�E�+W�Ni�i,�	su'p���N�T�Eu��KK�_ܭ[�	�<��,��`��@�%��s2 2�Z�N��ki:-3�J�:D~%�!�h�#�&�N��R��m��ԏ�l�<]3^Z�ɕ�K>&�J,h=n5"چ�&�"
�XSFMI��K[��j{�p��{�A�`�������*��YZwg�X;n��(�����z/eQ�t��?����(��Ѧ�Z�Ma�0;q���S8MU.�}s�R�Iقr�P�#���ăD�~�̎D��KN��3��D�5B�>��|� �r$|�8��T�"õ�x�H��:�z9;m� ��y�ء�ǃ&��U&p�%���z��J?/��W�G3?�|@Jd�����D�rt��G6ݼ̛�Dfjv������pM�k�K�>����� b-��F.1��e.�m�@MNL�a��Ш�@Z�.�:�m���\���:�;�K蓰PA�=Ds(��U�f���޾�FJ�ޣ��v+��+�P����d�^\CT�#!"W([���i�j�[�K��.3��!Vm�x��V�t��A��G�R��0}��S�|�M*<�M!�R�=?�qn:�-PZ?ޥ;�-�)S�a����1vw��q�/CM�W�d(~A���V2��.�I�,o-�rqh�0�g�+ݯ�XR��A��Rsm��8��?^�#�*g�t?E� �Y�\3���3bSt�bbh���<$<8���At�7u�l��7�hcsgf@{��塹xz.����b��Lĵ2#��"����,��d�����������@�IONp��>@irj�h��@���3ңO�z�SK_�����ϳX�
�<n�������5Ɔ�x!�	CNõNܦvKcH��k&L�+ �W_3c��<л�ĥ��I���|�.�6�*8�Z�mE�E���G_����uʼ������B�)�� �����~���G(�v�b{��c�B�NG��A�/7�d�'��%�?�ǯ�$<�R��9ѭU�ţ��ي=":���ո�(�pp
�m�Ϲ�R�R����9<1�^;r/<�0Sm�	Y������	p�1k#eqEO`;h?�~����)D��0������9ʁ.�Ï�}��k!��wn����v\z����N��ٲ�O
}�P��d���0P�����S�'���	Ԧ�~�C��&� ��:
�Ġ1��" �k�)6����d%��qށ=I��X���/<|��mS���T��D��	ĥ���j���2�UYCN�o1��h��3��?5�ZaGm8�O�&��g����0�c�~3Z2�9/���g�+?���,������<�\��i��d�Y�Z5�*2�Nu஬ȶ`CE��A͂Fp�\R����WUn�s��ό/�|��`+�I:dn&���b�[:e43��-�vQc�D��N���9����s��_1����#ā� L�H��� �G�%�L��K[*z�\l�a��*-����ϰ��yPUe䜚^#:��8=^�^���خ̙#�*�c��6gv��g�޹"�A����c��B��%8uo�c�.��;�]t�����O�^Z�� �^�M���m�*��	��k$c�bџ�,��;� �8��fq�����Kp��c�����1�MW|Pހ�>��	��p�mUb���u{�M��'�u|��6:�қ�g��U1)��lO-2)��LC�ܺ�x.��MC�B���*'5���F�Ύ�����>H�kC�-����}η�#=�U����>�J�����|�T����E6Y���=��`L�o�m�Gq����e�M)˲�b.u�!�%ip�D�|�	A��m��9`t�{3ݞ�p��V��֐���f�ii*I×�����
�6���l���1�O�J*�0��r1�҇�1��WJG�O��R�j�Rx�_R�ų���Ӄq�>\�^����<P���q(0�p�0��le�D�\T[Ƽ�U3)KN��RB���f��d� �O���m�.��䔶�?� ����?k+sܣ )}��DƄ!�O�.|rɎfL����
�E�>��WmY��\�2fI�˃�Cd�Fv�Z�������ɫ�d�k��R(+�~�������W��^��fm�c�y��`�B%c��}"���hO�c�=��n�0^��KB?'�jK�x�h�6�|!A>�q��#����+J�b�R �s����[ȽVލ��U���#o�Jl�T2Ӣ� !j������&1
�|��tcۨgR1�̤�n�]�����j̦�G��m�[՗� ��X�Q��vI膋"`��ĵ�� դ�V�֋lZ�>!�Y��A/���R	�暊�S����xIUC�ݽ�-�������Dŕ߰�Z$�A]�4k�1=;;MO�m����9�d��6��a������N;�B4E��S}��c� U����O-?�����!�Ez�m�*�� ���?m��?g�*9�)͢�8�rm��1E�-{ �g˓}0A�\��|�rf&�����;R��9��$������0��|(:�}�;"�q4�	��ڥӎ*ebcfJ�庡���آ��p<��*l/���F�^�6	��{?h����*�p@;�B�$�Xh�w�㭓�E�,�g1�1e�'K�Z��.�)QX��Y����9�K�+�NGF�NP}+ g'	ES���
=�f7��h<��.����L<O��XS�)����_*E��	%�~�!�Oӷ�U�5�A���� *XbU-�^�����Q͞(l�������e�vj1�����$p�Z�%���n��)�f�7M�y6~��~�a$G��KPw�� 5�>�OEC-���ӷ��#�/�`���W��s�z�)b��W�4���v�_: $���$`��js�y�p�^&Źg��S����sb���G�h��g�.�ׅ�x��M����n	�aV0Yi������n'�z�;�� �|�\��jD�ȼ���]�����6棈�].�Ҭ�Q��E�8˔��k��߁��X$��������:��HpXEk��T���U��ĝ�P�(���w��&��Q$��%K^�lI�����.N�L�J���aL��-��T�>�|G[�#�?@��!AS9O����p�%Ӈ����V� ��O���$��9�2`�VE��;�S㉷��`�u5a��}w9�q5�f���Xϸ˽���u��D�\dr� P�wM�[�4q�m)�_B�{�,���_�|�8fC�@y�8�p��'�N��J�h�n�9�G�[��4�4}��/���>�钰߱��lV��50�w�m���m�U�I���Y��ȅ�'��z;O���I�Hk�4�|����lH�9O�i���[R�H��OF��QT�3})�2� �Z���;}��a�f��=J�\�=�+Hƛk)�Bݸ%�P+}*;�WA��TZ(����h��[�I�O]T&�h,V��h�'���u�W�2�9W,�ҏ�̙�L�X�6���A�F�S�>D18��~��6�'���0�Aj��d�C���-I�a�FU.�^��Ӂ&d�R��Yb������ns����o2A�Ax`>�Д�3,
�~{r� ,�����ftO��i�z^��i6��%��$U,��e<����6��I��AD3�Z�2g��jϻ`�3�Wj��n���k���:���l�N�����1t��@Нu|p��v@�	�#n �k;����_��n� ~��2̭���LB[%3k�Su5/�&y���v�����g����D����:�-��n-��T���O�fZ�^�'n�+.v��ź��x��dg>a��,��R�hC��Ȃ+�{��Z�/�'4?���X��Mzm?��S�0�xu�*�R)�_/Dd����8��MEh1e���w�yAN���p������[�~(�A���j�v۹eD��J+�r嘝Л��	&BG���mI-U�.�7S����g��`N��=Wi��z��2�3�WЇUdf�⬽ˌ=�5�Y�ۦA����j���X<�����G�Y�N�V��@��h��D?�fS���I�Y<t�zs��Qj|9�AӦ�$�'�O�-��7A۶��S����0uT�Sg�Y�d�;�F��2�w)���_@x�'y<��x��b�
��y�6e�5�ŀ �b��k��tC�~$S-�"��f��*/掤���W�H�c{fF{�`���t��?'H�~���ז�`�.��g$A ��M%���G��	���+
�묯Ţ�x���(��
o�ج��`v�7��
�=exC�w,]��-�њ��Pp��I�3�}�m�#����l���S�s�ŗ�ڙ���N�v���;�����:J�f��/	T����)�:iM�y�`Ʌz;{k~k�,�<ږ؇�?	���Y�/���}k�����r��^�+�>���D��w��4��)�d���ng��N<�zGS��)�Tǡ�.�����Sȋ���"�1ݼq��*���W�s��w$��CO�qX����cCԛ*7���ÜWK1��NP�G����3�wg�eC�t�
<��h�ƶ��yIdr�~�[b�����d��������%U�,Ym0C<-��m�a����7ô����(,]5����<�˳خK*c7�D=Q{�������4��hR�V�V�����ۨ�o
Nq�AW��HI=Л�����p11���|-�`1�b6�U馿������Y�3ޡ���Z����3�=�>*�yx%\�]ڸ���fɷʿix4�0z���,�v�PH1�����^䧰�jc������ V �_����NR�C��:��m���G�u��	�I��|�4䔉�D�W�9�fN��B�k��Â����Z%���qy�WS�.�AI���Χ0�`7q�BV�{8w��������2� ��u.�����&KtO��J��}x�(*.�"�t����B:�(#�O\��q�kI���@�DR8����W��[VJ��K}p6JF�י|>E ��9�q�{Kg�=S�2���q�2���B��%��v��`�â�3G������i�mX@����fI�E}$�D�	"���o7�*4U ���"&�b�������P�e&aT�R6Lk��g�Ff��7SNK��W7��r�=�R�N��m|&�](����U@|�U5;�0=�$�? ?9 R>N��r\��S����D����	QξY����J��:E���,NݲR?=��s��0�n����Y�;z�4љ���ӗCl���&a$��,j����&;��w�^@+���Ch�<g@VA��t�Ht`��>E2-I�{n��)�j�T/o��v���PÝ�P*�l,�/Ζ�p�
>L�x��	O��^v"��?_�ܢ��J6��|�-ҿfrl�M���.���ߌ1��w_`on�r�rx(�g��9ݩB�� ScRW��޴������3�tb8�Yz�8YO����kO6��-�9���uk�Qox_{Dcm�H�D�ㆬ~�M
��T���J��I����b��d�Fea\�tS�` | c�Չ�}��&3Wn�!��kY�v��	��.�Ͻ�G�B�����ƈN7Y7]LVe�?<)q
��?�?%�R�>��	D��c&�U�d�׉'ˁwu<��nVXk.7]^$���iD��,�
�CY�@	�E��D��Ty��AJ����}�`j��'6Y���EU���Bp�����c�ihuA۔h��V:�(��>��<׷�����Rh�/P��Ɉ�jx�,ص�wA$&T�>%.C����s�=!bʻ��w'@e��6$s��_�� =y���3�(���H��	�PU��*s�=W����A1��zlˣ��W�Y���U��s툺F`��#4[�8U���R�\�u����?NJ����� kν�x�O�U��7~���ڝ������r�.T
��|yT��G���EGy�����h��hA[�Ei�lR@����3~ ��]h�h���1�N�mڂ�):�%��u�r_�����B�4ˠ��L�j��'�9�n�0d��>7e��@F��F�,��F�@������j��Ar�I�(�,���'@V�k F�j�)c�:'"��+s#���4p�������Phq!������	G�o��`9�j����G^g�� �`�x-B�bw�Ib���>zάR$��zR���0S�6����Uf�Fy�j���s%��P׊=�b���N�6��%dI#t�o�Bn��s����Ч�IIP�/�=l�ٻC�O�Ҽ���m:�E#ؑ��n]�$�
b^�B��ASAZ/���qE�����:;>K�+2��q�ٮ�4�	d�a�A�۰��e���h��WH�B�X�D����[!A{;���.ș��K�c�	u�ꪦt� �-�̴�`'I�s���;W��k�D���!���.�c�/��N��L����>�+d����?M��L��.O�B�'L���=�f��s��J�r,�?V���І�x��%h��l�7Ւ�J�Y}�ys��Nfa)?L�Xs>5g��	izb������\�I�4��8ي@�ζ����%Q6Q�lןJ���J�_PuI��QʢD�p�cg� �ԯ����vֱ��������������L� �?�?����@���{�˱�쒞+�$�L����Kd����7Wy;����Ux=���+�r���wN�v�E6����s�a����Ek#4[g)���TQd����Y���@5
�+�r���;����9M{�p'3l,�ְR�����E� ̼���������icyֿ�z� 4P̙ �d�Q&�b�Z�%Z�]�]7����'���؂0BW#�D���j�ϳ1[Q�gS��y���v�b���uU$��jx�X=!p��-��G��#C���;4��sz/i�}�ER��p���
��UJ1�VԐ���£ճS��^�~�|+(�u���3�3_��<!k�8��E:[�):/U<��,�?�������ڨj0�	F����8��]=���:����/f-�R��kP�Z�.�jKL1|�bx��,w���n���n+���P��ԋ #�F�>� ���.���:�;~�HHCY�>�h0�S��)v&7��E��Wf�6f�v�6�'�DH"mhO���?������TM5� � f�XwA�xoNe�_G`,����̧�GJHo.>�#RS�sa>� f�[O��O���J�I���4�r��"�7�yJy��S^_��-C)��D�����ʵ.�Z �$#J��h~��Q�&
iN���1����	9)^7I8M�=�n��УB�Kߩ�}VI���6�ߡ��6ņ�+)��>�o?�õ��E�&EA7���>Ԧ�Ͱ`�,?��t���M�C�<'o���2gXWR*�4������V����&J��N�@��3I���m��a�7B���y��w~l��azW&Qd��C��7d�������N:���g�o�k�P��iN��k��f'Hun =0_SHb�Q�� Z��[N���&R1����[�[	�_������f2
�6���[�Q~��]P�]sH����JdrB��?�`X��1�ݕ;������G>�AʥZ9���S��
���R��u�Kø��)7�hx�Q�L�]��������v�(e�nFY�D�DW���`ff�G�Sb�}��crl��oc�%@� ��Wt��|�e���e�`*t|'r���M�w���zƀ^hё�p�8��c(z��=ȧ��p�5�0x�ڄ#�ں��«X�Љ�q��_�	�{s�ڷ���y��:J�JABD�!���+�z�>����	�d)�q0�ؐ��b�l�T�������uFWD!����Ok�t�Au���Md��h�Sg���[��v�� �h����uTn� ������U�D(��GL��Y��t�t��m����o�H5�������T2�s�W	3��Ձ9p�Z�$�F�f\H'@�4��y�������������������%wdz�ɐ���0��7M���4Ӄ�i`�-��9o@�Joc�z�W1��
rÂ�`{xgp�،���EG��ə"��rW�Ž{�goyE�_�w��|w�����5!OT� �#����#} ���w��1���4�Y{���r{oc[z�jD�> x��xl(�\9���k"m�n��&���w��n`k�l:��cCN��F|r���}��e�<��t]:���ur�ԫtc"Y��F��@U{K����[���ba�O]"cɚ'�݌�����L�M��O����v>C	����n��_��w�߿��|����~Km3��.����T�����Ic5B��!��xm�y��g���HU	�%y����ƉH�{ŵ�)RJ�&ˇ�7wA�&� *b�l��!B���E�"w����-�����)�%v�;@`K��>���5MӷS��Yi�}�6�L��:����{u<0R`������چ �^����L&��l�ܠ[X�Oޒ��t��ة���9^�OQ~5�Av��ؒ�?�=�m��H�Ղ� ��^��À��+���ܒ���o�3t<�j���4��}�@�,�Smp/\�ū�`���s¦g�d��όV�Ǌ!)�ɨ�;��-�U��,c��/P��_/h�b7���2��uz�m��O����r�G�L��
 h���Us#K�\(Jߒ&��ky��C�*D����F=B��!C.�	]���*Sot� �/����np	 �HǼY(�1�v5_��l�6hs"�C�y�dZ�)�hO� ,O����gt�3�y�\0ʐ��י�v;k��TV�7��ɨ�	�K	��i���E!2����a%K��>sT��`7F5m͖M�8�m�%+	;��3����"`�FकHT�}ɢ���}�c=�[0�(5�^�Q�v򐰈Tf�#� ;����C�҅X���R2�p� �
�]�����u E�{��0⽪��W�ϱ��S�&��Mh�u(�(3Z�jP5TL�����K�@�AQ�)J��丫�uf5y��c��sG�������gf(��a G�1G���`B�S�~}��6ߋ��[E�f1��ʂ���8���)@��@��+����y	��Ǉ!�e@*<�f⻗A���1���g�} u�:3�F�S(h���c���t:�
pA��ʨ7������� "�t���o�*��%	���g��}K^� �Р��Ew��թEZ�W��wZo���/Q�ݵ������jp$5MT�܃�:Cm]JNԞ]����H���LO��X�"~R_7�La��Vg���6����@��s�Q���56F��_�+c���H?�G���íp�8�w�k�x��ea)�d3�����g�<2|�b	xk>���!T��RDy<��+jM��sP*��c����imW��h,q����fgHpe0���$h�^K�{xI�
y"1��٨�lV�j��0��J���-�{j�._��X� �\t�X��G
����E�ӱ��h�͠�Q�t�<��j!a��-�㋚	G����-߿h�;D7~4���������b������͞=�����߲�iTv(�q����?��6л�L
�G��E��ּ��O�ӷk��N��H�9g�8���M�c���nUzƭ���ӵ�{Xp'�9R������&
L��$��`M-�А&�X���fM�L�����SR�~�L�䌄���&St����i晏t�L�=?o I`>a_5���-��;��;�E^ςx����X��eGm���(rMg5SY0ad5L����s���y�I`b�_�^�6�Z*�H����������_r�C�݊Ԣ�Ѹ86�<��2a�i�����(w,�2�v��?
�z�Y�ٍ��*�u�7x�S�j�P=��<&H�|̔綆E��0�*��B������l�e���v���_���Kv�y�[%zАn�8�-c�w%s>m|�Ow�<9�b��|�9�"�l�Y��{\��x���d)Ud;Z�mos�Ez�nW�;}C��aDw�(�$w��ǥv���%�7-�wKT�K������/g�I�N�*���OHJQ������0G�%���Z��d��OL�L+N8p�ÏG��}�2U6i3�h�2"��?���󛨺;��qb<���1�V��9�:
_�n��a㓢;�b/��*{�qV�JF��:?@���۵��*������(ڻA�y0GJ�}\��*�׬��Xdi���o~qn��a`ӟ���t�3�dE?���A=����8G�i�̧��"D�	>B]~�5��S�R�֠e3\���9\66�(=�}�aA�h�=��ujM�w�����w��E�R���w�+��{(n�H��g�9~Kxh���� �a�	$�`K��(��<���F!�CA�-8��P�"�cZ5��`c8�Xe�� ���?�
p`ӱD��9� ���[zƥT/y>X_��>�����O�z��z*�AS��ay�Y)U���t���׆!?���Z�cqM~7e�j����#ӳ���`pF���I�z8ea�0���dlC8Q]lVR_q�����tT�'�8�"�L���fW�>���(f�˾Yr=("w�-�qG�iG�e��%�^;̛v�~��������\��{����J���!w�6�O�Na̡Q�yX��d�������'�'5����1��ŷ��}�[��y�'9�h-�|���>Γ�^H��i�k�b��qz�T�6u��>d�c�́��}�^��'�K��F��t��vMX�}Q�7V�^0����^�|D�Ȥ���8��s�"��N4�VF	�� �4hlX�����Pl�Ƽ�bi�?��h��2G����!m�\�vW�y�V��Л���i;���GM�
�Yq�TMk4W�0I�鬨��Z��{�+q�5��G(�4^�(��,|�W���IϿ��UC���"m�:���@ ��fi2���ݽ�U:�In��cH&���@,�m�P����a& ��F�T�3��G�m0����M:N>�|�0�#�)�O�	Cx� 5����n��[[�(,�,�e��T�!zn�8�d �������cr����k�NÞ\�M,��a*��G�L�3���3��(�}�/X4w�T��ﵭ&`������?"�B'~X�����x��$�v����W�o�ѥH%�����)�O�P2��Z���3!zi��J��)����T����WH���y����[��H����)��Qt���6v¿]Ujѹנ��	ƫ�3�O�8\ �q��z��+�C��G񲥕i �uP.�:�tdV�1-�T`,���w��zz0���xa��A7�>��6:̨�̅��_�\EH5 �re�!�v��(�Vt�U]
Q��;�  �d��>�t����NC,H)�p�������������L9��!��c���|HPvB�& �#�ݸ�$a}����
�z&����z�|n�^d~cNlC���'zB�;���+��BJnsN�(���MhGgu�c�=�QYT4L<X�vm���)�67�q�j�{�gK��f2 �|�C�^?c�c(om��~q���2��k�0�&�
G���v�9���4�Ђ���_�ѹ�P����0Z�ze,L�~V12�e���l{0�Zr1O�q��n���}�����T"�VtH$:�$�6U�P]�cyE=��K717��f5�v���)��_T�!����2n�s$%}G��j��Ai�����st�"��Q���-�m���x��HAuj�l����g&�Uv���mU�d�Z����'[�k�1-��� ���Sy�>���Y�qbm"��e�N98Ԣ�4v�s��Gh�цeq\��w��P����7]r�u�`װ9�����5z^�1�gČ����+%��"V����yhꗢ½�3�|漐��$�I��I?8��T����鐱��g|�К4A,�4űN��D?�����*v'$�J�f&���e��N���LnE5 �Z��9ApK7"4)C`Wih��h;Sj���+I�0�XBM��M��R�m*R0����
Uk��i0qwSݷ::�Y�g߃tр���{��S3mL�-F��!��ܰ���Kt]��jtL��Sv5ߠ��Vg=f-�i�B���$�G]̻ӥIJOt:;�x�s�?���� Y���N�a��E9$l��ŝ��M�����MKZ��b��j�:�����q��}=0(g�s$2{�O�9�p*O�7���� Z�Vভ��n�M1�,^�����E$Wr��7��6i�f��b�N{�I�t��Ӿ�E�M�v��~��9�oj=�XX�8U�M�-�j�Y.�Yގ1V@h���b����*=r�V�W�N(��h̢D"J��
����;����I�������;�G��=�-���%+p��*��|#q�A/07�&a��9���4��/Z��^K��V��i��ȭh��9�ȕC�ς��Ic�!e��� ���/z5��N�\��A��>a*-.�Q�G?=���{ �֯>b��@s��SOX]:7�
}gyw�U@m9��r�{�r�o�c������F+�����kFi����5�U��|uS��[����LMcY�H��G�aKp׳QB(n�hf[��ɜ����$MjX4�~5Q��yA�\M4�:5����(�W��z�"�;`�Z���,�:��^���:\щ-�X7o�� ��D���Z����(aΛ�So��nd��d��g�����9jA�M"Z\�7Wή�C,���/<ј�V�E�.|z����]X����v�Z�0��#���J�2{+����SUo�3Z��.��1؜�kʮ[t佾j����#�3�SEhI��F���F=�0����<�<֜�.D)���L��\�%��J���A��~�(�_p9�A46}<E�Ç��6�	��5vq�klO��)ޝ���*������K r;s��AoN�(ٷ�>\�<����Y���v0q[i!4�n��	�`;v<sj�wWb���p|eR9������_ݻ�:C��jSuTNz4����!�?8��}^�\k��
\��-�f0�G FVL�:7 쯃WX�YW۟(����Է�jƙ�Pc?A\�/�E��.ޥ���e�J��A�ʫpɏ���)�\��t�;���@kc��Qd3E�î�I��^4�^�r���*��i6]��� �}w`��s�ٕ��o��SzP�`��9���`�T9���A_��Qe�C���u6�ɀN�Ζ,��Q:<g��W�
Z�(e���BM1Eжg����0���͏�P�����F8�����'�F�&���U��wd��S��T�5�2��B�F?4K��n�����|*ˊ֮ܨ�2ۻq,�/.�����<#�r�8���t]�b}Tk������.�q�� ~��W���&���C4ն+O�X���tm���Ƚ�5%T�3?�jȦG����g;�F�Z�7���-�������.���X��2�<L�dYNzG}�Y�L�(~ݼ���H.#O�Ȟ[�m� k���SL���.6�(�k�՛���x�����an���<6�,��3K��b�����z�H(d	ɃH��@��T0�~���"{'�U��q���3O���ֱw8�dA��ۮ�Y)��k��^�˹�ax�@����� ��y��|��9��!G����VJbu�{C�Q�7�Z����{bC˱]��$�x��8aP�'H���.�z/�A�|��A�K�`�(C�H�A��Œ����J�/%�'J�ӟ1��Tq���Q�o�n-�p�\�u�X��w��]y�&��g���$G&B�3����d������}*��ā�Ч1�PkB���9�W�1�әEu�/So�G1�fS�ke���_�˃VS2�;��q�6�G�F�)݇'K�I�]אR?����� �&�xl&����9�=���1�����qI 	D	})�6Z*��Xl�<K�t�'�Lqu(�� �# �%��.�A<�=�0%��]w�I�'v�1[�U~B� ���Dt/5(�m�[qA�j|Bƒm����ǳyZ��@SǭН��o.��y�>����Yn};f��i�W4V7b��_��2�w��ؐG�O����9�L�4y_:�i�:�diay[N"�ZZiCD��뉛� e���O��yq����%�܁��d$����ɭ.�p*��jB!�Q�`��<��{��̖�tn��w�sv]�b߃K�1���}<%�oǷ��������Ϲ��<[k� �4��K�bZ����BF4�a@�����~N��UCmW���S-�5#�eY�� W�-G��fܱ7ʤ'�1z��fy(���@b����==���?:�v�؀����y�f�����/�64��tZQ7��seM�������g��uE2��/��6� ���'mk��)!��x9+�<�庲L��v�`O�Q���`ޙF`�����Jh��y��t����.(D�3P6��[y���:ԪTG����/�=Q�O�g�D�[��`h��GI�G\E���O:*�O�8+��`�?�sc�gok�>'A�8��H�%B�ȭhI� ����[��b!^�{b��_�P����>�h�n���K�SM�����1ɖ�׻C�����0��N�N�Lu�V� V>�^��Ģ�Qu<�����;$��ʸ�z�#��MUk�J^P���8IZ�K�,-fɄ��e6���M���^��F�;��@5�x\8��3����{!&��	E�(�z!ŮXxKyl�|i|��?�K)�+�c�ٞ/y���0m����c}姸�|1���x��g�������͌c�5��c����%/������1��˸q��!��}ٺȖ?9#���yU�*�~�o���T�"z�_r��"��jPNoλ���A�J���J�?u�C���j�]�~bX�%���Z��3���y���%�sgRH'~����͉���o�������Lg`mN��x�0$��t�
PvטB���D�����1�\d�0����"�r%X������_j�9,F�������j���d��n[4J�7Dz?���Z).�)�{+����� �j�S,��P����VrH�Q��N4-X#��5	���س�"l�:ѫ�xɰI�D���^y�`�@<j �3�d��)N�n��]Ah5U�\��I��"(��(��UdtI)��&�!��Ĺ�笠�9A¨EɐY�Φg3�j,1��M���i�>!d�:9�<��U��^NLΛ���w�y��FX�xt]�vB�}7��B��_y�Cޗx��%#��y\ȉ>}/j���yIr��+��$x(��=��1�b�YpZi�Us)��CvH4P��Y!�2�g�Y������I:`��Q�y�b8��<k7�c �l��v�
8t��=	�h�3�*[|5�(5_�:���P�ԏ�{*��ó~�` �� b���F�k�[JX���w���1h�G'��Piq��W��k?yz��oޕG������@��i�cG��q���<����:�=-\�삽�<H(c?���������ir�+P���,0��*/C�̗��W���	�S�;IVqYm��贄�b���JKV1�:U�k�s �"׫���V�8"��آH���OE+j_�r�}�x�K[�#�J�Qu�L
r/�ĕ�Y/>���:A����*$�͡d�&s���T�/(���~&��ޫ֬��e+��༕��'N�a�|���j�e̤#m��`i�Fu\j=�}|�a��T�A2	�i�D��OG ض�k@���y߉�L:�S�~�x�-k�!y�Y�1n���=3X����K�x1�Ԅ�:�W�Ne"rkV�6R�3äb��M�E��$�C��͢���O��:���6^3�{�^z'j������Opp`�f�����T���X�a>�B����百L�;����j.��xӠF�89Lb�{}����� ���O��|<�g�����#���,h�����~5r�����'�~_�ж�;���[�<h*1�ny����_�B"��.¿�>Ȁ��A�:lV��0�e��X�<�-j���ף����ms�4�8�X��0(!���9"42B�K���Yl��(b}?J��������Y�\��M����-���9�?���Օb��h4~�⌮2.�2���&A�b(��+�e��b[Hہ����!��.b�9ёX�a,�����G����1�����c�񁹆ڻ
���YJ�Q�<:8���\�vx7�@abѥ�؆�[�`+!XM)ٚ������Q{t��5���*�F��;�
����PY���v��L����ξ=3�V/L5 n��$��e�XU�ui� ����9.G���}.
-c�#$C�f���VDv���l��gH���	�ǫ��E�	�j�6<J5�8af��j�_�U�AL�g�6�J�u>���/G�Q�+���~�@#��rB���H��Ir}F�[�t���T�D���)*��9�35�7��tTT��8�&�5�1,$�|���J�eՌ������+�dav'�^��O,9�+���?A!aK4P6�s�gR�^���_̶�4%��8��?:k�_�;����5N�Z^$�t������!�~����YWr</d��\��Ե�9��k�?��~����U��3������g����8<�5�2����0���i<��Ԫ����K��L*bb��*���Uˌ�]�?��a�1���^��<�(�2Y��V�)�Z�Y��n��5ڞ��"A;�=�ȹ��nYo���Dx�I��\�]86P:}OB�ˠ ��ɟ�+�1!L1���Ѝ��W[�l�����QK9V��{V�?�z��]u�5��F���c�1��64Q�s�m�M���j3�k1^�����Z�bC�.3Ԥ2\`�^bh1��N~�X�ɛ��^ �㬒U~����=�S@���Z>�
-��p/u�{�gy@yW�7 ��'��0jk�qɔ��U���3KxE�$�1N����4v�}��);�� ���D����q�6��:0!�Q� %9n$9��6։����)�:�?�yy�V���e5�ēɨ��w�v��&���O���Q����z lU��(�����(��g
B�mE�
YH��7X�yn��WX(b�t��꠫A�jǻ#�s,cy�5i������`���Ihg� �C��q���O�\�z>1/
�Dh�E��U�����o#@MC���M��<���ތC�@liwyl�T�uB�is3L��H���j!�������ҧ�4-Hm&"�H�v_��n�閊؄�e�Z�r�_��˃(k����O �;�Y�]M���yC�i����}�h�8b�
���J�LwM��g�_�]�����"la����"u��#�����p��"|��Z� X�C�T���WK{����^p�D����@��a�1��T9���F$�b��H�PgJ�;*D�?}�̩`E]�b��B�a0<��{��Ѡ��(_��ǫ�@����E����;\���9���'6�[lm���9�J-AX�.�h��ଳ�=4���(��`���>�Dߍ�q7~�ñ��v%��[��*���ʱg��������4�.�X�ՈA��̃�N;��C�����D-�h �����㑯}�ʝas�+Q����1@��ԉ���S�$n?E.>�Y,"'�ڡ�%�r����	SPn��8�$]ZX�a^�����<�B���.PU/=6c�8]W���\۾l��@=�AgN�� �9D�jn3s�`�=������������D�~�q��;
m��랜�t��Y2moE��x~��q"Yר�g��[�T��}1͕��o�o�w� A`N�鈶�w↻��j c�:a0C>�K�`� �`+�kyC�y� "w����v�3�U~Sc����^A]�I���P�~���1m�9̊��1NT 3Z�RK(l�.~�w����8�̧����'�j�)
+�z���I���^�۰6��)�����<�(����R��哗Ӱ�����T�.���Aw���x(�LA!ޕr��z���?����2HG� �j���uIU�ͬ�F-��S�V��Ŷ�ģ�*{��
{�xά�eT�+Pŋ�U����,��K u�v�	���S��	RK��jF�z=c�/n8�n�
ѩF�1[�{�f��J�9�b�אpt�*������$��Oc%�1�ڕƤ{)A<�ƅ���Z�@��ߐ�\���@�����'�1�v�P/�u�����"i���O������
�
�G�{��V�J#� �q 9�.��,X�7�6�ܔ���MutO�<�~��I~<U<x�ƛ���0��C;l��	_�3=S�4��T��Gaa^��8��=;�� �D2E!d)��՛�Y�y�Zo���o"�n�yS�7��('߼X��b�� �Q���,_�mE_
J�hσ�@9 �+AY	�^�h� ����hz	�k;%����C�J�����Ž& NhX��/��Y�Vq��dd�n��2�w���V��: ~P�s�@��d�xɝH\�!s!����}����x	�;�"J��"�5��#V�n
C�/Ls���JPD��,{��=�
�,��;=q�E����}�T�fcF�l0끅�o0C��u���\P�
��ҽ�"d�e��7J���T�$�w�ɠz�6�=��j�A�/��ϖ�YMZC�M2d�d���x�C:�k��֝l�)�oש��!��1u�$)x7ߏ4��p�PPjM-b���}K6+�ڹ�+�<a%�$9V;��
�G�x�Z��ig����\H����������5��MW���B�W�
�P���]sf\�S�_~P^���e�����`&��\�$q�Sl�V������I������_��U_����RӼ�/eF��v\��L�K"�rA�.z>���;��+�2V���
����]�JI�����)�8�;_gh5�+jsR)�>�ㅈ'�si���r��VYS\�v:��Ww�l�s%������(�z�	��;���I�eY����6O�_��I>Zk�I�^re���y�`^�Y��XZ�z�Wia(��wl��#�n�a��\+����W;�w����`9��Y�(N7h��:*�hsA[#�h�}�*��͊����x@[��$ŠG5Ӹd?t1�1ă':]�T�=/���"u�~����~������@i��>_�2q��<��z��dD��G�|"r?��ɪ@T�b����p��P���{Zɞ��VW�7�	���)�`�����]}G1��B�H����Ky��V�Q�k�o��QQ<�����l��������]��F֖�	��:���Y��)vyp�,�ݢl��r�k;�����Ydk���Ӎ*�^��>�Q�J��{�Y*�w9U�~��y�m�H
��q����������a�®>�,?U�8�y/�ב­�B���v�[�O�� ��|E�E9��*tg���N4��n[_j���Ma.�.>%�l4z۬w�y�U�b���@�d�&��dR��V��/M�h�����X�΁Yf��$�(æ�C݌����{����ܔ=:�}!�䉷r@C�aP_]OOop�ؙنn�8�ׁ�NEx.���=�ț��'T�*�`��^P�g�s�������:S�JT_?s���ߓ",���DP� �.y'�r�]�]��Z�W6��G%ܘ���F�?��Lwʮt"$bIpd�/�l����~Uz�#�n����Tn�q�(�T<Aw��Կ�v~�LQ&��SY��e�t�	�������^��V4����d>�h]�jH�j�#�d8̗��@
=���������Ga�k��O˂�EH�M�*l_nXm�S���=�8M�%��6����NH�����}�$8�d��1wӉe�N.�V���������l��siEd+,b-ߒ�׃�0�\)�/g`������纑~����3����E$$��R'�T3��ք���eh�� �� �Ś����3�0q������;�hu��& ��/�9���W�\-���ڷ�?��w�����<�c�w������S���<��y_݈�X] �v�*�	���w���nC��SR\��Ї`��1��|�}m�'�]-�iG�z_��lb�O�����d#��r���L�s8|��<3u ?��'Ǣ��U��U�QsPcs�r:��~ߖ�F��ꢃ���v8ro�b�]���	ǀ�SQL���S�H����)3��4bΏU�y�t���ZB���;q��b����vF����I��b�YaT
����:�� ���
Ծ�@~a�F$�N�#bt�.���į�94?F�����4}�{?|���
��kB��"|�2�D{~����t�q�+Φ�x�����w���<#�wT��@c���A����]-�����p=�a!�RGXi���̗� �)� ���!�2H{^��:T�D�s$���Xx�J��Ti]��B�P/7$�m�Bn�.^��X�����"E��T�jOX��n$� �;�p�Y�do��P5@�_�1Ȝ\�Y�һߊ{���6�_K�˦j�����o_
�(�A}�?�����wI�����rĺj3 ����vK5����5Hl�^o#^�v�+�IZ��x�,2`=��wZΦq���-��#֠6p��!뒂��-�㩗<����H&� bH��d '��mv�N�^�#Ey��l���V����B�ao�;�e~�Ń�v���WG������q\稡/���iB�;s�uD}�獐�C�Ҥ����nI_���4���8���	�F��3��e�����*K<z����Q[R}D��1�e��CG�:\�rB��vq��}Hc����}���A$��s�u��@8�i���G�o�AG�1�]�5�e�&��G����,2�B��|N�|1�ϻ'�{R��-�4�Mq�yC�AI&�z(Hp:gd�(�p�b��J�J�˙��W����n�&Ԧ��	�{L�=R��f�8�qrl_�Dʓ�%��0���}�б��LS"���>���S9I�E�5��k��v�T������� Khm�R�e$饱.Q4��P��nS'��p6�q�	O^�f_5v֖�d?ƄOR� �Wڲ|�J�;.4ꐲ�o�چї��]�&~�r����t�2��[v��� �CCL���0K��Nef�Ǚ����L�ԭ�j.Q�:�'@�g���2�l��m�6�m}+�/� :�����~�*8����A�$�E�_�ܴ;�wQ|U�%aVbX�jWP;Q���ۅ��B���fO�R�,pGy�q�r8z�,=��L�ǻ�6�'���9�����e{�!���q`�5W'=����&��$�(��3�ޕ*k����l|��e��U�QT�!��!�F{�ؚ�p�#@ѶkoDq�1�� \�#T0�CY[gx5Y�܃���FmԎ�p�b������ �V�ݼ�\�͙p5��%��G�˰�#ոm_���p���p�Ec��ow����o���ڿ\��&�^g3(�?F��Qu܊:�tD5|_j��z)��S<��l�`4~4����,���ʅjwo�n�($NULUq�]�6w���lYn⾼;�����w�i�&@�{�l����|�+�gǩ6�V����a�����Q�f�P ��s�]��~ڝ^5H%D8��]
/���hK�1s�uO�/N8v!"(B~��3�_�y����q5<�{ӊp�a'��+�`�j&6�'\F�-8�h!�A�Zt	ZL}�P\<��?"��r�SuD�a�Kz{�H����%��Xm�/��bk*	R����{�0D^�����+8v����(ʳ�KI?+ϑU`��; a�%f)�26�{�ї��}��˹~?���
����X�����t�6�%�8y�'����8:H[q��N�ҏuy�(3Qk�UΛr����3����ƭ��]��CPaO�̿��?~�4�7��}�bY��e�zT�M{M��K�`�����P6�6�$S��bZ�*FxQ�h#B��F�t�ag62&�〵�w���K��9��9%�c,���)KS�m��Q���oj���T�5�j3�ˠs�
����p���pig6�bɍ./��VJg!�L	��W�o2���֕��n�|��X�Hx�y@��6��0,��<�r:y��D?�b��Vb�ۑ��Ў��@�����<)���xL
l?Nƻ�pܭ�C���0�sd{�Τ$�S�Ή���F�q�5��uW?�a�1�=��e�5����?;r*P�6���sA��ӷ���<���i 
��NĬw�Ԥ�c5;�E8Lo�"����g���P��k��&{::J � ��v�ְ���C�?��)��'y���+�R������� ����Дa�%���Pڗ����vYN��N=Ce�ܡќ`���=�i��-$���*�ݩ����6��N��QݐtT'�o�w�hQ�{r
��M"�(p�{������מ8�3�{��ߖ��&}�?ensZT^��c�V��8.='�>(:.+<����`n�8Lʹx�������������������*�叨�~�����xu�כ^+�ʬ��9�Z��V-H��j���|-���D�}�,�����x����#�S��3�K[*6�����R�b'��z���o[$� 邈{�v��u/K�u�-C�aew���LSģ����h#ֈ?Z������!�ގY*I/�3'�Y���F��}z#�jC�^��-A�S������5>׿d�q�\�$�u��H��o��Jy�lKL��^p��GkI8d8$9��$�d7��B�*u��w%�e��qf��c�G�"��:��7��Լ��꧉���sl:'/���D[���'���ԾNS���b�VA*�hfqV�f�'��n���؃/V�#�L�k?N�|��W2�X����'�Vб�"Ѐ���{}��E��*�������'���L�y��"[!�>�/������B�[�y�F\|�7��ҩ�j�W�8�U�L�B$'��
�t���<�����dD1��2�|�������t����%�Fze��	��G=��ҩ'�h���J�WG��UB	��K�g�GS�MJ�����nƽ$��Ƈo�ڦ����G��l]�g�ܫ��j�7�5/�8Lx ��]ewdj��w�z@���A��뫹��j��=�ͬI����yl�Cpy��"�q���d�k����@�}��/��~�U�A���[�?���n��V��l�ږ2��]�\��֟6��p�:���zԳԽa^u'�Z/y8)�op����#�������;܃B�Sצ����# �a���o`��ss
�!��q����Y���2"�jdړ�����s�)��O)��ޭ/%S��u��lGв�N��R�[?hl�E1��W�/�����7����KXUu��h���NY[hQ��Pb:	��)jZXื�1��h���D����n6��x���;X��|J�{I��l,����7�m�l�P���ڒ�HRڷ���{<�c���-��l�������C������Y/��ikE�g}���2йY 
�VE���.D'���!�^�1(�Y�Y�~U��ʠ�R��s��c���>�Q��ɻm7�Su 5G�,��	@)<�5f������"��t�M���ʒ�YN�b�qf�+�#b�P��G�T��.�Y�Χ�v�t��6��S����4Q��W��=�����Æ��nJ=ʋۄ���\;$M7���:��}�N�M0��=����E�`�%��O�N,x�ۄ�- ����v]��Q�[ {#ݍ��H���d�r:$�޴��Q�x��Ea$6�b��Gd�����J$�"E)�t� 7��|�Ƅm���� �۫WϰB��[ Io��^��+>�C�Ӓ"rJ��GO�s)�&>����A�6"I�ǁ�]�q�B��)�F�7Ѿ����}����<w�
������Yq�i�i��%��tt�*��k���jl���k�?�{�?�5FL�.AuF�*��k����Wb��q�V���q�#<r��ƃO[	ʕ�����	�AvEyN�N]������H�9"���\���k��%��rA�����#T��_��vae�)��n������V-�8L��cL`/)<�F�[����d�
��.Wާkp���υJY]W��t�������H�9�`���!jo3�ahH���R��Ǚ��t������ً�r�?Ef�96��b(�{� �0�v��q����}���;�냧��e���P �9�"���/��CYi�s���m�^���ʗHC?L�枦[����,.(���0�ix־�0Kj�Y���vaڽ���=]wÑ�tp����?�A��$�0���;{��*� �b��1��7ݧ̬e3H��_I�:�%�u�g��Z��BY@��la���!����.��*(�z�"���qڡ�A@S ׳E5_^o���+��f��Ȁr����|�]�b���]_˫�i��+��`��d��#����Zsď$�@gDݏ3��?~�(��V��=�_�UAP��<�Ȗ�
����R�8:]1�e��| s��,�Iu?e�@;��x0���q���-�ޥ��4f�]i�4@̮���P�&�,o1Aj��V�4��W�g�Ea��#��l�$#�ws6�/��h�N���!5)t��#νd'����+�M
��(~���3�'�4�x,l�R�h��E7Y��@���pv�ߥnN�xT��D�����D�*���j�-����ڵ<�@v��B��2��K3�T"x���cz��s����A8ǥ�v+������o����&Snک	�Kzl�bJokIj�t�I��j]\�8�E�ژ�N2��D�}�ٺ�装a��沥��z5�V��t���x���	���}Ǆ� x׶d~�~�9�����1�>s�:��@ȍu�"B��ܗ5��bQ7�|�C��f�V����<�UX�k=��G�n5>�J�Cc]��"��R�P��;gM�������UY�AA�b"D���G��C�w����dJ�g����nnl��,2����!H*A!��\ l 	�$S}^��Y��l�)KZN�4@����/���6�Ѽ�����£GG����Hm]��[R������!�z��R{4����Ӄ�퍌q��B�h��s�H����d�`Z*�?�n���P���_V)^���	�4��鎀Q�+ͮWШ���rk}����\�&�w�\kZM���:L���G��G�n��Zo!&��<��� ��=��J?gr^��yí��9Qh����icEg2�	X:c�C�|/6�ːM�a�@?S�u��Lb/_C��,�q�4��ͩmJ��˿�;,��ъ�K��y+��6�ѻ3T��A^��g՛A�VX���Kv�J���"���X�V�m����{K�`7�+t�y �Lc�	 �~�� �dC0Eṷ�z*!9]��k�E�\��
LU�ֺad���ƃ	�ɪ�Hݨ��P�BJ�Qf�{i��/u��"��3�C�&Lcs��@|ڤ�.["���|��4�T�?�����$���[6V֪P�~1/�O�����8�v�I�#mԺA.@w?�c�&*���
?8r�@�����ȫ�m��I�-��(Q�� :��OY��W`��D�߳T�g	������dE�YD�fzE���l��* ��F�wyT���ٕ��?�E��ں�U�>�}\Q����s�� �Ș���s���`ꅇ��(T9�1���S�ʃ@7�f:�w:���P����:ݩ�&���m�R̈́4�m��K�/�[���:S��B7�����.�-�TY�����8���Py/A=65���iٱ�R�7�$���@A�SY1�#}�]t�R3^~P���g^q�ӵ[��P��9���iY�E���iU��Xz�f��-خ��]ց9g�dx�7v��<nw�ʈ�1�K��B�;�l"�wdo��@Jￋ�� ������k��K�VmטE,�[�Y��c�&;���I2��������ze��f%��C�sm�Jf�n~�d�3���m^s��X���g�\ ��w�}�����|��L���ֲ�|���%d���^ ������<|J�]oR��R4큆��+/nP�������X6p��ג�<���DAy�)�F)��(po��:跙�b�M4T������ƫW�ƚ������lRHf�d.v|��N��mk��Paʧ�6��+���$��=IX��n�G��,0ȓ���e���w�՝��=�	��Эg��`�}h���G�L�
�z3ԑ�����0�
��0Hi>��Dv-!�j�-,Z.*�E�ԄM��+��q�$������c*��YK���%<���*�E���z�٢r�[@J�?q���]��F��bq����7��
 ��$K
���tt�gңů/���AYu7�	#����P(�p����)ۂbQ�h�{s��}�^�9�9�
�%���k���ia<!)Jۃc�U�����z���F�U?P�ܣǪ����<߱�_hlv�k�ӣ�ۏン�m�ȘΘڼ�8�m��x��]�}r=;ʠ�:�cǇ�͐Q���b�^������Qy�����Pbm��{�L@a�˺���'�}��O#�"�ir�{�LB쟗p�ё��7c����wڒ4"t�Ћ���|L��5�A��~嚯����6�P�q��>M��4Y��$���s����+;�bf[4k=^�Y�!�؝��V3c��V-U�f�^��K��o[$Z�_ip_(%�<�@ݡ��\MbэR0� �Qm3aVh�4�x�Cp��~H ��F?*
qI��*K�;��M��Ʊg�J�Cx��2��;�߹��Sg��7��ȳ�������Nna��w�4����I�eJ����x���%�,����� W%^7�L4��mZ���`��G8O�7�&�,�{��H���Sf���5�ph�j��WX*��)��O(�����V��R�e��`�T��j����91K�A<毮���b��F;��;��)zx�	:T�5	�.�
����O�@�+���잽�E ��r3�B���g��E�k���n�3?'�J�)�Nv�@�A.R*&�e�R$�"���� Ǫ�J,�Qk��I�$��e��`�ʻ���j�/��%_O����gB`�DH���X��D齱�	(�%z�SC��J"��Nk������G/����3��trY�A�,�6���p]�޺���i�Ű��N߅��v�Z����(ld����Bh�?H,���ѴI@������W�,e�ɩDM��c@�����T�R�%��|�Z�v���ia�-m˓?Ȼ���
�$�	�^��$�Voݞ���Yl�����G����P��F�Mf�8��F�:!yj�b�Q�Y���V������! ���z��1��I�����7�	��)s�.r$�g+�\��7�ە�V�E.@s� ���C?� pGqH�J��K��,>��&� ۔ֆ�]��B���~��b�E*"��L&�.z)]S����<��|���>ZTh
�Vʃ�ur�Ѩ��� �o�vΝ�ɎC�^�?c��)-���ME�֫ﺐ7�'	h�{:*YF���,���\��Ȧ����f{c�Wt35-" G�4q�ЉX�z���h��)u۟�B�,;�1=�fd�N_��� �>*��x5q�D1��v�Ȥ�r3�'�qRP��ql�g(*v���� �Ѹ�����;ذ��=�<����棹��%�z`&I�t��JO.Y�&��r��\�O^eiS���#ϷGz��^g�3�G,m�@���d&B3��Km����kzx��o��
�&�������^���f"�����:�h�1��P���j�{���Z�m�+�j��D979�8�?|�!����ÿ��i� �3�0OU��?�\�2u��8�m���Ra��a�8�r����d�劄9k��-�H���*v����Y"�dt��븯�yS�#��� I�3kD��q ���^h`��="(�UG�m4G�u"ȑb�Е��L65o~��}��D�0�2*W>�U�m	ʀ��)(G�����q�R��|,�g`z��^�����w2ɹ[�1�$�j�Z٦�vsRNbQ*��|wc��D�<蚢B��������e���5�4s
/��M)z��u��V�灰פ�@c6�b��4�F��Z *g`+������n�����I`���%!��~�(�j�8�ܯ�,eU��c��'���`dsX��V:p��n�p^[:=#�0��^ѝ][�~��d)�g�c��L�"%ݾ����Gh&3$���Z�E{��c�������eߪq�d3j^"��7���i
-3f��e>��>�����:��1v0��yv�hO���(y�~�%�]A�g>�&�t�y�Fq=�bo���O������*�����ƾ���Y-]*�����-���w�����el���H4�-dGK�qO�z�&�1�F��mz����8M
w�� �/]��/�ˋ�DP����*���Oy< &~��.�ϓ�1�%��	��v��k		�O��IT��} m'��4�4�{5ZDD�����DZ��S����_�:�H������	�(�Ӊyc�"� ь��T��%�M8��W���C6A?9�4�n��!%��]V.d�,7��A�u�~�	!���������^ww^C��Z��gYO0�YxP�8�n=�Q�*5(|�#Q��W���<�w������3�!}O?�
�+��l[�57��z���$���2�ϋ��!/�,$h���+�ltJ��E��:��jfe��ڪ����uᙖO�,�+/�	�x��Z��l\ŵͯ�o�n�]����O��G�'�� -%�֤t�wWe���#m�cw��Y���Ͼ.�/#�Q+��.?^;u�LƷ���Hِ� ��|��b�c�&�� Ϲ���AbaȖkE�I�$��֊l>�g�'S�rP[F��P���!�+0�7#��?��(�@�}l�L��,(�j�i��AOo:��l��d?{�\���d�+��/��t>�J:H{�:�2��ꯨ�s�(`�\y׼ ��mC�"�-6��.)����o"?Y����>)�	Яz�}_��֒Q�K����La����k���jU���Z�yT0��ҫ4>}�}#�����%�� ���ܝ�_1��nR\�?�q�&��D�$?$7:�����R]'k5��}�n�N�)�;�YT�a�G��;EB���Kv�u�W�e�U���b���0�����#`��9y��y�3J�T� ���D:h9��V��a]�����FRz�B�
�z��2�f��B�GĹ���5�u�^�ka�����ۘ>�Ԣv��u�/�����"`2^��&Ϩ?6�1���7R��Y��&]w����0��0��Z�2�!"�6�<�1�P��;�u�OeS��,����N y��rD�š�,4W��w��6��-��J<�gZ���Ā_
�N
m��0)��Rk�e)��$��czw(o����H�o\ �e�a�m@���v���Y��T�Cj����9Di��렻Q`m�x�� �R��F���<�=����S���݉����!A�K"¯�1Y���J������m��}Պa}�����B�P�C���=��J}~�9���S׌"�Fc�n4��,��%�1���^C!��������æ%;s�Ah��1�y�����̙������Ӫ|MY,�to�)�2w���0\���j7<�:M|�w��e5A�s�#������<h Vc�,�^W�I�xZ�[ ��~?+^Q+0�q[�B�>�k#���}&75�ͭ��L�M�����*�=�w�:����f��0CE�"�78���#X��م���`�6�D[��<�Z��ب��,�Ҵ�%�-0z���Ԣ="��0�� ��w��>����z&.T[�JC��Rd_�v��=]�[�\3bbd,���b]�4�O�e��!^D�2��`U�a���D����1��NGe�y�娭NLԑ��$��D�~�.��K��0���F�E\�tH�s��-%�`�N����nӬ?DN��l�/�,m�%��>`����*��C�e�TC�	B��� ����3}}cV��bI�o�7}�m>�'�vK�si�Y^G��=_�&6��Kw	�ÒO����"����g�[�����ޱ=�[���+�{���o�~Z|��w����@o����� �?/.XCP(�:)BS��L5�ma�6�`�(��\��?��2.����g��sL��#}���j���	(V�frJ^�`<��"�g!���82b��]ve
Z	J�E(Y�Z-�s��V�3���_�4��g�]���5Mq������Ͷr̃���#_SD�����	s��!R�w=L?�9-�4��RVc~j�f"�*{�u�n��_	���AjW�"!l�nEx<A���z;�:֘S[�9��GXU�FD����_~e�򲿣R<���^�T��5�7h��Jp����%|ً]�7�|�\�B�p��9i{�3Pq[�G6gҰ:5n��^�>��/�b�n{H 	�-(=V�)�MR� 0����S�E��q�8mC��6�S�g��$t�E�U�u�*�R�j���޿|�}Bݔ�U4'U��8?H��'q�v; ��ӣa.Q�΃0����w�
E�3�b�y�DޔK���f_�
��q�\�2�JM��z�C�|�@v[�$b�S�d��ښ��Aңvf2�9r��	O.��G�/�T�:���H��L�!8]���=�t���Ct��}T���f� @�ն�P̚G�&t.,�dC�jv�S����]o���)�}�Iٽ%ݟ��i�V���5��0�.a��7����8^��l Pӯ�evfgJ�5�s1����6
����y����@��������{�zL�ۃ�W?%�#� �=��X��Nf�1ъ(G��-�9�����5WtZ�f9����*����b֋��PMȱ�&���rӈ
���n��\Da�!������W��-�rK�����9E���'�F�V�<G����1�����Do�g_�ԅ������JVX�@Mϼ���h����m��-��4u���ݖ��;��Ӊ&O��8ͼ��>���<�vtjs�*�#XnT}6����\1�I��rٽB�C|�&v~��ũk%5�]Vf5?4@��40��Q�>+Z(�xd]�m{�T�h+�f^f[����fTX~���X��J��z�������dyf;��������Mb��ڦ�*K���x��E���w�����cn�׉��ݽ����7�|��.#���, �<Z�E�jA�Z�ybz�)Y��t��F�ǥ,�� I4��s[@s4H\���>���E�wR_�P�1��/���>�?�^�	�?�����T�}<9mٍÔ Ă:o���p��0�t�8n#��M���!����0���V3)���^�m����)M��vwr��J�V�X�EXge2J���(���S��E1�^P8F����d|���h�]V��vp��s�XE����z�E5y>�����M�'#�p�pߓJ��e^�1��eU�Q��UҀ;i����Óp�S<�6izU��3����9J���P�~-c	�/�j�$["���Ĳg�kU�`Y��ܒ�n�)�{>L#�R�I>����w�4nxd�����PU/O�i�8�c�� �m�"N�5^��<�b�W�ϼQIb��;~�5��K�~��{v��/��Q�;MzpT��_�m�i�U�@|�Px7���^G^�؂�'&v�Ð�"3M�HZ*z��>��*�(W��wp��o�u'3`�r7k�A�#���٩K��K����V��/���I�gi"�n-���H)����_��gu�:��M��[^c�BZ�K3~��kp�
��3��0��63��d�EH^�S���2�w����=׍�Ql�}�r����a������N�;l�:��]�2I���O^���؍�'8w|@C!��Ԧ����� �� �;Z8�t�f0��� ��9�T�5T�h�:�qZu��>����N�^=oE Ц8$���ݽ�7_��nE�=��YVc�x�b~��+�2�	��*�w'l�b���RoU�-�k@��K"���-���m���ru/�Y!��N�h =Ϫbm��0g#�"�fv���x�eP'=qez�kOᾳn�фR�Bd�S�Uph$�Lejj�g\�%K��u�)؎��Ж�C���x5E�?�	A��;�dX�?�" �
ON��:	+����E[��{v��O����{My`�B��f��/Dpum� iٽ]���pѕ����Z]/��ݒw,E���eme���3pڹy�#o�H�)�:MF#�������l����?w�(=��<f�����n�/_����|w�݊�/C��H*cm�l�v���?>�:�����Ũ����Y�P�Ţ1~�e��J�B4�O�(�c�������G��M���h�-!0%v��Tx(�;�*�P�3�q��Gģt�d�������5�9=ah�oD���̩ K!d<1�D!�lڙBr}4���2k�YA��sH�c�!oƓ�u��[�L1��%��~on�jjk���*�x����[T�f��f��y.[�̐=@����[����]��ʡ~+7?&z&w-v��+�c�.=�l�:�g�^�f*�edpB�z�Ň$|y�\w�C\�>�`Z�#�q����6�H&��d<s��tu�[��"M��}�2Y4�5��9�]�=���OƢ�U��y� ���
�r��ε�u`3`m�U+�L^�%,����-��/#a��B��{â���Oaٚ�U)vZ�I��%]<�7V���b�F7�Զ��T[g�%���vR+j���2?��6G�r�2�a��)s4K:}ƿf.�m�E������h��1�5vR�a[���H�Z�M�(��ٛ�^M<�n?#H�:���Y*(ϙ��X#��gD�� G:�������v��2_������OMK�FJ�����	���0�L�������j��-L�����ҷ�\�/�Qi=���#&z�R�#�~�vo$�2z7�z'v�U���`��GU�WŹMt��5��p�2�m�BL˕�.ڭ:���4�W%�BР���AfL�y�������Bw.����Ւ�t�{�H9� ����4B�}uD���|%�/1N>YxG�1�|߇0 ��������u֝?���w|t��4�4�
g�|�P.ۯ@W�?�
K�� �1<c1�jT��oEG(�P��zO���7����ښ~��;_ �D�s��_/�i����a�&u=��O���A镏�f����>E��<֐���{�8ڍ��E[<(t�Q�kX��f�F�O=�?������E0���j�M`D8�4��$s�\k.�&�~��P��&zSU?�<|��'��'��}
�T���i��קQ����i�Rk�P����/���4\��eT�``r�(�$��\�d���d�$��Vm	<�tm̾]�h��DJ����88c��LKg�N6�eaթ�Q'u��+��ׇ-�.V㌆�S��<�ք�rd�F�6��>b&�?E���$�Y0��xĒ�)�'I�t�UKu�K�PO a�gf��bp~�!~S�Yעg;4`θ~}����~iXBZ#��-�\���ǒh-���E<�����+d9�(˔��r�X#������⌭f"#�jڛ���C�=�97��ɶ!G�����^Ǎ�#�P?��U�<J�ޚ� a����@���sJ�����F#;V�-��`'�q��3:k�ml$@tԧC�UU�W��쳠<��B��~I l��C*	��`��d�vV��A8L����|<zR���B�����R]N������{$�[����Sfr]��}���@��5D�34(���}�I�s%��Ö�B��8/S��7��B@���H�
���&��u���eҨrBt� BK 4Q�X�]��D�'Q#����v���Tw�Q��a�]�yE2��a��WJ:��o�x�?�ѫ�.��;ra�$O�M��6��N���r��������2 u�c��k�%B6�	b�T�]����i���Մ���6���
�&�=\�R%����-��Q�v_v��D�t��^�m���YBe�����OE����6�h����t���sD������8&�U�E\v-��0���j�r��D��%A q&�=�WpC�Ժ�ו^<qXT��2�9Ջ;p��I�%	�d:&F�ά&��u�)���t��UKM��!�w��U[�^�_�[�I��:�|�"۾Q	Jw��N���-�O�u*S��OB�~��&CC
�-��!�fj]Jі6ȹ?�&�A�'�Ȱ�Ħ��ii�R��N��Bէu ,r!XgЃ�Q�3��?���\Mה_a�����_M$@[��G�$=o�2W)KLx_��X�4?r���xW"�s�N%a�P��*޴�\Cy"B�Iz]��T��+S����;�+�ը���
���� ��BO���J�AS�1=�hFc�����/����
�T�A�k�)�����)���Yx����W'ȧ��vU������374����4�
)�����;�+""i��	��N��;M�^q�ɩ{4�",Զ��[������^h_���h.�⫈����@���R��dV�L�@pk�j9O捊�J���t��{N��JIc6�A~o������HC8�>���?+�$!��u;��t��_�̛��NB7j8S���%o,p���D���N�ϳ�\q�0t5Au�yfF��B6�Y�5*��j��"����.V��]ږ+^As"?(m���>��)��RʰYr���:G6a�ƃ2��Ͽ��Ԗ�r
Ο��Y�6)��GC��}�8euF�CpJ~�D����]gy�]>�rh���Hs��`ӓ���:k�`�;����	���-_ɏ�*=��`�'�Z��EsB�U�=�T�fAdX����ULռT�"��h�b:�������A�y��,����?ޖ�,��k���$E�H�FMr��3
�>�L���pQ���kY
Q�	�0��ϦҎ�lT�m�"���U �:��VD�?����rl4��w�+,.Gn�/u�k��撧�l3���ǩ*�i��&���}�"F���)�5���ta�L.�z��^0�${��o.��
r1�y�r��=�|���T�y7Z��\Y0��Oq?��{�L�7p?p̰�iH�(oK_6�p�`]w�e�+��Cs~�p?��r���R�m#�^�p0�&�glitZ^�{�8P ��Ì:����	��q^���J��WV��Yױ�.��(vZ����d-�X�_�⊰C�2����1�ˣ|�O�h���۸G`q�|Vp�M���w���4���B��cQ�qߵh�����QC���K�C��N�B���j�>YM9!K��/�}cX��)����G��#�+��8�� h_��Ơ��Τ�S�Cn5iz*���\�Ƭ�%���Ν�a  �\-�"3��� q�s�8{z�<VۊQ�o` �P��E��chb$��};'��<X x��cw�޳�`����Hz��%���R`���+�H���b��
����Ҽ�B�s��U9��A�LoY��ê"Ǒׇ���P�AV�{����.��齿��920�O�+�Tsh{/����2�48OiO�0d�DE�7�0!
���us�M܀
q!G]�;�\��TB1J�1
-��k��d��gB�s
sݡ�ӛ~�<�%�ӌS����K���G��+����K��dd�`i��;�.�iK�R�^����uzv������!���_#��!h���r~�~Ea1����� _��h��f~(3S�lu��[y��|��Я#L��lLp�BrQ��y�SMp0�����|4�u�L�0,�IB��2�j����U�!�_�<�o�������U]��W�4�i�@�����R�n�Yy� {	�F"z�l%��T�t�aK����ǒP(7)��H9��y��L \tm#f	P��P�Ѕ���9���2`��Gu�I�u%����AO���r��:pae�Jg`�d�	�9Tү������5z�?�d�o3�n�,VJH�u�\,�w2:�}�u�ST	��0bOn�j�ً�#��(���{�i	O{����j!�h�Li��?�[l�rU��{�U�@' �;q���î��R���
����.�/@<�q�����R�|<(Q��S;�E�16�Jb&��ɤf���2COH��d<JԲyqV]�>�=s8e���#��o�;�fi$</�3�1B�һ����03�wbV��T�¨*�)E��A��X��&���0+Q{�����0�s�Pew+w����Y8/�u
Rpm�"���B��G�cB�c�ɶo��u�A�b�|�m�������3ȳ�)�B��5�/����<�E�ؽ }~J�E�� �Ԣp���qh�z� >7�pL��|d$M�0��'���9�@e����m�&,ӱ7�΃9j.�l��W��y�R=��]���0�\OB+�Ϛ�Y���n��!��ѹTg�Gp�,�F� q�Plp�s��Z�YG��Ø'���n��T�b�����$U�ϴwi]��ѳ����k�R�6~�D�Y�\_!p<��!��,���<�:�Z+G�l[��Q͵�sc�>����@d�wv��g��.�w1x�w�$�|\2>q6����� ��_[���E~z�V(	x����9�7��v;Z�탰�Uk����g�a���G��;²wt���<|rk���~<ؠф �#��oG�j"����`I�ņw�b�;O�����d�ka�۟���:��7�������G�R�+Zj^&un">���D�Ӊ�W�'}M&]�rDB����X��lS��4�
f�N���5)
>m��D>5� ߔ\Hr��j�b1���>W�M��Uv�9�(&��|Hr��P`�eF1�<9�S�U����|tӊ/`��ʨv�5K1=�H�b3��7N�!SJ���=G�)a|��L��Kyt�*���U��~}Lڢ������t���Sv��~�)N�t{5%z�j���7���	<2P�5~����ѩu$x".�ћ���/�և���ղ�.r�
��*�Y3Ep��÷��=;d�更�����3�e$�Y}v��y8��j5����zڳ��qJ5��h�UJ��2���J~A�˻ۆ��Y�Z�9������J?���Y�#'�]��M#2�+�\H]`6�49��;���L���j���z�[t>��g˱4��R���U��
̼����so�U��=�۫|B�+!'��&�;�p|�u㺁��FFZ���
�k����$��=*(fdTN�<���E�E����k��1����̨���̵���G���AOۃ|�=�t��R
%K�����x25�,� �_:Q/\R�FC@�|O��U�	�^k*h��wٺ��Ѩ���c�>8�~q(�i6g��8�9o�M���5��5�x��p#~�VeS�&���]��������N���/��ל��ό!Dz^J2Z#VJ�3�����
�s �;#a:��g��(/h�8HŦ}�t\! ��m:�������^iV}CrРrbCj`��U�fD+}�l�csH
��B��{�)3K�r�6C�c���:��k�B &��:[!�>�Օ��x2�c':�snz��'B��"���Йjy}ǀa%:܉�p}���r���hh��K���C�rn������;ej7b��5�)�FQ0��m�Ő׉���'��֎z5�-��Be�6~�p��Rݰ�V&���VϴkU���	�j_M9�4�վtE+nK�������<̰��2�<��pR��H��-���¶����}��j�M�
>�� ��F8Hds��Ad�cD�o�j9fM9`>VVӋ��	8�NR{7�$�t]� ϙ
����Zܛ��5��h֮����@>���{������s���9a�u�ͫ��u|��/���B�)X_���xL�5/�hr�k�>�nbmܛ6������ŷ��KTݞ&�'g��8s��w�=��'ߣ�݆��7�8�{T?~쏌r�S�|]M{<a���=��l4~�h����,�'����L�o�(���ރy"�^�.��t�Z~����%&��l�څ����l�S����;1Gwkܰ�u(F)���v�2;�%�U���7fۡ�Ķ��7QW�Lf��/v�觅0}��\evl�~r)QlL�h�<��Q���{JBx�l�z�b��"�Y�Y������'�2�!�&>���g����K�K�.��U��J�£='�1��%�a��ѣ!�̞<f�]��k���Z�d@G1�3�L�����s1����y�����*;���9a,�(��l�6�q$a�궲&��8"h�q�vK����1���3j�ʦ�LR����:� 8xN~Y[,�XdÄrx�|���S�����x�N���p�y��}]�,y*'��n	ղ
�R�QR���aE%���tp�ʍ���V u9���Ee�r8�s8���l��A�,�svd,����n����qi�����0� ��k��<�+M���& M�L�Lx������()�C�]"��&7�v3sN���Uu��(UT�Q�؉,�f�'�r�gV�7P�C���Yi��`,~�.���Y��g�G��dyB<R�F���|\/8�v���-���.*%vb�X�C�������O����������:�ER��瓇RhE�fm��oS����F����(i�����纘B���iQ�~9��]�I%�8&�K�����d�P�����˧��|Y��Bf;5��$=,Y�]ϡb@�p����"��?��bT��}52�[[����,L��<H��s;�agc'�q((������!Yv���40�Qu�>35��@Gu���������64�\��i�J$-tDTk�}�\��yl'�$�@d��0KR�IgI�;�ڇ��>}8�[�%6o�`�ei� VyG"���:��
�sD0���a� �����@���ܴ�ზ�G�0w�w�b�����'�p��mu�8MRsw�F�izT@���&�~ϩ��.�_)5�.�k�%����Q���IɚƇ̴����ѡ�}Rk�y��EP�� �\�P�t����13sE��+�t*�495+[(��BhN_=�^��@GG�a@팱��WA%��pXl�g5EV�3xqjjJʦ^�^F���O�S*k�x�E�����ǇJ����;�X4��������o޷��Rǔ��7���_�7��Y;�0�:�ȡ�L��n����Z^���g��@���{���!"�U��9qr��U��T54x��U��K"�f��Њ#�a���jF���Nt�B~�����rG��c���9��vE����sn2�KF����U�4{{r�8�!��:��ٍ+ �wrY�G��C�����|�2uO���o�r�K�a6���,p�Nۈ�u	B}�/��:z�4�z��%�R��礣��j�p�+�/uq
�H��A���� � �����á�;��h�2(��'�X���ip�@S8ySa���G����_|��_�jy�i�����o�$�B��v7��3����\����˞:�hn9�7��Tr?0*�<���4����C
�А�L� ˎ{؝k��׆�d|ç9Y����X�����a�E2�g�׌y5���F�����P3T�z�*�u�o��4Bx����T��L�L�%�Q]��E����v�Bb>1��8|��Ô��"7,*�	f����i�t��m���a���5��~�	
�xq�'���6����`Z
p����`�Q)�?|�$���%���D�4xyǯ�?����=��Qgͼ�5��/�_ �G'��TD������S���UmK���u+�>Q���md���%�Ȃ;N��!3)rJ������֮0~�<݇��"�8J�[����X+S��&���|䇓��^q\g��1��[MY������DY�y`'����|��}pӒ�N��K;z �
���I[�vh�]����E ����e����3��i��.���������!}���됵}_��pbt���=�tRe�����X�z���"�N�h-���Ɋ6
����h��b�F�����9v�O�݀ՄGm�[�6��ᾍ���X�����/j9��Px(�-�K�;ŦkI�!��ʖ'�m'y��% p�
F�o��9� �����;%E�H@"�p����N���"���$6�<#9�R\��e	��6��x�%����!�{�F�yd�V�ۿ%g��G��,�V& l`nI ZA@�0��L�v崦.]��GD驐ǖ���#�=;�^dg]����l^�3���u�9ڲ�ꄔH	>���y�?$KVx�����!�9���kB=��\�i/=���qJqU�Ao5�ՙA�X�<LZ�� ��`�𵄷��]e���N<��U�(>(��yMґ��pTNw���_}}��������Z3O�-�6�L��'y!2�-]�����G�(��ڼY	��^a��D���Z��Kq���4�,�B�f�*��!7�8 ���Rf��A(˺�i��׹1�Z��;-{��V��o�f��M.�xT������_hS�O��R�Xf����0�ٓg���b��a�w )����0��n�#�A�9�Ei<e%X}�z���30n���m8ܔFꫨ����G0�Kޓ��\~�i��6r��3���?��t�s[c���<L]:�
3T��=GY�pv�d )!JZ�?�Z��Jx���(}?����]�]�O�B;L�T�8,%��7�K֐��XJ��Luz���)J�pә���B��� �A�̑KIz�Y4���n�
�5|�O_�f���[�5.Rs����{�ˣe�$�C�.m��BE��0Y�Q��,�x��������h���
���BRU����&�I(Ռ(�]P��G�W!���:��Q��-�C�Chw���U�7ҷ7)�Q�/��Hsx���\w�)�܃!\��M�v`7�.��kh�5Y'N�'k͌��~��θJ]zDN�Ɖ0&�5R�n����*v^t�`VK��A�Q0��W.>��E����RK^���g��a�K@4
ě��JrJ�]ZP��˿��ǃ�fm��]�p��<�b�,D�,`٬��:��$K���H[��zдv����c�����2;~9���������0V2z��=��j�JSf�i�K���~�U�W҈�������+$�P��m��i-�I�`$���a׋&L>*�3�E���ħ����@�PP`�6�t*��ɘ�-N��e^�v��Mؗ�z�S��TD���L�!OEA�Gp�.���↹N��!��T��ùY�wHp4c(���Q�!i�� M�O�z�q�t��>��_�Z�V��L$��D�-��RO�-��!�Y����̼4!T^QAΤgSp�L� P�i�M��`qƋ�u��)]�}�ũ0���0on6e��%��崆�F7�}Y��@����r#R���;j�4֩��~$CԵ��djd��3�낕��m~i����Ȓ�x�S�/`�IE��,'�V����B��䨵�*���(�.K�pX��m.�wb�w��z��W�S��p��q����u�?�K���ʳ��)%v��@�.z�5M���tǮ�S��̃at�C15��Y���<�4l�2�p�;��l�ِU`~1��t�QR�/!K�ѫ�q���7�_�=�vA�-gE{���8�9�<T9����!�K"m7�����v���'��&`��G��F�Db?С�g��4�W�7Iz��#��p�*Kd�L�1���R_����JR��f�	.��6��C�N�5Ò	�g7y��]18�}醝�{�}79Y��}��d�\���j��"��{�:�n���J�6h��91�Y��Z���5�u�FEe�5�I�:�����z=`�i��NZN�����ַܱ*,����*��ڨ�cLN'� I=}�橄�]����d� �s��E���S%=;f���@=o}wNG���J��bm���Qq����/@A���}�3!�����2�_�ZY��X���J_ڲ�|5��:<n�<~;s����%MȿV�R�t�=k}�����څ�S$-� �4�4�VXЁ5)#�r� �(5Ņd���#g�u����,,C��p!9�92��F�1�x
T��kȴ��#~*�����6zF�����ƨ�[��%$�q:֒H4� �9)������>zXXԜJ���n�]�uH�dG���/�w+��X����D�g�b�F�(o��~߬L��}xы?5(����+�@�%����t�F���E�גy4@�����#��CB����8���!g8H���j틋�+Yv�*��������W�47�+`�vu����Ζ*�J#[�YiO�5�RΦE�א����,T��\F�{��_ {9<ُ�v��y�o�?	��8T���]��G��D���0�6�.KC��Q��xcXp�w<�t��}�����:��~�>O�*�9L�?m�4R����f#�0���LaX(N~#���@C���5+c��u�4�=��:`�,o>M}�C`��VY�F��A�_.�}�7���,5WE~"��WO)${���M�{q�C��rt`if�~�S�,��@ߣ��tXv���X�s�o�5������g/�@���Y��vF������Mu��%������Wj��Dnh�1�a�ˁq�N��IHU�~������V1�S�H�]x�C�H��Pp���QDC�ސ^��B�l�<4A�;�o"x�͏4�J	�\�-���g���J�b��2!r�'��}��1us25������q<l���I�0<}"���Kݭ���������O̩,��9�y�mĈ!��/��u���x�k�U +�!��r5�_ΎX&�s�*�o�����X�l�9���b���o�ր���^e�Xpv��&���W9���x���1�El��_yә�{W/��p�������օ�q"��$��� 3�\��k�Lᨹe�{�����-�8K)Nz)�H�������,,.�<���IX%��y���"��j��q˾f�3�;z�\�|��[�����%S?D̔@�y!R������+��	N�,�O�R��~�.G���=i�z��i�h�y�q<�6��Ŝ�/�tBYM%.]�Z���Jb��ب��U���D�Yvf�%O֦?�����i�5a��b9\�Hћ�=���A�N��"A������뛀�� L"�O��4��D%��p�JE�,Ϻ ,E a��h�}�8�؉[�K�OE4�A7�Oh4���k�Q�8��"ƹ�
f٘29r��>Z!��+���n�g��<��V�+�o:�*�i?�1#�դ�z����i�̑��[���C��iPa��|���xR��:���b9�|5��5���5�@+~�+�C�dm�pj�nq���������dg��X��䥨���|Bod��$�$_៭��ӷ�#���Ʊ"8ۄ7�$*���50K�l#����l�ւ���"��3WNn���qCzv"�ik�$x�F�0	���VY�{d�D>�6��<wn�6pP]�d@Xhת��]����W��>�Wƺj�'�0X��{?����;]a#����pO���j�~Ko���+|7�B�5#�u rԥ �Ηt3�)��k��I9�]Q�3�������Dfщu�}<�bW��c'�o����R�@�ܼH�iKI��n�e��v݋�kG3��@�i �l�?h����f�Y݃(�s�}7ZDQ8�'�~�GV�^���|ǣog_чP�y�v@|���b��d^W� �m�j�2-�Y��� 0�q���k���*��4�eZ��G=�pd}39F�L���/0�O9������f}��⦖K1�@�5��R��G�
�KK� �<e!jJ�ԍ�#�+Oɇ++f�{ѕs��֧�X\t�|���\	���@�z|bu��I�j0]j�W�H�Y"��>M;���
hT�tm����X;�����&m�c��N��ڡ� �<j���h�FˁE�̤0�u�N:�@�cOᯞr	k]��YA���{߼�u�aW�{� (�v�
Q��`�g��lNELHnl��y��ȀC@���g��`g��	��?���3�Ő���%��I��-����_u����P �wTgN�V�~��Q�Gb��������y^�ox/���������_aPX�W:U7LXiQΠ)�����Rf�l9X�j���C>1�$��~]4��U��$���ehLi�h,E2�����o�jU���F�*��40�O�+���
�| p��3�{�����gcd�Ҵ$�ڮF���z"����'
�4/�*���1��rv��p�U�<K���*ɪy�9��>n�}a�;7�_~�c�սV��Zx{�|����r8����^x����<��L`��Ϥ#�!��ٮ�|iVw���^�Q����]\,�"�⥹�qx����d�9Z��f9k�*XR��t�I%�Gb��{I�u
�]D7d�񌧢�ݍHh�r��+f�Ҹ����*�{������2�[�R�1G�_WpF�TY���� �׵M��ϤNL�,�� K��#揫콴������3c��<({�
�R�U�RO�u��u����f0�g���Zκ�,Y��8�y�Q�ȕPן�_�H�K�ֲ
�z��$�OWF���Se�~�b#�SkB�3�a���6f'��"��A��B�>t��aa=�zG��ux���������IR�mi�Q4P�B��t'bǐ@�{1K|��4�_r�;Ki����o F֦)hQ���% b��:�~.�I[��Oq]J2^�U)��v�EktpW�1kzl0���� �5�f��PP]]2�NJq�oD:T=N���w���X�`���B-PdiR�:kJ�������ka��C(�����㺔�νq��Me��n��{Y��e����Y`-���q:Kڊ�<>[�m������@Oe�J�Ԉ�vд����d&��Rh"�� �]�v �đ8�"�e�Z��&�@�87V*��`�wEO�#��$�n*��JB{; t �L�*ٙ_���bb�}V�����M�տ���O�݊�L�n0��)!{�5`���K%X�S��%��`�R.6�˯ey�q�#�r�f�8B�{܍�Ȑ��݊���T�gC��YSa�烵���V��e|dz���}U'R�H��5��5�
p^~4)�� ���i�j�ڮ�z��Z�Ba��(�J��-C���m��ᙻ`���l�!�G�F�����|⼑va�N�
�;g�ZbO�� ��!@�z�%p��Q��W�:�Z8���&k�n���Dk4� Zq$zWr)�n�<L���Ko��yh���N>��X8a�k�ۛ��NK�0�M����(�L?%��@���E�W�|lL���\�%dma�K��Og��9�P.`���ax�pS��t4g�C11��VKP���<���&���G��@j���A�A�a�L�#���:@���N6�׎,8^g�M�y�c���.��4�=�#����fGc����5be��7�"�d�C�N�pN��!�O��+��G�B� ����i��z �D�lX��=�e��k�=����
*F�]',@!���[���vFc�`��Ƿ��-b]��%[�ݨ?'C�-[��3
�4ph���*ǒ��E�w�k����'-u�%e^߆?�|q�5���	���U$�:��"8,�#|)ȿ�}P�T-Ј�
�0�"�q}r�L9�U�6k�rMq1�C.��q�H��Φ�2�+�el�Z�3C��N�HN�3`L�N0���냇��W�ݏ{�ִ%���~N�����מ�'���Nb���W�(8�6���� M�.��X���h@���9zw,���z�<����{�Ŋ�B��ґ�f��L�ߟ ��2sϿ����<Ƞ}����1��Z99�6����t��a$����*[�խ4�x�\�+�{�	�@QI�l����h�Dy�Kx}�!�"l������:��@�݆ч9p�S�;A^ ɀBa}�������PrV�f��:@r���^N��k���.`�GeI�w�JVa����CW��9��d�Pd�K���j?�� �e����l���|Y���J�
�3(5|,/��i 
(���}�%F�n�Low���Y�Q�mBy��f�������b\��,����T7s��U܃ܲ�*:X��.b�M�VR.��$�Wm)��j6�`Ŧ]���ia����X���������yia���z����j*;��1��p*�u�v��Y%<�SIk@�Ph�TT����y�j�@KG����nNw�5�C0�:$�a��:1����;dq����A|�Z��1��*K���=w���Ao*��
#�t=��K�Ez^�㛞�f*xY����1#�`�K"���y��U��f/�K�5��!XIP����s����O@���A�%e�p�->G��x�����4l�U� ����g�?zc���!�L[=ң�80U6^,(E.���+��eB�Sҝ�]���fF*?|�Vk�I(fm��"G���Y���r��"�#�G����rR2��r@$� ��
���ת�k��}��������?��c$7��J)���9��dZ~ꭻu9Fn�{���v|��xi�a�h�Ls�t�W|kR d�vy�Х����ߎ�k觚���~�n��q�g9Ag��U�Z�jg�$8g0�<5�r�`�F��~,�5��ޜ��R��'�i-����R�������7�<���D����R���l�*�s����X��%ڋw��2����f��:P�cL1Ri"��]l�,yP�5���{37�h�f�P8چ�D\U~	M���K"z_v�$�Y5saB����ڷ��~�o@���>ۚkFy��<�@ W�/����.p�Q�%P��r|��814[�@��3����79TgT�G{Up�Qu�)����ӈR0/Ⱥ������]|��&�IEC=���7ez�m�,<��1��垴��>���r|���ִ��uX*�f��%���_/ϫ+E¨4M-��^$zpR�xk�i�
�]����Ooad�M֋��Z|J���\X�Ҩ��sy�ސܽѭ�˛W!��FI���š��S�ɄI�$o`��{Ù�`u�]`Km�s>�|Q)H�"���$��bN��Ђ��U<2��#��l�@�h$�s��ݽ_�a� ����_T+ϙ������f�~*�����[��#�fޣ �Br&F|W���+�w�r�g�r�.H�C@�ZN���8':vr�LĚA_��g����Si�����ʏ]�khݍ;h���MG�Z�K��{���*q���H�D-g��!�Eσ��%&B�f�k%�M%!�@�v~W����
@���o�A6� �(�,�f���7sN�f3#�j+y���������O-{G�qee�C��`(��SϾ,�,����sʁ�i�8��G�_#�\㈍�L�JK�:�B���R"�?�D�.�Qdm&g*m���g֟����gj�l�h5-�r/�c��HIn��R�w��x^�Cg�[;V8�V�l�#�vRt�4e�+ۀ!�w���/���G��AZ�u������ck�^��v��i�Qh�w��U�b�J�;��g��u�v&�F4�Ed$P�L�<�
,�1�#C�H��#lAh������M6���qE"���T"�tŐb�fǷ�#����+ș�i�@��G����M���p�}�������Y�]�M��ibUrxeL�����Tj`X�Yr�\�Ymu$�����V��@�y�+����sݣmz�0I��}�.��[@g�:�%��)�>s�����e��#�'�?u��Nn�w�ժ��zj����$��>�C��d4�q�<f�$���d#x�(���}2����Ӗ�	���+0��Զ��4|�w
�.��,�+O&H��q|w����Yiu�����(-��v�n���I|�Rxx�q9Ո�]���h��+��p��sȕ��^�[���������q{Of^P:��_�7���?/�WW6��]���_�q�%媣����]��J*}wR�F91$o��K��&���1#���!���������t%�Գ���[�@$��������N���4z�K�����~�7��ϧE��s!�r�����(fU�8'��vʫ�S%��V�I)"ת�#�F�������qg�@����/P�0���X�7q0"�5?r�,��Rw8�i��W�P�]�<�&mqW�+�7#}�X�5�i����G�=�S��:�ӹȟ闿c9*�Oޮ��7�Lg��� N7Z�+�y��96ص����Dż6c���������N������|���c!v�I���Cffۼ��/���������~��: ��x]D�H�I�ٳ�|ik!�#w��$���Ѥ���u>�_dLy��$U�3�XL�� dS�^�?� �:q;�����$�d����������Db�L��i6�!>�ʓ��SP�2���:���HC�	O?��v[xп:t��W�4ߛd�}�� ��'���f��IIh1A�hO�>�@�x���\!�?8|-�ϣ�T'��XJ��%'v��\rnX��Ӂ�-I�sO>y�m��Ř:�4a�Hۆ�WB�{Z����o�F�%2}m$*�e��q'���w�yL�v���X��:hn�"����}0ʷP�F����1O��Oj0�*(�SÝ$`��	�?1��>�.�ene�G���A�M9�����7i�XJc`�t/!����cI, 4P2%IV�Y��Sz-i^,�����Tj���������FA���3`�
�LE��o��)��<A��1��Q���UQ�5�s-��{-�@P�?�5�Q��"���_s���m��S*�u���m�W�]@yV0�O��2:7ׯp�7b��㷤�3�*��L���eE�P�Z���2����`��yttӉR�A���B�]6e�ڸ(Yu̗F���5�NSc���e&�aG�1k��Tגљ��J����S Sԡ�5�)M7-I�Eժ�_�5�&ZH��s�����U�;�/Xӓp͔�p	�H��M�A{�|W�� 5�SW��MI��3��sk�_����5��a�x�Ѳ�.ثg��q��D��)���0܁>,z���d���>�}8{�ht�L�T#9{��6��xM?7���y�zĳ �HJ�RY���iv3���?���wMFb1T.��7����W ��t���\�B)]����_й��p��>��W��]��5+����H�����b�<b��'���3��6�q���]�J*��9rQ�A��%wM.MɮZ�;�PO6驪ͧЦ�<�dM��V��\�V7�V>���˕��]�g�3��F�Lq5�'����@n�o���������-��)U�]��]֋�x�r��u�(AC`���f��#�T�hɣE&�l#�3 �$OMH(A`�Rʍ�o-�Jܿp���������~۝�p���e�W�\6�����1�G"<��O��ݺ�-t�L�<��jG�Qm�{�Y"$E���}�[QQ��9�����@�5%,����g��t������5Z�������\v��Ϲ�̜�Qc�H�eM'���e��&cB'���	$���&P%��;�8J�@��
���ċ.\�aW�Ÿ�G-3(�V3~����Z� C�-���Q��G:QD����齘D�ͣ�I�$��(�>L��� nit#F�p������|��'/J�k���3���c�@�I'|����F����o�7�Ǫ���P�v�;)�z����e��e��\�����`���葝HO�U:��V�S���@qN�}�&���5������ր�C�Ȑ!"d��9_��Ⱥ2v�ό���'n+gԖq�)ˍZ�����4�a?sG�T�hb�9�t�C��iI��Ԧ���2#j����0N�l��C�M��J/��e
�	k��'~x|���J 8�h#zc�k�,�(Q���9��:eT�;�֥}�;�\�X(��.�}��';nE��%��s"�as��H���`�b��tӞ��&���é�C�o�A�,�uInpGz�h�`�ݿ,¤P�]��L�/jz�~�p���������y��RT�q4��"�%����E�zB2���O���� ��X1�e:e�'�'�(͉�G,�^��` [���C��^r��ޤl�j�R85��rw�����D�v?I��D,���ju��B�~�z@���B��#�����ȥ�m<Q����tXi۵W%��ٵ�$X�}1�Wr�|n8ܔ�LL)�N���	�WC��.`[ʫ;�bPT_�8r '[¹����h �u<� W_d��,�͖ +�`�~����(+��l�S(��à՜��������	��,��5��]��gDӠ�O�g�TZW���g�����{X]����ӎ��i�aӑ�`���K�#�0�s#��]�9&�� 7:I�Z4��`s��8�r���$�	�ߏHb�E`cg�OH*[̵-�ϙ�d@}%�VSܕ���,?�9�J�KVDv[a�$�u �-��kͩmu^F޽1����2o��<)h���O����FE>�K��<�I#��΁PU���ǐ<�Hdʍg�����-Z��y}��]{nс�߅�.�s�i��mm*�0��R�5�_
çgOs�iBa��'Y� �=8����M�L��b��@ŕ�O�`]�Z;8�,AY���W�~PA�����@&N�|����y�����QcPf���k ��Q*�}|Y�2��p�'3�T���h�8��E�MS�.@�I�~%�?Zь���N��R���� ��)�G.Q�J�}��o�ʉy�Ai.D/��"[�� ��$i#)�����D����0ֻc{`��x=��g�ŉ�!K��ǿ؟Y5n�y^-�I�o��J�ݒ'�sq��ҝM$}9�XL�"j/5�SG^ĥv���a'�4z^�̍���+����j#l��C�$֥�&l>���f@lЭ�.���&�m� s�C4tsXh1�c��3]�=��x>s�M��g��;��s��Ǣ��Wش� SH 6U ,s
|\C�5��*Y �k}7�حr�X�[�~6]6g�Zo!t`my�M��f�:�ם;�w�r�rL��c �lV6Q}YȜSc!��M� B�0~���H�\�[�<�b6�YS�68c
�/���ކ��.�dO�߻9�aXKq��\��K�8������3��Y��]����N���+��~9�!���z��Ms{��u@̨;H���p�� �|��M.� zB��������r���yŦ~+-n��
����1A/�P8�������.1�r���5��sh#_�������t��{R M7�\ۍ�- �K�����RC-M�}���ۆ��ۢs����'���U۷�����(�i3������G$��V.�&~_��Cė����+�ŠL�䶭�n��x�o,�D�K�!�ezZ�����)�n7xF����?�)42�>��?ݷ�d9��0���چ�x�-�Y~77�;o�#��Q����A�\�x�3�i����c&U�Fɣ�=B� qYQ��,�Y�RRpu�A!���=ޔ��+dT�7 �a�>M&G�L�+0����:�"���*;O���K��W�H:���c!Z����}X��d2{�[�q蘷"g9����6���f�cwk1Y�������^SF'�������cܤ�E�N2o���"�Z�cT��V���	����B	IٵE����ˍ����z)L�y��|�YG��b�RSϭzY�'���zы��H8��^����hJ�.q-�����*�䳉v�ƭ�e�]��t6� n8X�A�h�����9�Z�>�9��qp����`�o2��gK.�zE}�Y:-��T���&�Gc����$�<�5�`"�uê� �Dj����k+��=�-���ll_x��hJ��;�(�!�w8[2+�B�z3l�����:V�G�^C<5�ڨ��V��-ĺ�Z������`r��匏�i�}�{�����+{<ȟ�<s!����!4�X2��X�vj���snn���+��aI4d���3�;s���WBU�J�PF��=޸Z����KOCIȳu`�3&?=��vsq �O�̣�S<`8˙��]L�`���q�0�x�~��F����MY�n�GK�&���
m!`9�Վx}Q��t�W��9�H�m5ŀg �۔��n��(�4�?Z['��Y�l
��YGy��J,��.�|�<��������4���V]zP-��O
��ޠQZC͕R+ցC��Jj���q��-�Yg� tU(S��Uո����M����Q@���
I����eBM�)��̧��3�"�F�f5F�	�㘗�����T=P���=�)�6}4K�����q�;Fo�'��u�9e�T_ ��/il@Ѿ���%�3/��&�̀�tb�pt�E*$K2.��p#����%s��`�e՜�K��j�l�UL�C��|�C�*va��GI����w�-�Z�uV���9�D+#��T�2��D�'Y��IQo���&g��o��
���L����_f�B���RK�t2�+���4�^�=�J+�o�-���8G����Ƙ�>!�me8�Rqu%|W�Cʤ����A��]�Wh�@'��ق������7MN�^,[�l���F���">����a?�w��Q,?}%4��3J�������}��xE��`a_{��C�i�L�[�3!Ha�8:7	Tmq��6���2A47wem�f�>�ׇ���g������4W�t�(|VG�Z��H=0�ݷ�K��OD��D*�8�6� ?��>�tH�/�ABO����u"7���$�j2�qbrB^��Aէ�p
���>VѺ��y�R���z���<�<��_�\_�XOQQ�8Ӝ�&������Y�N��ZivmL#@��B?p�ڊ�N#c�*�Ș���^���c@}p0*�!�K��D`64'K7ktK�y5O�(�C% Xy1��i�bem�ϠȨϣ�N�9���	������|�VF�B�2<��i\w� (/%�˃z��tw��)B��	H�
���8�r�F����@��t�@M�P�^�2N�u11$,���$b���3\�-5��'sur+���}���M��P6_N�w?�t��u�o�᠘kG��N�zWj*��o�k"�\{E-i��a������&��$(���;������9�@JAע����8b�؂U�O"A`CsQ�� � �������U-���~�<�>�AH?D�!3|��A�ӄ&��l�:�L�-em�ۼЅ�Y���O1��p����;�ȡA?�"4�Po�>��BK���Q\N��%;�.�s͛D�v���p���K�t
�sCI��[�0"* ���,�߷O��B�hY�޽<��0�ēi��]���R'}O�+�͵�@���|�Z~0R�E#
�����*����W���h����]�/����~��u�7ǹb�P1ތ%8@����kr !���"ّ�\H��۵̌��:h�D��|���R��)��RKqq�ۂ��%��Oܹ��U�t�+7`�
Ħ�.Z��d�������H����f�y�@��B�Ţ������R���:�$��ֳnU��R��G
w�@ �b�c��Lpĳ,
�V~$�F9���.r�N���Y�n
T���28!��|�{�8̢Eٮ�Ixǡ�8�Bh�@htR��Ƃ���&��%��ל�4�nC.N|[�衾[R���!�8o���ޘ�v>4��>!���V����m�h�u/Q�_�n��C��vj�.�d/V��K�T ��M��=pw~��U�i�퍑�M�y�v�=�)
��2�ߌ<�����g�ַj,�0OÈI�]�Џ�hM�̗-��Wu��3
������R�x�ِ^��Oz�S�t-��W�t��5PL�E<j~��>HɨK�u���u�;�TJV�)��L]Y���r��،GD�h��q��m��c'$P@�W]	������!�d��x�K�p�k���w`��kg���H�ec^6b�����G~��Tmf9�뼫@^f�W#�Aj�+��E�\!t{�%_��3�;�@q8c�XAd?��ͤDNč��łᏦ�=�]��Рb�T�J��]�UD)1���+�"�.�[�>u����u�(�l�<m�V62�V6��Xy��.u4��V+�Bj��㪏}՝S��X-P*���s�X�F,zpl1�h�D���bD'��S ĵ��e`�������o.�X��d�]�M�7���v;��_�Ry���D�Ցs$��A��W����
7�X^�/6���D��Q|e��;��D����}/Դ����c�B��M@|�Y�*U���l��"D_p����A3/�v�⏺�`�
�HOz�����|IT�+��o��{�5&,��C���Yr��v��qԘXO|�M:�%������zwDs����]�J�WA�٦�1�W��)����&�J��,��d�c����p��mߍ{�ذ�������DD�����Б�IE��q�e�1�ԧq�TE�a��^~@F�HN�oKBE�5.�]^z	L[��U���Ni�g�*W����3}����B&!S�Xx$8Z����C-u��P3����iZM7�ڊ�w�j!YW��j4�pX?���m-Y���Y|>kdo�W�.�-}c�_j�r�`cr8er�tĖ{�XZ0	��+=ABϽ��i�7��g�Wy#7ZD�P]�X��Nx��l�g@'y���j#����WNa�e�4�ة�G���\�y��O�>^ʠ��C��Ro���+~ ���ʤ]���)HO{^��ri:Z�3������ ����W�]��!�x��I�N��%V��i�l(�~=	Ց�����U@[�q��abFZdH9\�Ѵ��5������3 ���ˎ`P�I�9�{��kp1	�j^w̔[��p"\ݭp�N�,v��"��C_Qrg.0�!@7�,[f��(�Ň������F�͂@�ׯ3#�ak�p���3��4s�馱�Y���k�ˉ4��5g�U]$A�x%b`[emqyNJi&�W#� �Y���M0��t=[3Ͽ�G`�Yf�N��t�P�)��x;twWS�/�mf������2ݩ7����ݫ�xȍ )R���d ,�4w�0�]�t��Wj�le������ߥ�`ª^�E�w��a?\���B���#����m��nH���5��+�.�1 $r�f��U_E��M7�dR9��'�����~��4�=x��]H訔�"����m�2Oxy���g�� �DA��6���M�z�/�F�/�GxO�o�hr$-<�d�Y��К�5��܏QR�6�K�A����>{��	ǅ���v�U,rg[Z�K�^��^�%9�z�ʙ���\��%�7��./A:qre&w{��_� �ݙ6',3Y}�d"��m?��#Bji+�oT3��6���h�7OqB�=G4$>�vY�׳d�wfeĸ��Krr1n&�}x�ĩ�2�n|������e1}-�c��7k���ů�A8Z�i��:r?VtPu���3D޾�	_��4�Q�18�D(�U�G� �*z�W78˦�>yX{Y���zo~5.�d��*U��&����a���nw3k�\1�J��[qHes _����0���;ol�_p�U�ݱV�Z['���6r]�Pw��0?�yp-|��![�;���1���[�=�Ӽ2��jK��>�����!ī�E@��*�H!7r�{è��z�k�M��b4n��3%f�P���?��hvL6z>�v-��P�O�W����\��E��5O�j���Хa��giZ��`�ovb��T[߿�a� 0Q[�NY�:�kt�zFc�%�q�mSs��lПVY_HD_�%�C��j`���?R�ذ�z߁j�g��?\T-�D���J#���ݴ�C�_�Cp���y��>i�F��t$q`���O-:8����>�v|l�����u�� �w�H�O���M#3-6�K����c�;���h	I��&?f��N�
3�#��40�}��C�-�Jo^�j:޺����>�^��{�#=t�����`����P�X�_|` d���	�}��_�������Q2�� zP��M���jkǂ�J�r��.�j�JŬф��QIv� ����rLN�Ӈ��f���i?�����-g�s(�P��u@�_���|�0��m��w�E�������,c�;-��\|�K�Om1�q?V9��Ċ�Di��V=9�?�*�`~c��;��UQi��}��IO#i��f>�\�?�;,xLfXK�?S敏�Ѱ����np�'��B3�ĊMW)�����p �xhI�J0Md��M��(�a�M]NT)��%.QM�{<B��!�y^j[�{�^)�n��=�Q���k�_�y��fcu5Џ%�ʏ��^�H��*�y�6��C�~r
iM'��nB#C|҂�[��BwoyzKpյ�{�7ǊG�"���^/>���ҡ�!�%zE+�4�jt0j<1s[��������%ס��df�F���z�������z(��0c�Z;X��񛩷���,^Y��Ǎ�ɽU������):Q���~��N�*YB���^(���;� � d�	�`҉=8�+����1��Ҥ���:�b0?�T�d��������^b]���"�%�m5_����z��CQ��2��j�G�:��I��0��Dl5�l屸i�1%�N͙ЫIl�`D�S��X��Q���q�[�T!�ZFYaQ�D����]�b�t��ӫ!�_�_�ɨ�BZ�y����$eyy��W�Rp�����|B��E�4�at|ɏ��w���\E����Oa|�R�f�x4����1�y⥑j�8�xH�%V�u��-����#_!r��TNR�1��-�Y����S�q�XS��:�Aڮ��M�0/#=�����e�\LQU����r�v��6M�mB�$�yg]�)�F���~�{��]�j[�7�b�5O�mS��\=fA(��Z���"�ݯV��TFW���'
����g��G<gr�#$��-X����E�)�3�iy�E;�JD�5`�o��MY��g8
뜥kw`��5H����u8gL܎2�0(-�r��c�� F�
��E8�����1�bƠ.q���E�v�ئ�߽o����E�1{��yU�R;�sT��GX,�X'��3aX�=�T�D�v=G˖sA[�iG�$:dH�i��xf�J|r����|l�"ozz�sW,��7ς�>�=�k�;������q{+�������WĹ����hnd��p��0M�|s#��������X�l���'�r�:Y<F�I��@ۜ��I�Z����k\��`E@p�8=���7�Dg�ҍ�5�Y�_E��\�� Խ�zt��c�T �k�؂ݬw���䦋h_{xT\S���0�$����+b\�(�>�l$�Q�O\M�y����<�̛V-ؤ�A�c�%Z�:�Mc�fIF�=d����ױ"���O��i7����H(ذ�VYhԟ�ڲb�����_��8���h�M�>�-��B|��k3^c�5�E��=R�
z���^�bJ����=��� �V�?#n퉘�Q���"�e � ?���n�.��nՑ��:�VZ��e
9_���5�+�|�ڽ��]��ES�^VD_��q�����8"���p{y=�l�P�b��[��#��ag"y)_B�^D����%�D>j:�T�{x�����}+z�N6t�6ۮ�|lF���$���?f���G���������yL$�Z�Nhy<����-*{J?���CQ������Y�W@�x�C�Ҝ~Eģ-�h��4��`��p�o_��!�b<�3��c���ר����tbZZfT�S�4I[��5(C��U��w	=7�i%��X3�Z$��U�S�Ȳ3���HǤd=LE���F�&��b3��{5VL�ܳV��C�}��'�K8e��;�E����Y��.8,�S}��MG&#띦��#GUEٞ۵&r�3a_ic���N)4�pl�u02c�v;�S��#��)�AK08TFɈ���?4�E�uǤ`���z�VJ�Bڢ\�� 0��>C�ܒ_�۞ՠ�c=�|S]A�3�Am�}��Î4:�׺4 O�X�n2����츠)@�
e�A?0�er���{�Mw
l�`q�mqHІ�!�6m�_X���Ʊ������`uUV7��b0�0�`��{�]Se�����r���0D���{�`�κ�H|n|��Ʈ~Y*��x��ڝ0V��u�B��z�F ʔR:��w���w?���� ���V;+;M$p���
�K�tv�s%��e��W^ԩ'��%�8�y���k՛��&�.3�,Ou�C����prE�(�ϒO�mC������j��f�D�~�Jz���lfQ�y�/㯘�� ����2\�v�>�S�o.�jrۑ�X�f@z�x i5->g蝉*�8�H^F���Y�>���̈�4}��1J�0O���ҫ�I�� ����ۺ�����rG��7�>�C�z�9��%��$rު�;{�VKUǇ��ds%x̒�qn��G�/Vݐ��̩jo�v�i�Nȟ�LO������Ԏ�q�BZd�/t�+����QF�\�f��\2q���s^����:�̢�	��#�Ej���Z�!���wq5k���}:�]�:D�é�x#Pd��J\pW��k���3�<Ɉ�{�w��N��cpb�S�Ӌ���B�-����U��k\c//)����Yw�`5Daٚ��-��3o�� �^��a��k3���b�ɯ�[�;���C��O�k,�
��{%\�ں1?ۥ^�T��k��=�M��C���!�e�3�ҡ�_z:!�?�YĞ�H<P�2c-��nK�p�@|����r9!��Re������k-�÷���`y5�:���j�7r���p�!݈�X���u+q��/��y��h����4X��V�r �-�'��Ե)d����|I[	��}op�DӽNd�Z�~w�&!*�7ב�zͼ!j�⑗�:���4���Y�v��-�a�6L���8"H%7�4������;X�l*nYF���͒��ǋ���8�����a-�����'��m���
}*P�Q�����2*�RO+	A]�� )�f#�5��Y�.���2�p���6�q䇄,�	��d	øL�����������4%����pEf�'�u�\N�s��|;�� �˽LTD�d�ͺ�}B,��W@���z��Eџ�V(�!����ѫ%����k�\e�pRg�*H� ��b��!IS��?B�-w�5��(T�᪂ݚa����X�p�[�=&K���A�T!��=��5�%T(��P��3���r�~�����	3r3�ĶlgiD����{�|J�~�$~���P=��]^�$k�=5��g�đXC��sY4i?�2�R��6��xǙ򏢁U���~N��ԫw�Ҍ��ta'�1��gnb[R��X0���`:6�'�Wb�8B��i�	?�/A�{O��j2�Zo��������T�������Ub���B5jA��q���)+�l1���dT������2*��{=p]l�,�D#*����_1����zq9��H?�:�n������Ų�U�{�D�sX��2���\�)��a�Kw���U���+k�QI�W~E]ɔgn�v��	,��lR��%�Q~���,�u��n�e�t��u��bPś�͗��	�XE4���_Y�������魕�yU��r+h>Q���Cu��W�\��C�$�K	U"O�
�e�.yZ��%����J�N.���;���d�ڴX
���X��[n~�)����|�QGS��λ��o��2��1�Y<!Ia7������fK�����ˊB��I1��-�4RZ�� ^C�Yďn�>m���.F�M������U����I_���abC�M��u��`��Ր���f��@�qM�mD��i~,[����r0]�`!�L>鹭2��R��M��c�+�� �[g��k���ஔ�Ԝ޿:�v
�&v��	�D�Ce_f�K�,���}����Ug������x�T~�7��&rXݛ����:묽��S'�p��C�HA5�H����0b�(��4�3�L+��]�xM����|pg'�e2�I�ݶ�<���&?kg4`���KG%c������gd]IlL�y���c ��͙rd���{�y½s5���ߢ'�Q����;�?��=��q��3��y�@�Y�zO�ڄ��� ^�e�Q���/L�@�\�;�L�2�*Fɐ�Сڿ'3C*�kIh9�&����G�u�]#��anY�F�Ҳ�$w����L�h�׶�����w��_���a��o �Rc9�?c��Zkm���4�W�ִ��*-�T�G�[��ǂ�\
��3V�����-���8�A
1�C�n%_��I8(�0	Z�Hl�2�߾�D��O�F���'Y^���u�=1-��0����7^�3���7�����|_/QD\�ŗ,Θc���������sE\w?� �GS��.]��)W���v�Skɖ�2p�ҫ��w��0��(��M��� \���^T��� |Giܩ1;�3��1��E�Ҿ*�k�-�D���q�r���!�",=���KUO��U7�$���v���W�&�z�t���E��h��������nD�V��D��G~�"��a`���8/�Z��)
�]^R��q������f����b��c�(�4׿�g=�Anp\a�ɟ��u��g|���%fy&i����	�+B꿌
b-�(}a��t�������'��Ќ�.\�y����V��M���ϲ�>I��sm�]b��>�Q�q�S�q(M��U":��I`R�������O䅺4���)��U{�K ���&�<�P(lzŊ����%����C�����Ci<̆��əN�"�ol;���"nT���	�U�%�Xw�����l����^�hw�Φ�|��6=�d.�:���I�QюG󺶵�%E@�R��M0���Y��YbXq�X27�X�
x,�-D|�YdN{�͟�f0����4= ��s�!���x�������>K<��M�� �9�(�X��Voݎ�f5�7͖�\W���\�������6�[5j]�K>�?Rc�|M� ��0�P*�����*��
�-A�G�<�/�ɤ2�9���<�m�KG��2!�P_�ڢ�B���Hg%�E�ZSؕ��C�C��*�Ig��"�r�W��Ɉ�t�#��>����ID�}x�7�ޕ"j��
#�0�.��,��Ń#s��p�oD�/\]�9Խm�=���M+����֧͘�@�� ��;d+�p䵉EZ!�o�ٯqO~�ˁJ��x�D*�ٟO  ��H/^�l�����X��-5��O0�p�=�Q����}��E�\.�GȆ�ٞ~dA�����͉t��-t�-LN]�<��'M�m������U��孿ٟ�����}��%phX G��Li�`-- E}`޽y{x�G��q��W�jefv{C��G:Ah��c��S9�T񢷸{�n�Rp`�@��Ho�u>�EK9�O ���=m4VYZR�ؿ�{:2��: h"�w��s��J�ݓ����1���`�v�aV8��+@�X�JO�� ����3x%�o�B�8GcĄ@����������]�.�e����:����%2CKr�k��ŔP��m.��Y=N_�4o۹����X�`�]�����s�[���S���*���a�\��m@����4�U�\-'k�Gq���72�A�,GPю;*	�VEΏ̿�����K����^k��Ʈ@��t����ʫ��~ҼU�5h�=r�*��D��Q3ǌz���	�%�l�&Uy}��U� �1��AT�6�xl<�(�1M>7@���}Y-�Z����V ���z�cn~͖�ޜ��
.���vv�J���X��eP�܏;
4v1�rZ�����.�v���_.���r,�~rh�.�oX���6.$�����M.��LM�֨�|��H�h�fmҋG��SlK�+'	�@u+V�V�����;�u����}�cg�m����EdfO1���W6�w�w�.�����]n�(f��w�(�;��ꌉ�A��j�e[6�C.��S$���8ӿ��Q����I��m��x�w�?���W����b�]��ϲ(�s�<�k%�s �J�He�~,�>k�����Q%"�rԾ��a���A$���<��ұ%0n�L��%~�B�YASԜ�O���rq� :t	Ա���ok�p�8��������jRQ��Dvo-Q�&Z/�Hp���j�e�:˳�1
Xڏ�Aѥm6�agh~�p(HA�����!:��PFY���ϬB]��E5|������`4S����H�F�}O������ܕ/&��ۆ|~/�|�w���+hc��Ҫ�x�%5dj�ut|��[�e��3%��8N"v�ȥ���I�]'�Wl<�H�z�w�s�\!�������G����1G�WAT�`l�6�"�i���S���M�A�Cj�+��l��v��,M ���11�֠5�����-q�q�1뭗;S�%�*�ůj�)��ViT�ӿ�Ǌ����z��5A�rS˓K��3�6x����u�iY��ZN��%�"���p9(�9ђ��!|p���D���:��Z�b ���]�L��w�9N�؏+�\��A� �҅kf�!j��Q��6�R��?��ǦT�[�L����J^
$�af�?f��ߓ��F%���2X��m���+�0m5J��KB�2X�|�H����m��K	�l���h�q@ʹN~*a�]�M�V,XF��>Us�����53f�G+\�&?+��?�dR�Wb�^s����/���i�p��!��t+��&K�|���L;�&ӃS�_iI����6X���2�4����$�%��Sӗ��{g<F�����@g�vUaf��.�4�%��ϵ羼�A���`��F?����~5%ӂ��*t��������ga��c}-}dD�U�IO�r�����}�?�G|� �4�v�9@����J�k�Uz��Ҫ���ŝ^�k��@L^���/��>�	O*���ؕ؜�fO��(^�_%�ٻ?�Y���@�3�9,@m��5�l.���	���T������,:�N��`=h�R;o�#��(`�e�r����5��W����8�!�"1��#(�M��nC=�����(���K�,�"h�u]]*���_���P�JaG�)�w�k�\X��|��A���l��$AC0J�xǺ�oN0�#F�Z�y�2�"�%3s�j�E��7R�y`&�+���y�Q�����>�E�=ۄ����.�[><Z�$_n?;��œ��:m��b����v��L��uՃl��>���r.�J�A�ڳ�1�^�jq-8��meW<:�Fj��;�`��t�����'(#��'�zʀ}'���plj���l ��_���櫸�8q���t�I
�w�,��!Xn��8:\����O����XTά������g��sL5��'ޮ1wG���v=X�(N��uM)�~�����A[P���F<�v�mn�N�u�0	���g���'_B@�9\S��j���P��h_��rL"`W@H�Y�A?��m��*z�:��M�f�F�����h/�9#=JvdM����D��h�v��z��w"�|	�WX}@����H|i����s�-�Č��d/��d��cƳ����CZx�o�j��bY�h�����M8}`TG@|޳�LC�͂�5ү�*�j]9�h"Y
r��j� �,6�,���������@G��l�aA�5�=�Yo���芹��uMl���t�wN�ݪ�	�Ś~6C猀��j�^�LԖ�[��c�Ӱ��hEj���T�a�Ʃ����\vʍ�F�JH��� �V�7�4�����7�C���=���j��W� Wܟ�	�!�rY�U|�LB���Srg �P	�K�Ŭ�u��Xj��Q�-���~>�&�-�n<�U�S 98E]8��X�y�󎋓5���9g�"׹8�	Vt �%A��N��/u^�t��C�+7�F��8������b��T"5�rAd���X`d�g�] �PY@lႸ�J�A��'+�q��rP�;,6��ȳ�,V��.PB7�?��ɩ1�$;7�U�{�C��[� +��xX'R���ݻQ��dL7�7��V~�O��~���"�`1yg�:�%+L�Bg�e��v�R7Ui�//�����%��bP'��ፒWp9[֮(f�U���S������`�Wƨ%y=r���m����w�*�ˊ��E{�s�U�5?RVwZE�8��X��י�L(JO�g�
u��p��:��aRz1�UR�2�TX���[� ���	�~��>�t�Y�j��+&����qoŧ`\����-�8�w��J�̛y�}�P��Y�~�ɩ��^? �C������!���bo��0���W�Z���j1^���r[�[/B���p�~�$h����pE�?�I�����+���(2������m=K�������b^�0ry��K��n'���}��m�ڎe�P´��+��ƨ����7K}HZf�w��9���Tfm�\j0�>m��G��ad��)r*'IbUǝ+��l%Gmbj��i��>�E��8yO�^$5Ԉ�%��E���_u���ۊ3���A)�y�3[���*HR�(]�G�^��c��Θ�"�g�n����Q~ ���g�ip�ûA^WIy�2��W{��c��7Z�����T� �3�1_���Z+��iX��0I2���ϓ���K�㛮�,�,AŊ�݂i��z,� =2�}$累0���Y�\���*�N�T=����YP��O�2�G'I7_�,��u�fGVZ���xc��1��є��)brS���Qݴ��n ��zb�Bջ�D͞qt{%�Z� {��*����LdĶ�졥�!K��@����yCW �F�w��SK�X�����׼Ն4g��Ǹš��&�3�֩_�.\�pو�(R���$�z{� _%j�E�~Ib��
�����x�K-@K�,����e�t�I�RxB;��$�b4[i�FOmH�`{��db],/��� ~�.�=g;��k�'�ʣc����l��T���� w��Wu�æo�o�ic��\���M朗]m���2i#��4�uV��m_=Z�{vFo�ڧ���~�ˁ�݃4���E���9��,J����#�<ڌ��R�w2)��ȭ�Z���[�����D2�� �Tڲ0P�P0���>|rF!6u"���H�BRI��\.k�|�������5�\�i��P�.�}��T�Q	�����'z���f߫<ԟ�P�|>�+x�of�c�^���}-��
�)tT�w�3��2*�
Q$�">Z�(w���̛)�8��������X�CW�_��i��G����b_��0/��K�o��r3�h� C�JҐ�G.�����Xig��!��z1�v�a�)�Wo8vZ��I��vFN�V2 �����q5A�K퀑+�������K�Zֽ8|aP�G�Ԑ�����c^�d��X;���o�df
��UA�5���0)�����x�ﯢ�1��]/�P��.q͟�[��B�ఋ�S�:[1���௝��bDH��}B�VQk`?���]�f�bĦQv��Ɲ|�dQWf��Ԇ�I�U�JC�QM9��nqG[>��01]��~�[;a��#�{-��\Iv�f�D�zN��&�ř'�ӳ�q[5��vj��z}���3),��rڈ�v-l���-�:��s'��ϡ��qW�87������J'�+W�f��>c)IYx�AQp�_�.����"i	�4ge�=e���ڀ�D����Svtv7���'W�3�]Q��5?+��	�8�$����ii���1���w�`����I�Oҙ�%�A���툮G6�b�c�+�����tt%��1�8����x����Us�t2D��kv6��`�ە���A�oS.��:f�A)�9Ջ�y�2�B\O��ņ;#�����B����F�}X/����V-����U�A4�������:��EN@���Q7=�Vq�m�0���e���Tߪ��6�v�F��u���H��e����X��Dj�Ə4Q���[���Rl���
9��k��(ci��N8"�Y��b^P��i�Kv��_�
������y��Yb�C��8�Fq��"��h6=l�_M���B�#����x=gRĝ\FT2�/��$�J�ބ��l��џx�{@��ކw7�!&cc/$�L4�1ŗ�����=x���v�f�a�zn��5'���)ާf���m�%__⍗�4%��7F��K��O��vɔ3����-��S��4@�x��R2�
��,�R��F�&:TH US�T��9#�P0uā%��ZF�3��+��*�������s��&�5=II��tZ��p�o���~���/'K���6�VT�\{�I���δNM��y���ʅ:���gZi�w/ �X���!'������_j+n�K8p�<�ş�F'���?aK��G̺���R����W��t|��@�x$q���T��|�����Y���h���}J���@(��!v�.�uQƓ�`�{��P%�R�# WqS��B�@!�Ea�-!�	Ѷ���m�N�]���> ����\L͝�Q�R���]�g��LT�b&��]"���7�7�q�F/�ZQN�U�󡒩=�k�Xoٴ<l ��GG�7����b_�jg���㰻��Fc��s�u(� .���T'��s�yE
����m�������ǰ��n=���˴�A�#�+$TL��������N���fЙ���DN�`V�V�/:_4����e�����#������[&�N1�+�9���ސ�����u+�����uF��ńب�TG[�h�4~�B�|��ʸ=i�������{զ��`��Z*4D�����:��=�A�8蟫����f�iB���c��<{~��şwQ32P#rl�b��ipӺɫr�;�U6��V�P�0�ާ�`D		e.�ڨ�#�/���Ӽ3e;��C�Z�r�isQ��=A�+g�����Rң0+VM6������x�vq���;a���0�dr�v��We�$B��ob����N��
)��c�f{W��(?�� -ք�H�O��P�X�d�!z۪@}�	%�n,�������G��A�Z�N�om4�՘��/r���𼌡����o,����ۢ:�|%a�=Jo�'Nz?T��>��G��o�Sc������>�>�;�
i9�L���|�O��,��Q�
(�l,X���p�6��j��ﻘ_��&���������Ή.}��oX����y�;���#�Ë��Z�aʰ�w��$�#r�i3*�����!��n���_a�qNw]20*1dF�q�a���m4�|ލ|�(��{�(ۈ[�f��*��ٴD	�+�&(ae#�l�v��y�k)~�� ���P�,��`�I��#p��~��@Ģ��Hu�{�f�������U�ڲ��sM��қ�C���4Մ���F�'%m��QDD��O�&rA�Ϗ�b�������U
����x�i�!;jәj��Eκ~��c��R�,��%@�6KL��w<9��U�%�?z��p6xp3:X;|t�Y���}C������g����VS��{5K���ī��=��KJö�-\�;��`�:�i�p/��!�ڭ��ZD��J�S��K��	�B�%��|X�gy��=*Ҭ ��0j�[p+�Y��A�"��B�TY�%�4  ��ꮺ�T L�4�V@�nf����g�?%���ܻ��R	#�B�@��LP�h�e˓�����'p}����Z���"���3z�� ���<����U�ĘP'��Vz�@<`<o"�؉���u�Jʳ�]��7q;.h���D-*3��5�0�mmH��܈F��b(�4/$���VJ���ʆ&��������Ů��\��7�\]�9G?�Q�곅�8Uv{��0;	-ց�jE$b�[q��$ݜ���W����p	j�/v6�O�����~�*��򂸊�M��h�ǇQsz"r���c��}yYN��?m{�;"�wo0��i 0 �Ij���L�	W��thf�=�.��ގ\��}�n{;�$;�+�O���"Ac�U��V�
����H��.вU���b�	��1�G���$�߈����K ����f]'�[��h�������V$[�K��xF�������+�;�iI�L�-�����?��K��e{sFʸ�.ӫ����I��!��P���RqKT���
�����{�H?O�w�.�8���/�?5�$��V�=�&w�:���4IW��:�!)␮w�y�8���&��50�9�����,"��ֶ;''k����!��2��YTAiH"��;{����_�د��/���"d��`ݬ@|��3��RK�(�%�[�)����j��J4Ā8��t!�n�{,�_�܎1��Y;�^ބߵX�я�����]��c�mX4R�W]�����L��ى�.�W��4��=�lp�
��>� ��5�����T�L�?z����f��}	O~�>>�����bubn�zE|,j(C)���K�:���s �Ѹ���O�U!��A7�;KNI�}y��f���F�5S���l�z����~M��� ������s ���ݣp��mB�W�?� � Ȯ%��Inw{%oû�i[KF3ك%gb����嫦�'�2��$?����l*�"� |H�W,�^�3��y���e�J��s')�<#�NLWo��*nD��pmE�0��������|nM�u.�TJWG����
j�z�'^2��s�yZ�RA�ͅF֧��M��(��󆔉� �}\���S��n{Z(N�8B0<���Q��\@����C�*C4����=�!̐��Ž��B�o�[������l}c�^ lU~�Mǘ�f�7���#��z���۲��<:��n�@�2�����<h�]]/�Q����	�-S?v)��쏾sB�:�HdH�$����N�D���A������62�Y�FK�����VI]�!B卆�1Ւ�j�Y#�B o���?|�3���ѭH{	�*ۉׁ�f}��Q��ч�9y!�y��Qv��B$�&|P�P��8v�;8�K��33awq�ۛp]����%/�41�'�)���>���A�L,�~a��ƺ�y�A�G&�Gkנ�l�y��5�"$Ғ�0��of P+��n{�Q �����x��;�ز-�=ma�6���Z3\�es�L:*��m�ݰ�I�eN豈�!��}F��^�We���*W�3N��6w���)r��E�Y`b��c}�Cӓ8��|ݩM���s�[�ŔG���.�cr��Rr1�� Ř&�9Ϻ���vd��ē?�~2ʍ�Aݱ�����=�b�n�z����mT��!��>5l���NO���C�-0^�E�Fq���?���F��&&�^��)	���]�F���N>�wR�Ƚ�&Y���{RH�Ǎ�{]�e������92�o����V���Ց#��?�0^�n;�6DZg	΍+�Z|���<����� W�6��9<;KX�kUO��?�d��%x0����Z�\q�<FA�K?��E�1�NW"��h	X�z���5h��f�O@��S��������UrM'�ƨo����7"�CY�7].N��G�8ٿ�'e�Lyz�]z�ފ/�W�<@q���1���&�څ�m��k^�q�3.�ؚE1c�A^#���ģg�לݓ�9�?m�a����rх(��E>7xA������@ik۳}��%L�P]��6���#d�o�K���")�/����������-ߕ�Ә�9ԋiq�4sar�I��t�ݚ������t�i������Ș =�|����1��< � =޻ m�5�R��P#�f����P&�A_�]� �`�ܕ��}��fH�t-g�?����W�d4����̶���^�^))��"!�/��]���G�T�_+�G��(jpK�^�)�.P��
|�ۈAx��u�}��Z��Q�.I�e
��ϐ8����JP�5���E;$,K�k���.J�����_\�G��CH�ǘ)���Y��=���k��4��!m8ۨ�vQi2T@�(��4�k!�b�`&���
G:���{Ѐ�F� xa�뱉~A����~�x�[�q�;����e$�ƈ�d�:_��S`�ڧ�fces�]:��ꋯ�(��؁� ���_\:+N����)P��w}~;c6�@^N[�ѯ�����v�Zb_�FC�]���uMN��.�������*_�H�
��'W��`�mؠO�H��d2Ǆl�EY��x2~�ex$�ݻF��	�'�T���,ݰ�����%�5�����u�5Ѥ�'Q6-P.�L�s�~��+p!TUPP��k�1
�,Ȇ#�B�wlٚK�A^�����V�unȦU�NY\V��H�=������'�M�j�НEr��!�kN왡��
c8������D���2��c�:i��K3H� !�]$IZ�����T��Fɢ;��2G��a"3���Zf���d�'�uR�~8���t��5�6���*E�']�{qܛs���4r�+y�]��t8���^�'�۸>��Lʟ��4�~:���z�D{.��j�='�(��
�
�F�j�z��0�(A������i�����q?�zl�+���A.�Q��}�Cء�Q(�V.l��B�Y�`_*���VD+�s8޺�.��bI?,4�_ή��!l����L�2�L0p2��e�X8϶<�|�6l}Z�&�6��|���X$N�J&u�b ((`4�2H��Z!�E?�/��� ̂���z;�g�����DMj&�?s��:��I�Uwf"Y!�}���E�O6�c���=�$U��K�/8�>%&�
J<�=	(�pȠ
y�-��ݮ=��n�8kЩ����ʉ^��H�O�PKK��VDao[���6W�P�C�Ztt�*O5U�W�(�C306}P���K�&�/Z�dn��a�/k�k�~f_��Ѧ�?����1C	�//�h��-��1���yR9r�K�#+�H��m*s?�
�V ��s4�N�pE�#���ǣ��2�!Z:�53m|b��w��,.CG͜�T7Rz�P�X=��RD����ND��CF���i�Ⱥ���t9ް]���3�%x�u�#�Θ�*s���X�dK�Q�z��˘�Y�v�����n*��ݻ9%Ӥ�KB3A�W�Ђ\-�L�/`�xJ���t�5�'�p]�j�k�p���lÿ�+��O�^#�	�X�]w�Ӡ
��a�@��HhE���įcsn���n��=�{��G�5A_X��枾�(3׎��]������tX��]�Q��7dʕp$�e�ـ�-$�MT8�fQ�:�{����������[�2��6o����h�#���Z�^��V �������D�gas�Ө�U	]�R��}����DvmH�ӱPԊ��媤��,S�[�G6�tQIx��^BL�6����H#��wtEDaZ�T�r$EY��o�UB��u���*f;��/��R�nb�vj�X���+��0 Z ���ƴa�wt龃rɄՏPa��2v��l��O�9����Sb|��\5��Df�)}7Ōb���x���u}p�Lv_��)H��<I�N���Vn�v���� �T����W?B�Pt�7�pP���
���)#�	n���tl4��M�������?�?�p}�X���E�X�Tg.�+2�
Qp�W>�?� �� �vR�$t9���f��"�Ĳ�'�ݮ3���?��h��Bw��N�%����Gٟ4�҈�w��ը�8!׊�LK���dF���$"/0G�R
�ֹ�P�Mj%��+4l�V�j6�%,A��י<�08lo�J��Th_+���%�ۼ�����Z���~���0�ˆ����M���ͅ����8��tn��z�|�.����ᴵ��T���%|��i���IK�[e��z:B�Sd�G�6\�7�'r���%��"b� TD뫢v��"o�_[��s�E<���!��ǝ�g��|x����ߴ*ҩ#,�'ч' �oVWl-n^_(�@2��@s�����hd�H*����pq�������
M�c�34����MC�!m�<+,�[�Sұ0[�Tc�����6*�*a�`�l�&�=�H��VH��-�'�̿I3/b�a�?1�^!��;OBl[ 3��2���5H�>�N�PZ;r5�<��� 7j����+OᲩC�*�,��=�B�FXr`\��[�	<x��(�M���Bb(C���D�]�6��M�h��@�	�:�nEӫԓ���P�&�dO��>��{��MWiVfɏ��oż��˓�&d܁>�Bm04k�H�3�3�M�)<��G����.4�V��� {A�-2���=b̸wZ��d3i ��������)��)���R��9<��C����­���o$�,G^����*��2)�{�������\�(u0��HK�=�%�7�E�b����E��3��̽ym����H$��p�+�� V��@�S�����Ce?���N��}��}LP�y���d��a~���V6>��l�Ǐظo[�,u�p�N��@���s�������=�$��Mq�5��r���m�r�d@ҩ�7p T:m;-�kP�6|�}�L�7�/QzgS����*p�A����[�������u�{��D#.T���jT'�n�+s�a��=����jl�pY,��D��ύ��T�!>�p��@Џ�����+>8�XK��mb�q�Q�8����$�N�p�$�����(U���Ԕk�&9��;m�;|k�JI4IсŮ�L�k�͓��N��mA�E�S�Z,S0Q9w�� m�1xo-��o��~�܌�4[�t��	:.Jj҃}��|������e��d�}�uG��FBT��b��e�fI�*A�����s�����I�C���h��L���_��>0
燂eX�p�$�ڟ��6������I=� �F3�A�㯇��)�����Kn����G��'��z�"GKX��6P�7C]��QӴud,�K�0a�<U����$Ik����7k5�	j�P�!�T{�i=�H�Ir��s�ܷ	 �q����^ّ���$"2�xI��
g�.|\�NS'��C�N�X�/��<Oy+6ʴ�{�i@q	!��u���VP���A� ׸�� 
�I�^�H;b�Du���m�A'?�����z=�6��9���̐?�� qx��Ս�������W��[�i��ϟ���T-�����ҙ�};��B����������(a/�����'���_�BK��<��N���4CW>Y�J7�4�^̭٠a��PL����%�e�W� �S���o.������dy�z�#�
G�Mt�(��3L�K��c;�Dn�N�e��|����!gԐ[�g�G?A*���pv��\�z~�T��,�(7���C�aN�ZZ�9�A�����b�d�u���U��Ȃr�667>1���j�2^mDtiY8q����^P��kI�H]X��W��1�[�03�.��$9�����;'�,�R鷗i��21�'b.��U��_�f���:������W��׾�	��?^_��OS�.�c�Đ�x�̴�:�;�-*��)Z���>��Jzn�������ڮ�w�HӸ�y�|��MʁWI��}룂M�'Y �vG��$S?`���<��~��-ÿ�'�?�OBy���7g�XY:O�)��O��5��5i�2��ȵ�s�\�^�c���Ph|�D� 1�~V�ڢu�u��q9���#>��STD��q-��D.@�b����Q�@@�~3��8�!1�p$�M�{n��	�B��sv�jU�ݕ�X�Z� �`����Z ��]������FX!:�B�����oITE�_/d��2�����|�s��8�m�@�%�y�J�z$�������o5ų$Ti��;q�=n��J^�G�.iC�w,�B�jL�9b?#��D�B\��
 ��J?�-��fc�T9�B��`q�+�'^3G�CA pn����I��+����=`�F��¼�q+�q-|��Į��ǖ�Y��=�t �iE^��Ap.�|	��o���
{�w���!� �h�A�h�*}}�Ӗ�7`��]�x�y�#� 7I����>�or������ X����[{1N D7���ǎ�@����&�<*%'�Ywy$��^[y�x�T�ȣ��w$�͘�r}=j�a �=R%��)��C�Y�K�$�O���[���:Z5�~��.�����x�6�x3v��BI���s$�j�>/��
�o�残���9Ha�m.�]�nXB)��;Wi�ƞ*������"���Q?ZC%;blW� V�:ـƼU廈�f�"̽��j�ǿ[D��*�вa�26�s3���_���Þ�$p��2A��~V�>\���>� ��Op��>�>E�U{��kȻY�5	�^1���eٚoCWy��D����8dP�Wz+��IK�P�ࢌ��1��&9����!AS=�-���|0J��*��g��F�����'����S�*�Eo-'��)D����7��~D~�t0F٣ƛ�r'&p��.�Ld��Z�*�D�R�i(pә�1��4�Ẋ�
mtM��L��A�&5����eo�x��;6�ƵxJ�I;e]ؔ5F�ڛ����?̓�D�@�r]�9xL3�W���cm����O�_�/l����-�
	��#1�"5uJ�-!���!e��B��s��-�/����l*�����@���5#��;\�ui���D]m���m=��	L�f��Rw��$%��E�E��,�d?E =w�s:���2ߪ�5紐�G�g>�&��Vd�qG��ѕ�?���T�:��G�֊݁��9N���@��	�Ǚ�2N=��F��ȀH�y� 'z?M;v�r��\�`j�'P�~<M`�[�MY��;��t{pO��&� ��L1'��
͊�`�f�tY� �"�w���t�π�F�,�䌖v֬,�l���=R�3�miX}V�>�P���gv�B��.���ٚ��'a��.8MWפGH,�S�g���`�Ȝ�P."�5R
@��
� v~s���ti��
�*Iw���a�M	T�G�f5����ڨ�WuB�R�a���Sy���-�}�*#�g[D^��*�6�{��L#f����ۗfyx�'�V��������?[�F9
�`;!!l��_Oj�{,^����Y+9/B�q2�4q�R"�����r ����u
.�bʞ�~ɧ���=��F����̮O�s>*8@8���T��^���.JɏW��+;/B��~l�+�'B�m1i�.�ł���0�_!Ƈ&�X�?3��u�58�/fN~��Ď(Ͼ���8�۽&��`���d�E^	�PD��rj9X�Ll�go-o7��0�����Ӄ��`v��֝Z��\��	��ֹ�wT�#:'QU�xjH��%7���e���yŌ'�ʬ\Uz�Um\���u��(2�ʬ/X��_M����t�tef����p��U-M�/��X�Lh�WR��2�(:�ՙo�Z�}㦅S�?$�(��\��
�[��Ӯ/�y`��cX=|(gLuF���gN��D&�*J�7p;ܞ۽m�P)�V��X��&�yD��&�DL�L�]!	����t��J��*��c47�au�0c�y�&�����ĸ��H����*n^<.ÓY�(Y��5�R?5���<S7�tX�B]	#�`&����Ǫ�48�7^��(�V��9���S�[��8���X�0���w�
�G`��0=<;��r�ZF�SM@Y*� ZwXڏ{�c]�j��Ͽ,E� _��;y p��(TY�E�h��y_��'w�%��?
$g��)��*�A��C�b)Kྖѱَk��v�B��X�������� u寡]i�"U�,�*?|�"�ӷ��^�Z�w+��c=��2��O���e��U��饋����hO��'�v7��KA��o<�
��P�4�>G�6�N�$;c��6=d�0����M	�����6�G���� F�8�-' U4�|�ɱ~c���������|AQ#����Y����PN0}p�8;��T1���
��)��s��!≂���#� ݇�y�b�k6�
���{P��S���#}ABE"�Z�_�����$^k|�6 <��v���!��z�����FO�!�`i,�L�9��f�;^�s�u�;�v|�x�[t8ݜ��!_W���+�h�U��; �Np	rb��������pcPKU��>M�Cn�|�_����5�ǀ��G�uQ�p=�z2�!`/R���a����s���M�-�UK��56n��p����\��o���$�s�Ʈn�$�㢔8�%�Dbֹ�9��p�q�[��J�BWR��I�:��F�Mʐ�t$bٳζc�Pj+\̪�X���S��`��t#yƊ6-��E=�J}�9©��)r�hX% i����Sh�Զ�)����:�Zİ1������01��4���s$ւ9���p6���_N���67�hjt�����R^mc��'�z�����$B
�j�D%q��;�S� L�N��a�/F�f�>� R�+ie�Wz��$�O�>�.��AHՓ�,��_���7R��{�+�!�s�r�����+�q��U,��N�c�U!��ڽ�L�H�����f9<e�������F��d�]mzDB�U�>�m򒆽�U�z����~᩿�v*�R(o=����q�q��7��w��1��8}S�J�d�nc���x|W������ D�'�l��`4B��������w�)k�v�[W��w�5p�8����HdC�����A�A���Eeh�῭����2�GS!uP��Kl�}�� .�ˎ�~6�m�D,�QlNZ�?���6���GmoV����R�9��һ�+c��Yh)űa����X�an��%HEZ�x�����6�;%�)hH�~�3�LG%�U�P�DB`%M�`��F�dlţ9���t���KRU\2`����_���Z@��@�j�H�w�y]�lw��8���kg�FП���d16���j���@��O&� ����(���a�Ƈ�,]̣�?��Z�rn�T�R�-է/�r]-*g�p�S5d�
1q���͋�@��͟��n�]N�-}☮�Y�(R�b�%������g�(��ȍ�nTb(&���b�c�-� x���(�`��ȯħݩ����T\SA%y�t�t�bC����W��,$�U~���;�3���R#������h���k����&zR��q�Pj��pT��_T��W
 �.�`�sD'w\X�K���ؕ��+Cu����$��"("�)�I���NZ3^�q�,z�1��~n�0�ƥ�j�h�x*��P�K*��X�+��4)��P%5��D�&�s(9�Ug��(��X���cj	�a_�Ū��������Z����e�v?�T�����܄�U�k���Et�ʤ�p��~*�h���\0�]o����s�<���,j�ce�j��=�N�k5k��ř�tG4~ �U	(D�uf8n� ]X^Հ$tq�/�E��^R���&2���AI�n~f;���6X�0�7ע�g����# ��H_6��+E��b����%��ɹM?i�.�Nm�]Ȟ%B?b����	��cE�}��UvrӸɘ�s��z���v�y�*�,e�;>�b�vVqZ���U�@=���˂�J�U���Ys��`�e �[!1K_���c{F`>�%��|�Ȫ�$�͛;��K�Ǯ�K��d��p%~�b��E n�P׉B�a�5��_	�|9.�t����ֻ�%���8:ji�1H�����T�W���:��������:��3E����$>��`o�U� ��H��4�О�eo�uBd�w$2v�\lz�E�������{����5�!������{5:��Ztgw�;P;S3Ep�H�8�����N�
�F�N�Up��J�0U'�K{�L9���V��̀�y�j������{�9����kTѧ?B�~*���2Ί�\�h_���r��1zyh�"H��+�/����ka�/ׅ]U���PM�^fP��q�����s�<)13�W�%А.�^��9���j����L,�3L� �%�e=��r��a���j�3��ޡMU)�H~��E�L偉
)�:�b��U����58&��I�V�I2�B�h�]�2�>����dZ�`%�@�[M�*,Yl���`�3�9J��׎~%ϡL��ifȿ&�W!�� :&�Y7�pچ��D �f��B|Ĺ���#+ʆԇQ�L�<>o`�Wv($���c?��WaZ��aᒒ$��C(�i~K�� �s�:;�S��l��,�㗉���D.� g��0oD\��ٿlũ�����QIjڴecH5�vh��4�#Zղ�sھR�f�ȶ$��ic��8�[Me�cQ@�X���p9��t�"U��8
~މ�z�D\`^N�d�a�xt5��G8N�1ʣN�+�.��6i����᪓��P���H�]=�y����rx�;���@�ؕb
�c�Zv��q�.1@�?�A�|����v01����\���z�	=18!9�����-���m���$F�"9�R���n���=���{�R�F���[A0�u�b���P���y}��/\��|؀�D,� ,�����,�S ��
�ml�n��D^��n��LW��V��6n����"�kjq��1�6����.V۩�¹d�9��x��8�Nֹ�Џ�֚|Gg)z���ޓyf����\�T�g�;�BV�gR�o��r�q��O�)��sނ���r\L�8/�3������LW��?�c�u�JW�m8?7��0:��
M��.;�L'Tvə���˒A�T��uS�Z��`�,�x�"M�e�i���m?�qF����5l~ ����2�]7���T��N�9���Y�Yڬ[2�3��D`T�l����L��1X��(��B���	���o���m&�Oy�9�"�P��$S]�`��85�Q���ݷ0x`�^>65?l�:�#�G�n8���%r����"�]銗!=_
�o�IM�ȱ-f{?�(�=�0��[PY!�%ȧ��wل򉸯)z��1T�J �'�nr4,����xh����:�"5����!M�<�0�U4�����4˒2�/ދǩ ���Ï��? ��aDL�fo��BU�ϙ-P��7��~ƈ b��e>��39;�g������&rQi@P�
&����e�Z�Ҭ��p�8(����TS��H��r�X���~P����t�Ұ����rc�t��@o��+S ��r�M���=pµ	��5�H�VYz7iʼe��2J�$�~������c�(��\;�
���a�O@Kk�(1�����8"D�G��_?�2�SI
r� S�ߺ���$��sVl���n�ɦ�L�i7���#VA��nkv�(��u�o;�K�����K��a=�r���/��_߈�]c`���#!�48���*4r�����I����̣@~�0�O�hv8�eP`:��2kVGʍjK@倫�����	��>o"aٽ�����k9���l�뷜o���v!:Tw|{��9��n�v�H,��H�&E�ƞ���*�Њ��8�x_��j�	q�$ ��1쟿.���7�x�V�CT��\���4��)�	`ќ���7����%�&r�F`s ���Y�J�([���E�g[�lL���ak����ڷ��Ƥ��[�mj՗�26]V,[Q�+�'��Z��U��Ϧ��0�K�RM��ϗ*��Z�����F�0]%8L��'��\ʓ-t]C�G� �ƠB%+
v)�O� �Q�,d�R3~��?�Y��`�^����������mc�G���Bb<�U���u|T�N�[Q���`4�$mhB����o��Ӯ�S�|c��_S�����ϖ��	��hZ1�����k�T�q"P���'����9����7o�����������?���$+s�}d��iƭ�*�E��g��ي�]R=l��6V�+v��qOO/��%�>�땬D"T.���I��"豱�!_ܜ[��ݟ�H�֖�m,_0e�ךPۄ�g `@��~3C��e�!�6�J(~G���
��|J`�����ƃ�qk&�Zg�md�٧��w"�Oų�������1)�����?qUp��3U�]Q]g��ͧšu�9��緉�j���l^u��[��f�x����Cf���	n��p�u��l�{a��AEג:5�aЕ9���%�b�la���+���#h��5"m�7���'�(
3\*u%�N���|@�_�`��C�	�Ea�0�mu��/�i�Q�x�t߾�w�B�4���� k���%6�
)� �����+[;TU��2�*�oY8�\6洐&�0�#�,%�X�͚T���,���-A�SD��78�&;�f���Y����U�]��݇�"y;�X�!?�g��n{��L]��bQ��!?He�>+&m�a ����K�����}@ʛ_9f�q:����_|�Y�����~ޢ����2Դ^��*᥿$t�*#e셮�Bj�!3����|Q�SF}XR0eG�g��[2�upp>�jB�=(��$<�������<Pq��P��jZn��z�°�#4�uC�1"S�[�j6�)Z>.~����F<Q"U��_�&{�7�ˣ���",�=���ᶋ������=H<�K�V!�h�����e7�h���Q�/eA�u>\�&�Y\dTΪ1�hzo$�gKv�7ī��ț/1�Lw#��w^62��kV!C.v0��*�8}|Erz��i�{!�٥�������`�产�Q��t�B�j�����y����âmU��@����߼���l�\�Խ��]V���։|�܆�o9T��ܣķ�G����� ���wzun:;��!m	�}LI�ji��}O�'tWȷ?!:������⌛�G����J�ia�m�r��uG��䌔R���x�PAr屹��1����k��!��ɸ�!\� f��/K�b[[�tԻJѠ���]�b��T5�l.t�ӫu9G��kn�HTPH�ע�^���[1Q Ud[E��_�lNX�
���P��>�����^���8K���+)HXZ1�)�s�݀�w����R��Hrr�=�Z�3��Ρ�r�����8���Ԃ�?���#j|�F���!s7b��rXRJn�����N�\	y: OE���T�0��$�"α�z�ߚ�S�kd(C�?w��*`]!�1��.�O�p�킜��������;�t3�J�9�7hN�^ �S���8 �5R'�r�q/��]v�͎ʋ��p�>t�Xu~��r��v��r,��܃���d:"X< �,!}���-��K��[DKXf�*��||�	���Y�+ �齜�y��%2k�-��r�	j͘{���m?D���� ?���	R߸���_��Hf�Ɇ���@O�k�f��j�ߦ � ��V�;^�)�Gd }1�]\u���J�N׶�%:���r�X�I1�4��_^�� �,8mw�R�5{��x���.K���zDG��p3�;���b���D���C�u�z�-��4c�a�Yv^P���_����/F�jrr�����a����x%���e��|�޺����-e4���/���nٯ�NFx?Q�<�;��&>�U>����ql4�Etx-��Wy�R�/���B���(���ϦL}���Y��T'��D5va	F9 ��YuvX8/`\���ϤfSM{;�-��)��mdc�{�ZF�J��E�$ǽ���M ���hq���v�c��,;2L�y���P��X~1@���Pw�$]�>N~"�ޑ��ӉL\&L����G��9�~=�(�D�'� 47�L��d�M�0.��z+�,^� �[(]缑��o��
��-y�E�t��m���&�Krk��y�c����4,���zL����Bǭ<b	H��Җq��j֐�>2J�5�͗�y���l[��O�`:O���$;q_e�O��{�z��!K����������_�?BZd�^2:��N;y
��\Zf#!(�,f'��<��r2O�� �����UFa�$ri�.bY4����=�q�k_;La �.O؋��op6_�]`�9f��9:�H\��&�����=y�(���K�D�q�Ȗ�n�Q�bwP���cƾ�a�K���߃����p<�b�5�{�mk��X���=d���.k��C�T~�R���"\r��!����s[H�ʟ/zM�c@���h���O���u��q4�z�7��R%O��"9�>�^]_�b��.VWJ)8,�>�]|Rt�UP�94?����w�����1��]2���p�35�gB\�fM�����O�?<�p~gi�� ����D���wj�t}��]�_gu�]&��9e�\���%���,<�v��Pwk�.����*��0cuj:ѥ{ߥ��yc[w�>�ҏ��mG,J͉����=�P��i����OxU�C	<'��4#J/3���e��r�/Oq �б��h$�1'x��J6���X�Ȱ�M�I����Ǫ���Z/��j �>/ךkG<�}*lO���5"�_�S{��G�cvf�H��y��VR��p����"��n���!9�p(�= ��u����n���چ�4 ��
��i�Bյ�)�P�5���p��*��t�u��7�9�48_�S�OI! |w2:aQ��G��Ga�j�T�]�+i�^$*U��9��ˠ^���-6�ٯ#?C���������4m%Ag~����6�\h]�i�TN�9�)�PWQ@m`��i.��9�/��tl�WC�3�Q�U��M��*��~� �@�C�>��[q�"sY!s�G����U�4����4׭Dנ01P����29��1�J�`�7 r����I�s���
�x���+O7�0e`�e��9�˻/I��ȹ@��t�%n��s=r�����v����HX��O�ɀ��`m��'�����{1�8,2ipb�<V�݋-�\l=�{$L��vz4$$�Y�<sղ��\6�i>��#�^�l�<����Wc����!�B�_�$60'c;[�%ǀ�:�}�=-ުX����o���w{0U=���j��#�F����
h	�8pҏ��8�����L��Z��X]��*r��?��^L�۔�F�l��_[���6��?{�q��7\�۞�Rr41!'��\�غ�o4�����w <r�C�SA��� �6D�
�U�*�
�YU��;~�m�����l���.F'�;�f��
��\%��83�����E+8�Ɣ�#��D���]QvO�g�K��4\������9�8tH����!�V\�S�5V�w�0}�R��KA|.����g�QE����?��MlBYp��Hj|XBJ�Q�
K�z��9�`�n$�b��f]��87�cҥ�H��6�0�R�<[k�ʂ��"�N'����O�*��%��Y�)��Țln
�z�HR߬yYUTbz�hc=Ͼ���'Cf�w���[�o��`\�xWcyP��W��q5p����SC�֧�:1������j���d�[�r�7�z/�F?t�`�=�G�/$"4f!��VMA��H�5�11�x���܌�t��p��-�!��4y���V�[ˍ���Gsax��;%u��J������m�Y�;��2��X .D��<2�Y���";�s"AMG�/$��e�~놏�_��*tHM��l�G˕W��G����w8TyXAq~kHf��Z?#{TO�tcG|
�sž�S��$���B�K#�*n��-�?dF�D����Q7����Ȯ]�s"���(H���2	�q_���[��)�]s|�������2c�@9��C����"⯆�v"Q��_YB�u����ty��IF:�=�S�*��W��%+��&������8b��ifJ 3�l��`�����YS�Q���#שL��f�^���8Y&�G�s{�-��_�=w���
��= �k�ì#5���S���n�QkF��G�`P�y��(�)�t��*��:���aenY6�Ɗ)�Y�A/;x�	���7�7�B��x{?�s�r�ђ��N�b�%�|� ���&����T�9F�jb��F��L�Hԉ�6z4؍c~|��A*S(wcW'���2a��(N��g�(��kg���y�u�1��j6�E��#�DNrN޺�@t���f<zi?��i�M��@��UyWjTn�����z�r�O���)���9��Q�T>�Í�ͪ�=Ǵ��9�l�|�+�6}��N�KX�����Q�#�|
ڧ����p�}���r�� >m�~��u4�2kG�[U��f�ᰚjTޔ�*]��[e��/G (�u��
�9���5�cO�W��A�������&uy�����EC�̪?T�q�C\U���9���Z�ͦ�S��g�j�%��/�]�+�eX.�ê�-M8�T��h!��l�F���JL�lu����&���=���n�^TS�*w��=U�� ։<��yK�.=̞�1WyŹU�`��Z�M?/�z�0I�:�9��8��k�k�E�-�3�b?\i�[��$����ck��k�'�,8�+Ȥ���!���$˙���%'�4q����n3k�����v%��+�������o�Q��<u�y9t��t����e���ZQm:n�H �(��T'ac��Y�μ!�u���
�������h1RX�*{w�_"Q�8���;�|7i����K���Z�F[��є�ˑ�WQ��ǽBD,�;���B '��LY�H�V �q��Q�q�:��E[�K����������鞬��h�,�_���/����4u\�{��L s�3��<t��.3MlU݁N�� ]H}�Z��#��V�
<��JT�1�LK�2϶� M]$�\gI�YL���CK�;��U5<����G�0+T'&��$���8z�_2���r�<=1�J-�%���l��F+�Mw4�S�(�ӫZ�ncj2�´Q7�H���,'X|�]�� Ɍ@Bߝ�AD��:��؟�|�����h�b��m�ew䈸�����O�$ifu�]��3u�zs�]9�C���rqRF�v��i��	e�h�H�/�b�A����96���2�+`��0kx�^���Bo;Rw�m�o	I�u�,��OÑr�}F�?V뒭��x�Ul�g��fl)��$A�ƌ�z/q�?��Kv	L���!�M�6��tW�u�����
��h5��@M!�	L�h�Z7���m!�e�同�H��2|^v� `�
P/d�d����i���P=ܦ��j24�i�j	�z4�h��.7���*u�J�uQٔE���K��2�d�R�1����[�8�J'��E����c�A�'��?
���&�	�"�Q
��y���#���ǖty��W���aK��)6��n]r�ͻ��B$��F�mҝԇ��.?��pU�#��zѡ��MM�A����v7�Gќ���0
/ -`, ��g@c١���~���Kn��L���ns+����6�����qG������L�y��`��wK��GIĭ��㧝�%�BN��%�1b��#9�o������)�[A����L���ɖ�;w �;P���d�e��eJ�9�2��2�;Q�� L�-y�ǖ@�I!�wךU��?A�{�"�z���P����u�q���g��wكG|��q��1Þ9�u&y���q�e�ҥ���d}1v�e�ɱ�[=�C?7Cf��5���4�C���X�ܼ%
�4)k be�r����k�T,�}��_�·V���~bjۘ�oz\b�A�m5)�{'�ݖ�*Җ��W� )�-�ܾkG�q�չ�q;Fe��R���d(�ۡyP%o�/�('W�2��G�V��"��Rk��J�eW,"μȇx���L{�,f��?�;	�W��J�⊦ ���h65��^hV�o�^O����Vb�a2�xU�0MYu�q��,C�z!E�v�\�N��Kن�9x�Ћ�H�ɯyaM��U�͝!�ԇ�M7�	���X1�Ԯ�hkt�<�1�>	WM���mg��iI��,i���w/>�h׫��`-�T>Th�p�,�"A o��Q8��I��k�I�(�Ե�ƥ�'�X���P�Oa2�&��UMx)��2���|����L�H�Uz��B���� $��Ջ�'c�8G5�_�8�O��c,֙����K �"˦��U��Ñ���������}����g��������"?u��B*dD9��P������j��GwU�Ỿ���0����'���+��+t&^'C�S~=�LŒs�q4L��brF��U×�u�1�
 ��]N�h	�����D7,|I���K:��v煢���%��v�gT��/q�ᱹ��+��My��fiB�t�(55�\6�r������pu���\�����z>Ly�w�g�N6?���T�����C]|�/���J�����:��ȼ��a�b����I��=Y��o�%�x��ȵ/"`ҮR4���p�H��xH8�HDQ�V�Jě���®�xn,��3���c�ٌs��)l6�5�Õ ���\.s�S��a�p�Sqj���Fbsﾵ|�|`2����|�T�ƫ��ͻ�q�oT��
�/aafI�V� �Y� I��7[r%�̢ϒa�4�ir}��аw�&��Խ�xq)�w�b�ha�u5�����"�g6L"#z�]b����R?S+f���$�������&��S�
�\-m�|c��"�2'\�oT22��K�G0�*I��c�	5\`���o���[��m��wDva��((�}��>�,xq[)��^�*�P͊�i$@�j�t,FR�������k��UY��ڗ��#n��]������1�9r[3��ƇЂ���bT[1�8�y��nF�)�����y&�	m�V���]d���>_ Ψ��f�0%�$0�M7�@Ӄ�@N&]O��y���r�#��<����e�Jk�.�c
�����񽌐��)�H3����v\�w,V�5�P��S@ϲ w��^v�a{H9���v�j~�K}�Ë�q�#��V���qB1�����Nn��InN�;_QH���̼�Q<��̩?ܲ ���sB��.���}[��t����V���xx@�I.�=S�K����.;�K��t�\.=!x����v�㰁�n����-qmWx5<٫o{�k-p�C�����]��C�#+�:�F��Ktovm�ˡ��>g��څ;���&��trUr90]���C.����U�w.��N4.�v��*�z���w�����͞�q�e��f �o}�q'&F��_��J��S��6Z�P���.l( ��#��x��OOi��9�!���p�M��/��Ѳ]u'���l��K;����d&rF�Ǭ�Cz���߶�����*��Z��7j!0)r	�࿄�	�H_�o,���$l���o�.�OT�+���mM�eE�v]���H�����4T��bBG���
k 腮*�����^�q8l'��:?7�^?~Zj���M�Dj�פ-��!�a����i5�9����9F����@��j�kl�hͦЋh��\�#����Y4�C6?g1�'%��ߑr=g N�Sg3,�P%I�c����ك�l�b=�J-�\U�=�j� *���[.� ��2_!��C%�3�m��Iz
�B�߸�n���ޗ����r�^-
�?�_�d�Q���t�<]n`���|q[d�G';��|�E��>=��{�o�U�0�@����B�tbZ���,-/��.�/���-pn�5���k��b�����rB�|a_hDs�?l�'0�[�ߘ���Ɋ8
]��*��۫��~(���ZxB�g�V=��}��8�~��s�r�S�4�ׄ���U�T�eD&{�:��~���ϒ�w˶W"WB{�N�l��3}<�K��-v�RD!������@���P㲯�Z��;+���vB��MvܤK�:��.���� w�N@�#�֍�>փtܽ�[�VU&]�\����4��3n�y�D�v���s�hSzғܼuDE�[ ���(���{��p�u�y�I�V�K0��v3�H��L��8�Ĉ�Qzܠf
��L��a6���_�HX�̬'�K�C�����
�0;vu+8*�^�	�z�,L�"�O�8Ǘ�_��J�{M��t7�7\�w�<G�gy�p�MA�Obֿv(L��ۊ�%��2-������UP�
��9x���Ѫ!f��-���T��@[gu��Oz21���~a��*�\�F~y=N�֏��h��Nϭ��#�>��k����y���^4y�''��ȣ�,� ��9#�	j�HdⱮ �

��9]ω@`�޼	����6���'L�s�KW%�~ZC�2��%\��x�ƅ&�q������[���{�1Y�{t����6�{�W;���Ƌ𬥧v��B�����(G�����kP��;����a�KrWn9U$��nPJ��S���
'�f�Y�7^�t6�U�Wr����w�E�N��,ST�B_�Q]��f�,H�����3��ܤ����b^�"�_� ���݁�9[�BK4+�鹂,X�����à#�����;	�m�]��W�Re�D[�w��(�3>فz�"_��̉��v��f櫲�ԛ��	���!�Ѡ�$�}�gv��Q����'�,���?pd�|�YV�I3xI|�+�E���>g-��#<��Ox�R��(��bD�3)z8�A�N�N���"V�S:Q^��av��PV)U�k��%t��[Rʗ%�����:��7Ͻu��)�w]��	1.,�w������d���xtR��vo���Wx	6Ŏ��k�yG�=��jW̾�H��W_�-�"t�%�}=	�^&�w5���B��P�
^u0��X���3��#	X�
۷�|�zz�$\��u0:;���lY$�z�ؼ3�q�<��:D7�V�X]�3� � �f_��)\��b���A�&J��&�y]���kcC��]B���Ϣ�r��i�itOlӄ]
m�Ѐ��A~y�Ob�"���т-��Sor�ǰ<���CR�o�ʏ>i<�-�I�8�y�y��sޮ���%��ߑ`ξ�tcפ?�~���CDH�u&��v����J��0`�t��2H�-7�1�������Y���6�2��t!gm+�)k[;c��os�������%:��I�H��kY�*�����EAX|$IL��xĄ����;F{�������z�����xB_VW4\ ?�*�����KxT�R��zk3��G�j)AM�: ���ᔽ�9e�n���l�3u��P��łڲ;1��q���^���a�}X�9��K!RS��j�L��G"��P����Ġ+��{<�q�����q�gl� ��O���Hc��%���%�̣�'�XiL��l�J��D�[W�J2�6��d�k;7)�F�t�ː���5�l� 4�y�QZo"nRy�P8{M�A4�����H��&���������������n��^����٢���>ƥ �'7ЊU,��(T�>��m��/Y�6�.��O�1�@衝D��nTWOP�4�����l'�����g���a���;^�ڧ��� T+(/�FJE���p���fqT|f>A� ])Z+Y�����nu�@����웶	n�:�C���jI��z�v �(�s���M5�{�����xQ�u!g8�*/s���J�j�i�"C���৔XI�W�)2��._ں��bq߼�J%�Q��i(U�N�
������`Q��؛]��g+	9�ެQ�'4ׅD-q�m^��L���� �Q������@�G�2J�ޭ�$0����yI�b(��q��ּ\�]X�A�I\�%<zZ�!�����Y��;V�X�GҲ�(a�b}�[���:�r�	Y����*�-�u-h�Fwһ��rD)��u trL	���՗}.�	N�'s@�̝��m���2e|\����m��6E>[M���f~���l�>�sd^�%��>�	��e���~]*Ϫǔg�#�jTXiW�j�V��P��t�i�ށ~r�͍�Nx(W˯#ƫ�����um�4����l����?���MOnx�;����%���k�+����r먃��f��.҄��4�W$;��}a�T�I�C�ı���a���8����M�8܏C}?�wE�����w�ҫ����ۨ߾Y�r���ɖE�B��4zv
��T���5�C���1v����i��>���!���	�U-�p�k��r�>&-��Ď�����B0mu�;��� V�<��@�Ļ��C.)g���4(���h/o���Ē��u:��y�@eL��+����M����ա�$�������_���_<��|
�O�6�K���W��Q�R"�%ؕ����"�Ӈ�[g~n��e2uܮj��!�˳U�����O7enm��~�_��F3�� V�YΡ}1���5��܊����	T�~���Ut��_�]D3���ᯋ�C;��7�u<��ٍ�7]��X��+�,��F�/�-����T7�¤f��(r^Lt��yv���/đ;����؜\&�J2�i�(�|+�/����zN���$�X��<��O��f��^��Y)��#DA�%�������:H���40Ֆ�V+h�:�ifZ[�����o�^t�TU�,Kv�̀Z�L4���;�Or���_>h��i{>|)�#V3����V�ͥ@��1L\�+t�Hw001�}U�����%�,,Verԇnd=�?�n��֏yy�;���{����w�n���v��|p�1x���I�D���g��cZ�K�a��|��ڙ7ǅ����ǈ)�F#բ]��f���b+jk?Ǯ����$|��L��p�gD��5�`<YA���"�¼�x�&�����d���#���,4���Y-*0�X;�޶�Vˍ	���ˊ��_�AԄХ�=�Đ_L�u�_�+�]çE*��	��x�Q�=��H[�>*@�7�u4
BJ��x�!٬�Xǥ��w���"�h����+�-�z��-���ZE�kR�Ym8S$H��G�n�O���j��z�5������gL�%��� �y��������F���I/=dơ 3��`��9��0>֭FC��=�,@�g����-pb4����|�9�Jdh�#i2����.l����,���I�.�����݈������1?���(`��xO눇L����	�V�̌xXƗ�,�ILa<G���F��>h|����+��	*��£�Z��3IY�Ꙁg�h��G\�QCf,|*�+�o|q�^˶�|���}M�f��$�Gc�&-�X��?�%I������+M��@�M�4���,(E�k8xL.C �
�o_[3�F�Sdu��#!�C�55Dް������:�'���X��)�u���`DU�Rx3�և�vCs�AU��6�Y8��{���oBR
3�B�Z9A�W�"T%Uϲ�Z�@<�w����r���NS��£�
���f�BT�X4R��BSX���i���
���mx���(�,%i�m�GG��������SAcI��Um>{̀��eL2&��0�-��RQ����Z��V�Y���S8���ݱ@��Xc�r�!�ά&��t!7?kho�&|Mq��]	g��aq�R���%kۊ��lމ���L��&��[p�O/��ӏ��颁7��<�ם����D3��|�������B+��:�5�7T��N��@of�!z��D'�Ǆ)�C液,�}At�{�#3�FMS�Q��Xy��0��Ү�>�W<;̩\z_~.�4ٕ�"��y ^�Ʈ���m#���������
���.�77�@E���`����ѪE���������ذ
�܄�ɵ�(���7�姥%5�����Q��x��l����5��bس[+���K{��)�-Q S��z�C�匄Au�K���#&��E�G�w��u�m1K9��IL��۪�Li�T�.�Rǆ|�,V��]��c����{��X���_j�����'�$b,P�|b��
y������3Q$P
�[�s7C�F��3:�d���dh\�K��ﮖ(�@^��������9���o����ȄK>�z�+���K��_x���6�'lr|�ȣaSmn����洵�@��Z^�@!���p�^���6|4g�������qQ�����Z���q��шX����Y��d(�ۓ��ڗZ'J�J�
�h��]��t_P�WzD�n�5,z��4<�SN���E�jSk�.`�!ώ�g� }1��oN�n�_�&-'�J#'�$��*�c��ۊqh�8@\�M�p�F�U��B��V�J�$j$ �I�$cg�;���I��$�הD�&S�xn�m}�Y��O�I65�*"�?f���v��͘BpX.x��e<(���7�ղ��YmIe��q_$�")��`��lqt�ͳ���k�`�|�\A��4m�KW�ԏ~��	{�$�s%+�<ʬA-x�P�ˉ�!���eww3��O���tL=�������j$+n\�ب`�L2�B� ��wP{<d��d����<�pQk_ �RY�S���%)d��+Nu@J5r�?���Cu��Q(�.�&��R9�r��TX��q���@����H����&ةI�\[\S�͌���5<�r,��{�^������@;^�`ǰ�F���T:��)6�$���h��᪴�U��l�{��ћV%#���s����R�es�r=2��O�8���,:O�4�٭���s�-�@���t�sC��ap$��[o�3�Y'4;9%�b���o��!��qh �b���b���X7o��Z�RK *
zaO
����X�z���!/4�;m��f�$�@iY������n<_�������k�l];��)�?��=�?p��D��������;�j8�pE T��Z0�����j��],,��g��]����gꢼǔ~8
����'Ky"�7l�2x��l^����֊��b#�ֿtχ��蝞U���VS���og�������� �%�~iTb?�J[X���s�3��|�x��+�`yH��E�#�2hd���4(��,D�fO��V��5.�@�G��E���=�@FdZ�F:
Lד�F�%c��̍��Mu�i`�.���f~�T�F��|��ޔZ9�u��~�]���.�l��.we�!`%4���������;ؔ�/�-M�L�4�:z-�5��k�cX�-�]�j}�g-%��C�_sǗ��E�|&���)��,<p���D6E�*-H����C���N���ZZ�@�`e�2sl�/�r�{��:29�-:&`�r�ط���O�+:Z {��D�G;�q��Sm���,��2M�,N
��R����Z�Q���}�i��J*A����O2�F�G����ª�X�o�M|�����Ì���H�]9�Ĕi�O�����@>���b�U�%�+b"�hs�=/��l�2�y��V�;L&Xew��t)QFg7NA#� ��������Ó3���_�����J�fQ@�T�5-��� ���4��4�뫶�!�g���T��TE���ڿ��}��ϟ��QV� X��\9w���;UQ.>r�GL���_g�Rw}�ϼUv{a�P�Y\�JI+���"�8�9�����ҟ�'P��i`��s�H�qiK�Pn�d5D/���5�ɚ���x�* `�5�l�ӡ0��H�N�)8��O�c[T�e���6�sY�M��@��.ξ{�V��� |eV�i�hD����SA<���^z��&
ǅz� �4�땐��8r��7���N�@ć�z����O�|C��)#��sO��t�
vT������������Չ�Or�Z,��m�y���T<�@�99~�*�HG�@\YnM������c��l6F�t����5��s��K�U8���~�LLl�NÄ]`U�����5
�9_�t�G1g%x�#��g�Xh�;��ۀ�m���5��*��{&�ArWr~��{؆��Q���&�C��v���S�eS�T���G�O���'�5Y7��,O�����r�/���Sz.	��B�mՖ�
%�]��/�ot�$�s��?!��9T�͉��Qn�6���Kn����:�A���)&���Ē�L9��Z,������l1�\]������1=����w�OD2�c:/�$�����Ujnzb��*�Z���5ti��3tL��$�?�U7��������·x�^��i�[�E�T�31 o�t	f��9�m-�����'������G2�3���<���������Q��ԫ�
"~�a?��6N���܌_��1�q��$I�*�bM�w�N�s�@�"`jN.��8<����D����[�{qA�K�y�Q-3��7�jm,�������=)�:��� ��bu�ou��ԧ]C���n1(������@�:5L@��s�����o?����S<��L=�n:Cf+��!�UWI�W�q���s�k�6���X�n��<E��,�6������!-Avܭ6��N�r2�������^Vֲ�rE���Zv�r��6o�L=ha*�0����ތ�&i�DۖD�$"Αj�ܑ�8�����R�T'��H�81o�1E��)
���I���^RL{�AX}m���O^�9�r ��\I���!�,Z���T`h�9s��0=�M8�5&��	�!پc�}�v�a��gbix�:D��� �sB4:�Y��j�Q�g��T0`x���Q��Ǧ ���mkV.t�O�_���&�FX�D��r�C���h�5_J�Vgq�SVu�i��_=�x�
|��z6vc;7[-͛��S����1m~9U�q۶��,�R?�+����!�B3�d�(��	����ű���Js�t�\��*�(>"[�6����",Oˇ^~�x~X6��/y[֒�n��_쐦^"oD!x��L�8(Î�Y?iM�����h�p���k����;��r<���	
���G��`/���`�U��0o�l�;'
ş��h�7#�%�@��#t��-,� C����o���F�,P�X]L�4�^���[6� X=�G=�i۴Pw](q�i�,td�7#E�"�x��<�J�O�(�3S�D�������Q�J���J#�i�1��$�f�=lp��8N[��_.L�;� �aå�.�5+���ք92s�Z֯��0�a\{�
[�{)�&��ok �� �ᮠt�?��8��^BT)Բ�D`���z�.�Y�Jc�.�?�I�s<����):�]k���AF�w&ƃ��I3q�#JZ�6��e��$z����E�J�YiQ�爧��-:�����X���,�w�e��׌�Z�ܜƹ+���Vp������ܼ13��O���t��:V�������LU^����A�o�F�����Rn�[�mD�Q��r�S��H=%,<�iS���sp�䆭�����r��k�|.7����Lm�������~�?�i�0���x���* ���j���l�w��e��S�6W�?��G~�XQ6hd�����e�Q�]c��3Sg��o�@�T01���ę�lV�Q� �t�$2:����vŮ����������!o{����4�=���ˍSD��A��`�J�DlO�uSE��0�+� �(��<r�B�I c,�%�F�}�Z��'����T�c� |�a�?����+���1����2 �n�bG�ر��)�ei��Ͱ�Y�/�ůEZ��U6�������v�vײQ��&�R�	T�֫Fr����h�>�D�����H���ɦ~I#������v�<�+V���Fw�ۚ9�A��ޯ/�%NU�R'Ӭ�����c�:�mV����k0�]u�\�S�*oiU��@%S?|�,��ۥ��`#lzF¬���y���<A:����'���
m���碝�3�s߫�w���M��0<fq��܄��Go��[NM(6�W_�o���d�JJ+����qw[�L�hQ�Fɗ��qG������%N.����:z(jv!X��F9�q��K(!u�j��C��:���PNi8�
����_�U�)���.�.@�5��;����ƃ>R5��P��O�0Bߖ��#�ɗ��ɫ�2i�����0�U�幺=ۺ�/��B[��3f7<�m'o���z��RŨ��>�亮��^�G��zӕ�!��f�/c�[�U3����ֿ����!݉4:s�d'��U�K����ue?�$6,����|&��}D��^ނbGu[$LH9��Ȗ���Ti������X>�O,��ԣ6�'co��T� ʑ�,*��i��N�r>V4dCv�+��?1�[O�3n.���
�Yt��y�Y�t&~c��S
�x��6g~?�M�����o2R}2��8)qu�!8���v^�5`�u6ŀ��o>�Xm��vV���v λ�xdn�ҿ[����k�rn&FC�&�O����_����н0PV?��LLwze����y���r�\���G?��-�N]��B��O��	�i��Ej���=�4j�P��A;���-x8����<u��c	o���C�G��
/h2{Ʊ�,T��_<��j2���Z� �Mb�[M5��>���Δ�����n%|��Ʌ����c�OP+�"�L/̩b��<�p�g ߖ�i����();��P~K:�/�7;�X~��@�r�7��u���qe�=v#���0��P�j� �F�hK�}ޱ��x$q�Ԁ�.j�A���1\�߸�\sDMu(ԊԔ�ڮ�9Ge�Y��aKZ�:���8���~][����yU��;���m�h}ҁ��l�^T2���r�B8 �8f�U5��.��(����I��߯�ڭ9u�e~J��V�ԕQ䵭�F��˰�g^�4r�	��� �]RY�O�K���C0��W���E�1��\����=Μ�A5"�J��Am�#��H:�5j!؇3"_���݆�߇ؾN�V���a:�����e�P��FE�9����f���_=�z�\{�+���J�0�X��K3�I=N��@F�󮞐��ϕ,�Ϫsc7�hw�Z !j4~0��K�	6�����RC_��q �xt�]rW��X�-0��<�X�֚]�,����<�����4�Pe�B������� �͛S�IN�\��4��E~��/i3���]�z%ju�2�5��wD�_b��ش���yC�Z,'.$��9��c���1?^��)ozc�M��F�� �L�H(����|~%���5���Tk�V���kH���t� ��=�#.�=]�~���f���>�	�1>� �lT�O��n�}��%l�-�D����{��Cd����B�y�K����^
�G!���W��jBi���G�_����9�q�w(�s'K��;B���ŷ�����y�n4,����na�I xn�(���u�Ĉ�{T�*���D��7�K��}*��˱S�q�:�^�z�T8���\�8-$��	OѦ��I��{#K���]�!�?�^��c��RL.�˲SW�.Tu�S0�|hH�ڙ�Oȣ�H �ܝ�\r��d�Fo���a�� ��}�kJW�Rm3{Zc���?0`���s�5�����ZH͘w�n#�I��h�i�P��k���r�A�(�;��������9�Y�϶N>���yO�"��?Ɔ%UǢ�M+K�I�&���5���$�M"0R��u��ё�f�n��~��P�"~�"҈Z`Z�,���U����
v%��{)�����e��C��5��[$oBS`01�����cVKK��V��� n�*�τ��Ϛ2�ƊPo��T=�1�ѿ���qM�6�k`���l;0��dn�2/���18@����xs�43�	�m.����-��e���=���#�k���r��2����i�ifEl=�`UPr�LRdSGE�ı�)��g�<FZ��۪^�O"�oY�7�7�����Xv%�C�s�ZWl`��n���`�R'�/�a�R���2Т}^��L������fȗ��M�f�&�'�:���&�4�����W�ES��mL�&���2�Mн%�w�xmi'�텱ڹ���ֹN�P��y�Wd���݇O���!@��!!�����gJ�Tc��,Q�9��v�pf(��Z]bt��l�o�?,:���ꖘ�M��O��{�b]�9|������&ܠ��?�L��Y΅�AVֆ<h�\����Q��B7Yh�c�d�cڟ�?\xf}���W���;Ƃ�?^�&��
�@{b��R��|C?r(0c;�$_#E:Sl]�*����T,H���:����J|xx6�ύ��B��(�.aӑ,4�k�m���\Y�g�_)�(����5�z�FwhY�����3����A��%�aJ;�D�0��N��>��<�W��'��㻣5���6�%�H9`���	������uxaI�H�g��H7��)8��yk!+��A�vw�Jᇹ���ʕW��.�I��i\��O��"����B��W�4�L��e��v�v�Y亇��EW���l��.�;�r�#eg߿�1o���NP�\`�V}V��A(��r����nG{N��霄����Ya�+�[�EQt�J�O�;��ђx��2�%�T�_��^�;f[_�Mn���OE��J7��z��N�G��$��� ���@������y�f���N�.��$8����W}ld�԰�f�K��a��(r�d<ȯ�X�@��-]�n�s�y:'��
ٵ�l�8��D,n�o3�V�O����/�GiEWǪG��p�hX_̈́K�SТ�@n�\���~�1�Tw�N����m��fm~�ǟ�S�t4V� \��6������d}ʌ��
c��*bK8߃a�?��Q�6J.�hh��O���U�ʻ��4�7�L9�l��'�RU�"4<���,#Ҧ��9��n�/e���zt�k�n��	%�1��L38��]���Qg�q{z �-�i+Wj�`iQ z����Q�����*�����w:��n��T�4Ռ�����@�JRhp�g��A���ғi��-�����>��Xo+0j<�ڤ�OO�ZJ��ui�q,ݳ?o>����}@�:�S듔��<��=8���$\˗�ݐ���z2=�`Q�,��]���۾�t���t1^X��O Q᲋�~.0���I"~�ڰt#1���.k��LC6�/���5��z��!�"����-�N���d��@�я�1Co��;�is��`��zE=%^�ZN�|����s�,e�hJ4g��T5s�g�Z��#}�
�_F�B���߾��.,����_�F���/�?tW����q�]p�F��H�.�C�l��,wЋe�̯�˱�o�f ��E �cyퟜ�c�k�~dm�HɋR�b���f*��o%e�������A�V�Ť�㒩NͧJ�m�n��*����zc����U돳�^�4��ը�ō�-�(����"|. ���d�ϣa�.�|�\�E�b�ʒW�)/��ZV]�x�e���}k����7��	_&�q�Zi���/����0w븓���<8��-.�s8
3�K�"��!G��'�S�:о\_ט!�2�"ޣT����S$7�$5�Q�=%@��>�N:��@H;N�}w��J��F���U��Ք��k�D�R�kJ~�p�ٲx���;L�|��jq=o9̬����\8.@����ۃ�m�,��ۨY����.v�cv���r���Ցx�hW�'b[LQ0��BM��&#2N�7��N�cu߉.�N�V�_u#�vv{
Kdsd.;��8KyZ*���3
-��<��d�΃�I2 �d[�n������tb[w��I���ɂ%�ȎK����Ec��-�w��L��_�s/�v_��f��Ŋx�� W�� �q�=����-�`a�#T:����.����V�`Jā��zf���d���_5x��>���{�w����u~�'�"��TΕ�4�0���22�,����'���O��Md�!x�%��QX�?��T���aI����5k�|�-��S��파��cjuОm�{AÉ��H�̼r��1sүTu�.l��ߢ�E��J���������'�>b@歓�n=��}�r�` ��Ӿ�A��w?�'XW�n�n�X�

AK%���.��fX<�j��/��7���x���j�[�Hb���K�2�e��������wpL�	�+C�e�����g{oV8u���'�/:u��h�Wd�D���ȟD���h�P��m���P����,fop�x�m1����_U��bU{��`sY����g�X�2~�wy�V[­��ifg����.���F>���1ߥNG"�zq����+�L��b뗉�䅏�Cz������&�i�l�ȴ�T�J�kֵ2�zc�XD�8ة�'*����?�k�6�ܺ��n�{jy��c2�>�$�-��rO�d�	I�M����p�8_8��ʴK�
g}��������&fh�w��x�Fi�C0�7m��t�#βo�#
$x�[S���3��A%�h	ܾ����f�k^���*��c����~ ���S3$#'i���D38����촠<�~8��M8!�K���Q��D��n~�̇4�F�[�:�)��.7ɩX$������L�O�Ufh�
�B3�]̨���=v��]W�i�ђ�]�h�7E�b�����$�.���t����P{6�8���0͓��C>3wd��M�.�jO\���x�y�Z�J�忬�`�<g��oin��J8�g�<�i��K�i�����I.�0�J����� L�Ev�*�\��U2w��u��껀�<AXہP��;�@z� ؐ��[v�����0��@ލ��\�&�/a*�u���W����#n&c ՙUE���im4�����ՠ�ꇮ���X����HB-���I��ݧ@�!f��i�@�hi�@T�D)�9H�?���	ԋ�5	I�8�S����L���u��S��k+��*�{�=�g��e>`6}thWJ�Ӻ���9��1�=��
R��P��r�L%��z��?�	�c��C}N����ؚ��WWD:꓄�-���V���>(�v���ґ������T�ʹ�_��|�@ս�����B`��~,t��������o�p�M�P!v���+�X�����{��OS�9WBL)m��B#؉9:��**�nZ�.
�����D�XjV��O9���d?��ob��m/�,�G
Nw��>�>�v�N@��%�ݟ4AQ��waL��4�u�c7�FT�ݓ@����GGǋ��a�l=���(F��� �8����)�䎟:��n���@��_TB�݃�.5Q��O�}�V%�x⏓�|�[-�ϼ��H��ŕ����i쉯��sJx�<K'����� (9Ѵ��ڻ�`C,��z���U���XZ�J�~������$�Ͳ�#�Q�2��1���[�l۵6We�R�JO�9�!�邡l��o�=?Y���Ee������#�s�B�W���8��/����V��Zh��ii���Ul���9��>G�v7ge8t;L�C�M��r�D�ޠrò{(�����G��w�������51(��!�Uv��(�g���u�ɑ�c����Fs�.A�I$�0��WH�ᆞ˥�]f��R�5a�n�;�v!��yK�1�YȓMXmE?�������G�B�@��{�"\,.����������^���_k�#��_� �Ҋq	H��!�e+5�`�*�鼤��B�4�I}��0��b�1��^(�"?�
)�����)X� 9Rw��f)�`�N/�G�خ<�Px���y�,;�����]�6H��-�pC�X�jP*���T�������/�<gDo:à�_1	k<��� h��u��b#h��#��������K�f
����
[WI�H��~$���֘5;���j��rMA����ȇ��
w�>�
iOAO�xK���Mt,	�T� <VqRm=�4Q\�Z��Ų1|��q�vW���� �&ï^���P7��]3��@\f���O��s���)� x�n�u��I�9�OX¥�zCP�; �m+'	�ʇ"K�!��=��&w����;��^�R[�^Ze��h<ӨpsE�z��H��k4_W�Y�4��������{.ݭ�����)��P����
�Eg
Y����5ū�MN�4I:��?Ʊ��H�5����� �/ٺ�>�-�@�ԫ��CY�:�8׼p��%W��p��-��5W�*u��)�/7��i��#�_���2lH�h�71�Dn�� >D�ϙF�
G+'&f�l�V��. &%y�f z���^���BeN��KW�|(��N��zΖ�#Z���X<� f0ln�)�|�S�i��I��J��{>F�I��l����$M��ȉ�f{����Z��*���990���|O)�`����KÓ��x�>_�Q}��y��s�ڒ!�[���
�~]��u���(��n.AԚ��YPX���jY��?,a� ���{��=:p�.���� 1�Y��薺tw��L.��]o������37��w�o���jS�6,(w���{2�W�;���)�Ų����9:ܙ@?Ph���?�3,e��2��>xź�J!%�~L)��#r�&����\� ��\�L�UW�V㿾���е-T͍T�Z�f:���@�V8\T�I�vx�����������,���U���~+ �K�M�x�+���T��6���}���F�γ��[��Єh�A_7Km�t�u�9JB��ߛ�3,��*�rv��39�$�����=X!��h��'S�#�>���G(����ٲ�L�- �+|ٟt#�P+?�w�h~��Q(~�76�X��h��&I!N����F(j����m�ݎШ/)F�6`v֠d�n��0���iF�A�{X���(��1}�H�����k��}�������}k
��΢f�m&���]�����|?�H��&C���L�4Ʀ-d�&ѫ�v��Ԇ��>��3�%��z-:���/m�]mM��!h9���%2)\��<8�tZg�/��V��~Ǫ���E_A"Z�/�
qДX�������]F.	uFc'�L.�b8�l;z%�?
t��q���JDjޝ���*�����/,����ԡo��� P# �%JUm]tz9">Sg����� �hO/o�t��V�'F���H�`�LW#���V�\��?�;N�� ��J'8@iF��J&��:	���H�{�֩�:�=��|�0���x����0�d5x�`�א���~�dc�Bli�ՙ�hG�x�8 �5m�v��2��QZ�Y,��,�5wF�
�2O�v؁f�l�qy�ߗ�\���%W�ً%m��h��B�p=N�o��� ��H\dj�<�
7h#��
Ow_���d�K�� 0�]�~xo0}"ّ5�:�V�;e��VF�l�.e����1������	
�B���D"���y���ߜ��d����x����Y��nT�
g/��z4-kZ��&�/�@�Y��}�6���_�x�fY���.�O��Ga���<;��2u��ˇ���"��Mdڹ'xfv4͘��,�]>Y�6�[��ZҴGj�-�c�5�V3ug�Os�	��v�Eѭ�Mũ��F�5�"JK%{��sb+Ư���{�����8�ev傍�p����0Ro~=�%a�"W�é�����J5w$�fF���H�Mx'\D�E}$ �7�����T��`���'x����~GWO*~�p0�}o��hFի�d�Grl�\8�?����v��?~��G�_�Y�#W/���n4#��3<���B��tz`�	SZ�D�`��a��`��I�|�>$*�1�C	h��m#��� Y�N����H4����9Dj�!y��_G<d�R%p2OS�w1"S�n2l�L8�<V�n,3�G1��>����/��j�/ﯞf�l�o��0Ԉ
z�bpdwP���9����	��V��P�=HB��_�<�6�'�<{�;�.)��@:��A��Xڅg+�s����&���ZEL�}k���O���\
���Q�B*Mǚ�b�F�Q�c:v}���og��_L[Y,�UFY��3њ̄p�A�;�'	��^�+���`�г�\��_m��&�bfG\�ޢR��f�+�/C��@��J戒��$)���7���G�b��Q�΍B�*���z���+���Bl2p�M�p��vsm�n��W�&~���,#ap�eo?��l��͝��@�]��x��iQ�ƻU����&�%�m<1j{Yn�'�g�����ߥ�)���.n��4@.������5"�ڍ���I1�a��cɶ�.���f�������z^�Q���9��na?j�\��jG���
1�j�����6�Q���M��-B�ig�PUv��6�I�@��J�^������3�~�,Xp��8��Pg.���k8���T��a�!U���M&`�h�����t��肟�V���4��� ��U��Op�Z�o�W��L�f���#E�n�5�߳l9խ�CF�����ݶ����R��G�}t��c�ջ"L��8��$@x�Λ2Ě"�Q�a�VK��o����J�^���R�8�	��\�:u��ǎ7�A$����ۺy�}�I�U1��rMX%٨)�W���^e���o��� l9�\��V�VQ���]E�z�@9:k^N��X%�돬�/7up,�@P0W�R���� r��H8!� %�eƖ�������9���w�}��/����B�p�����6���氩��g|M��OxPQg�iH��1Q8�|�居 ��ֿp����F�i��0�`m���H7����8Q`Gy��b7֫������13D�ъ�m�Қ�%�G?$�.C�w{K8x��?�����.�*68b�Q�[J��c�2m�b�/��^��C���D��)��2���(.��H���:���s�&��ؔ?�}R�@�?��F���V�����(�d6����3K�mν�!V�"�S�	��5An�:c��@�鉼�eg��aXH���b�`Num7D�ę��L���Z͹�l��l1L.�2I�%D"�SR�~��c[��(�+^�W"��g�WG��֪�'�W��b��w���:��E�
���ؕfQg,���oѤ;k@ �aX�\Yv��vy���d���V����M��K	��٤����J����M	�s�{�Nk-���,\\$>h��C-J��ń�O�l�n�ۡ6��2]B�)���6���U�����{�W���z�ׂ��N���6?T�IR�Lob�����-�|�Θ���L~�ͳv�3�RڕB{e�F���%�!O3��G�a(}�R�����z.�$<=����-�����R��q��NLYv㮊�J���G�hF5��<�$|��Й���E�G�4�	/�m�n�-u=�y�k�'�{D��j=����&W�0�������m"��쳆Z�o����/'�<Εo��G�G�i��-�+	|�?�'�̺��d���U�h�Qq������^���baSU��عn����y7�;�d;x{�&P��'�m�;#�d�<y<��n�
��䣹��� 粟{��h�
s�M�n�5�r����G훻����K� ��G�r뼺��u�f�e���������=�~S�����;���.U�R#�( 0u���P<���W�&2E4�<4����O%����&ؑ>��!�׻��v.7 sd���jp����U���|"5��_Q+{	/�(���F�tT��QP�[�^گ�F�.oGc�!�Gʓ0�����`�iv��M1��(XyX�����`�^n���6�"���3������ ��1�|�(.Ҍ�|�ylp�䰮>o=��ޙV7xC�N�S�o�f�\�2`l���;Q�Z�]}3O\8��6�O�H��:���
��S,���T�O�O�	ԯ��*�}�64F��w�	�k|W!`qk#0>	���Q=�0P�K��ٙ�ܪd����s�|�-if�T��Z��Xn
{�WF��$l^$X����έy�[�:��"�=�W�d�k ���E!iu���I��qKr���=S�������e%�hN�M�9�K8O�~'"\v{Y�­3)��^ܽ9/��-�������x0y�#�O<o2$?���#N�r�b1���
�+E";k�Wy�����R����O�{P���;`�3]&\*cq���,.5Xo�vVO/Fi0u��;k���&�M\����Sa@�r~�&�ƍM��2�畏_�蝋��(��l��ŧ�l[�f��i�yq� X�ed���C�6�<'čr�!�f�ͱ�h����7/&;v�SS����c�i�M ����CǸ(S_�K����L����K��Bghy"|����2�8�T�2F�a�nKkK��q��X�/���9��(bG>�Z�N��d�d�\Y���goz#���(�u9mԚ����xkfᲡ� ��������K����=�DV~������Qy%��
����X>�z���k�Cx.�Syh}Z:N�B��*�aq8P;W}���*ɫ���Q�ň�_���<��zN\jo���W�c*��:���<�I{���������weŠ���^�,f�ǹ?�	_�����#.v�L	��q �t����$U���l�F1��A����� 3�'�^ɤWvP��� jÞ���#�M���/|�W`xL��@��-��ӭ��$�5�dDd���-YU�2����O�C��j�j���b�Q^����;L���P!t���+����a>�"k\��i�Ё"�������P0�q<ݫi���[�/�ڦ��^l\CQ�OT��P�PD� |*.0s&kv5yD-��]��\�ٕ'�<�h��$U��c�8���В���A�/i�4�hs������:�I���\!�����m#������_�:b�8�-ѕ�P<�v�7�el�8[ѫ�@\��2�2j��M߿����luإ�)C�y��`���^�n���`$�a -!"&JME2;w��p�D-��H����׆g*3��z�*ن��{�@����8P�H��ЀW�c�����:�a-��n��A]8Ƒ�		i��/"�h<.�k�@���]���"�3y.�����5;��d� z,kh�4%۱/D���������U}�S���8 !2�+��&��1����yk��"2��|�������G�zL8�p=XB�;�8�X����G�X0��ōf:Lv���Gh��vھ#W�:�S�x��Z�J9j��E���5������1����;ps����m�4�CMA�}��8��B��6@�	�]���K.#���.fE%�3� ڦ�l�N,Ph�K1�A��>��(��\R��N�̐VطN"pʟ�ک����n`7���1rʌ�:y8�� ��}김=�k�L]�,<��8=��^@��j7��ć��/�˙EK<ɸǿpc��^��nqJSy��{6�=�F�����GjO�����Sz�>-��ڸo��G�����C� 	2Kw�\4�����8�!�yQ��ɵ-���"��c8�'���Lb�
�+D��Ot��H���v��[b]KP�2�!�D��!D5���	��|D�s�"):�*��9����ǆ]_�T@EK��!^J�����ߵ)9��m�q�֡��Z�g�H���.,ߏ�Ǳ�ԯ֦��:��w�<Z�i��?����E�M�l��� <Y="�hw�vd�1	�65�Ո5��Qgq�U�`�v�N��2�1��X�B��	=[6�"�Gݮ�P}
04��q�Ň'�_p<����XC�Bc�~\��o
�k���-΅�7�7Ewh[=Z���;�����h���i�ڡr>f�d���Q�^�v_n��$pxA|���J�{������g̴(�l���Dr^�pV��@�?���,Y���_rH���e�����M(ƲU�K�`;�0�ᔻ(JB�Cv-FE�����$�5z F&��k�i�ۯ�`�)�2M*�����*\�#�oo=�ė��|������JA[���%�.)���]����'%&"�#]���_�OscSl� �wc�d�:��K��~5[`�M����9�y�yV���a�3�W�B��ǥ�B��Nхp�a拿��#�<m�Ӻ�v
�0Ni/\�ěڢ��PgB��ʀ���8u���T��c���&�K���{=h��5,l/����M��m�D�^+-���!)�4��`�)0����4a���/d#��ooi�������Nno�'@���C��.�1i@�ř�M}�_�5�o$j�����U��S	6V��1}v�b�5���' ��%͒0Όn֬Y�s��Y�>�)�������j8��2 Z��KǨ��á�O�	B)�	����S�Dp ']�u��&��>i����G��-~Y�>!}�1c.>�C�:���`>�Lx�p�G	%F�;F ^�:�Ֆ�<��E��`�'�������9.Ϥ��5u�
z����I\�)�G<�6�����A@���w
���t����c�����$l�F�pW{)��l�X�6p�_�o$����K�Pq� p]+��yz1��������'O��Z��qG�It�k�,�WW�e�C���R��	2���o�%�b��M���/�����B?Q�Xg�/�j-+uU��0~:كu�?���F+�%ھ&��$� 8�̴dO�'ҿ`�!Q��#o�8��٬wNE���۲�Ne����;���Nx��4H絯v�����i|t����!Z���b���\onܨ�5��1��8+�/���ʷ�����N�y��$e���+I��{�ÿB&m��7_�i����[�V�������'[j���lʐPe�rAoi%�c2Ǖ����(��,�>�#�h�8�F�R@�n�
�:�oЭ���F1�#��^%���I/F�]�Ziv7����(|�r�/OBt?�_��e,3qL?���k��D�|�O �n�Y��a�W0���g���r�o_���0A���T'�H����Q$,ҭQ�8�����o"��n���:M�c7����`G�c��@�[�c�f���5��l����9��z�XT.�7�j�*���m�^����zX�5��$�$�������g����p[�*�%�1|�nbK) ��-��w��|k
B�x,'���O�آ-��U��K���~fiO���F��P��f4�j4�} ��G�R�����%W�T����N.�������:��{�:�g�tgf�K\�|�,C,w�Y�pK�
�q��GJ�\5�tV��0�a�H9�!ۮ%q���%	�6�8P9�5�'a`�5���s�-����`��f3Z;Rs<{�1M/��|��,W��4c]� .�M�)�`xl!9<��#(Z^�u���,�N(r
T��E��S�j3��$�+���4n�ڃ�f�S��Ǿs9�~�Wy�h�'�?�|K�a [Id�+\r��:�~��`�o�n7�®s-�5 �q �	�>������	^ܹ!�R;��������bXD�+r��|��f��G+��Ͻ׺�^� �d�*R�x�C'ra,�T�SIy���Rx�s��@�|\�R$�ՕJ�����d\�I�'��{��(1[�Z������S�JD|��ʎ��~޼64Kΐ�]Ǟ�f�-؋�
@���X��k��L+鵓�� �P4k �/�>Q��0���A��ĉ�ل�I�m_a;~�aknl.�F���e��;�k����q�R,t�,���=�V&jXyGf���M�h�2�+[�7����Ho)s�+�a�0�'MY���d��ЁBDk/Ƭ:1��!����k8�}����δ���S�=ϙY^��l�A�������!�(g�(�N�:6�vH�y�v��ٙJ��A�Ky*��,�O��^2����P��m$�=�󢕅�~�n�#�DwQ�ʷ~�C�vVo�� ��>�5Lr���^������Ah�� 2v�Tg)5�S'���`!���JKAûSj{ �`�F���|͛)L����Ề?��bf�����]�l0��� ���6��S�L�Ҥ��o���>wIRf�s��;�Vy��e�;.�G�&�7�?���vCpG؜���So��J{<�r�Rlą�Zq��7ߘ�ّ~-�jL�g�h��:e{�e�HW1VC�/�lQf1��2���`��l�v��.I�,�x$�����Э]�6�@7�>�:0΍��)�G���&���t�� ��5{�jS|S]�)f����M.��������+��ѷ��%��B~6����GiI�:S��΃�ʧ���J�g0SX?~�3�+FG����f�8?��dĮml�0�nJ>�sW[��^A�

�}�.U0O�%ea����TC�y80<��ҧ�W���(�����!6�TnT����Q֋*�A�J[�ld�J����A=�����;����m}Z�4�ͯʣ3��Z�I˃��/	Y��13V6:G$e��!3M���x��K�DX0� ����;Ɋ���y<~�{�T�85�G-�,�q���Z�oM�	x3����-Q�Y�h)�
P��§��F�kP4"�r�%��@����� �����e����`wH/��\�c�/�N����ؽ֘�A��(3��E�:1����;� ���3;7��u���j�D?�f��O2.��1{��M�2��r��;U�X�l�"^���b���0��r��+��v��f�D���(3�� �p3Q,�� �EZv4�R/yd����:$4�#�槁&��u��׾6
���EY��7�JlC9Z�+��B
�����c���W�����b��r�=�`u�򼸆�;!:�ЍuB��cB́>�F���
�
�2H8�X��L�<�%ɪ

@���}�O !���_T�T�ߊ15/B✗�I&�~�E��\�j�em���w</c<$7R	����SSX��E� ��*I�Y}#�q2G�LAG��C����d�sAz�4��֜�7�g�d(�X`
S�Y:ղ�3�f��À^�PnAE��J�N�+~�T�?�Xxw�߬�&��#���~��аC��S��y���A���N�Xߟ�l����@P����9	�ͩ�hH7�zW^�i��!��'�r#�j*G��
��8�0�� 	���L-��2֦ƺ/	2GB>��D�B5�S8�ȵ��?0VF�0�Ȁ�KQX'x-�淫m��Te���JP��t1��cU���YZ�h��cM�UI�7���)��D��╷�m�/$���T�M���4!Ygd"�FnQ�)ظa���r�ُ�ޭ7��wӎ�ËKt-���NT���;�� �4˩4�X� Z���F�i׼���Y��.�=��V�[���>HY4[�Ʋ�%	�pl�	ۄ�ͻ_~�@V�ϧ7�ƂT�Ξ��H���1b: �[5/��7��֣�m=l�G��)i�/VM���>�����Ϻ޶�2Hĭ�5���5�P� ���@�Šb�%al�[ρi��������3jڛ٣����UԪ[U�R��T�q�R���-���lLT�Qu/X�ɶ�0���k���Ҥ�,{/��I���D� ��^��I@��`�\h��w{�b	����P����Nq_���|��m�ٛxg������[6O�H:B+y����i$�G���dA.K1h���3�k6��%�謲�Y2-�]��������HlM�QQ���$��,`m�7���,�	ò^Uy���`&`\%����k��Nf]퉧��u'��.��[fgE?�%6[O�+'�_�dU	�@S���Z�;
��z҉�E;A@��&@(*^� ����4�1��?n$��_W�<��=��)�M���9hƝ��z��^���_�E2���V{����rS1)����D@����p��hᶡ�. =tٰ��j�lG�ď�S;Ņ�V�J��bH��t��A��e�q��⸩�Y�z����Ł�騯t���Ef%ɉo�@d��談[~M6��k������e�'�F�5'��ݯr������V��TMg�L�ܵ�(���͙�_��~�h�F�`�%��pN�!]	�E3P��0�8���Q!	�hA����bab�[�i�����9k�Y�}���� N���Tn�l��?v�V𜦦F�s��=���&ع�E�������ok���eO����2�sĸ�$Y����(�������|����<z��P��Ŝ�����`/�u�8��5�k�ŷbI�"��	��-�O��&������I÷|�!p�=�=_�e+����+���~�]CF���S������^�Pf��������?*5B~8v��)E��\���*
,eu���y��/�L�S��z�^����'�R1e�B�~z���WS�m1.�
ˏ���P�!��;���o��vT���۬m�J�3��~�{�
���d���N�'�s �)ނN����	r�����:�#��n=��ΓkӡAqk�z�L���`8��4U@N��[�k�rW �se �X-�3(A����DG}��{�?X0F#4��#u����\iH0��\ s|��+A���_��I�2��ߔiW��1�V>�3v��!0 �р:��RY�N�u���|A*�Z�l�Qr��E���{R2e�������Y[$_��7��ba�3uƹ�Q{I�>�cda^<��!xd��_���� )S����PlB&V�읖<�]�\H�����,9u�� ��T��L!�2�ϭV-`���
s��y�sR���)i,|-+]��F}GLg�@��r��d���\��SM�[3�<�8�/�s�=@r�A�ݖ�MQ���.}�"��\���X���)&�4_�ۥ#K�`�ys>���n���w;�����+��c ���#c\qG>�x=X�٫j�{�"���ǒT�� E��~4��TH�f��|��ȅ���O�չm*�o歿`c��d}��t��#0�9eۍ�ϻaM����g��O=����t�n��P����,�]�	0��@�u���|��e�(0�w�֫���Ċ�2��c�-�N8���n�R�gè��fM���:����G�..-�oJ��}Ϲ��)�`���U�����r��������`"w�mr�B��咘T�uZ^�=�z�Z�F'No��.�kۨh|�۩׍6	�ӟ}:{nRۿa��+���)yV|�[�y����Z!.��H����cm)�_�oS<jc�r���f�f��^V"<�؁[�\�L��?�S��a��h7ZeVk���'r�u�b'<�P���)�ҺD,8�^`��,ʁ�V��EfLp|��&��[g��~�8DD��v��|�n��#7�Yx؉��9��q����Fk�֊ͽ<�H;	`JP7�`�]�������4㔬Yʧ�������a]�K;-u�2��*̞�#�2c	�B�]�D	7[ǔ���Ƈ�$h��}=�q�H��dw�#�K}y*�Y$��1?�?ED�c���*��`�}	�F�	pOD� ���b�Z5�l0UR��H5���� ��Զ{U�g"������)wY�~����W�+����B*'�/�?m��O�n��,�z%�Ȭ��]�w�݀_�\�Ts��  ��V��U��e)���/C�w�anاj=�sJ9"4�t��L�T�<��I�e�*�}��pCh���Q>4 i�):����TY���օ.�|#ZԈf�]�ڏT�?^��R��PD�Gpn���نlݝW@��'\�rx(m�E?����OJ6H�}��vq����?�O�0'�Y8�r�ҏ2�j�k��^���W�� �mO��@�8��%3pؿd`�8}b�b�R�R*�s�@�Dmh(�%�37nI��B����zg�\k�3T���aUPj(6~�M�Pg�?U	�����r����O��/�gI��:��do}�퟽����(s���ц�y��m�I�&�K�쨌�z����"5�y]�_��pP��H��7�w|�R����#w.f����zW�%❼�~w�<B�'��.���B�I�9��gˎz�l��N�K�yĽG	�"�-�PN��8 �\���AP��J_���Y��Ϯ]�W��"H���!s��;��;^��UqD���v�=?鑼Di�O����2��p�p�i�>qEw*(|�\wRy-U�B��r1a�����x;A��j^y�Ċ�^�v*�����O[�DD�L��_�@���G2�e���ۦ3�Z��nk_gJ����!�t%� ���)�d�6ړe0�$zj���D�'Te�9E�fH���T�0�R�m�n�.s�>ȯS����ΑNM�5F����Ӑ��5�qk���ĵܬ�W4�Mx-��>u~����P��T�j��j��f���5
�Mw��~{<�"V�1�M�<��)h���+h-�����f��Ib��6�D7=Đ]��� ���>H˕_�lp�l ���h��5X��!�z]�\Z� ��`�,�6��G�4�?x[�t��,Gv?��2P����x�6k/���Vg�,o�4�]�fǒ�):��7���0$(Jx2x����P�[QB[R ]�����5��$Y֙� ���U��%x���?@L��k�t��!S5��	˟��z�353*ݽ�hN�yc�J�@��s@2������5�#��vQ���śz��}�C�����h�ǁ�Țڊ�m���5˟�x3�4��v��K�t�-��|�����]UvboS}ڶY�}��R�"T�����e��ʺ��(�����g0%4�����0��
�߷<+�Ճ$;�T>��#L��#�y{h8_��w.�,�&�٢���9�N���Y�Dig�e�h�uF���;�8|3DA;�a�s��!/V��C�XТgd,\F���G�m�{�/�o�:�7�3:��q!�Nբ� "�t�2�CQ�v���{!�l�E-�}gȇ);��=F|�E�������b�0�L��L��T�����_�=����O��!M�|�]�k�T��;UC�̲*���,�����	�)�?)��܀$�ky��@>v��Ĥ:_��Nh\�q�1�Nб	ik4�T�!&AW��z�3Ιj�vj����C��tw�4�>봡����Ku�y���cƴ���x�Kb���ul̂J�Q-�k���5�QD����;�ٮ������Lv+0#o|U�ko�,?m:MC���F7�eF��b7^*��)����$�z&g{\c�uF�ũKʧj]��{�^��+C'��!G�!��ٛdM_n[U�8\v�m����nQt9@��.`Gą�d�-�;6�׈hg�M8|$/Ks��:W�iVc���zZ3P�A��z��F�/����a�[���<�e
ۅa����.������:M
c��}�B�ښL��U�|��v`�H��sWU�]̦=�gT�:�m{8!��\��oBO�H1�+�[콥�Bf�P�4N{��l�����j�B.��yF�~��p�Q��`P2�K�����ӵ��E�4T��p|��U�K��7�� ����$�F�(ܞS
ZayXD��j?�WT��S�b[�Ytep�D���	�|�����F�*Y��51*�'��� �ض�.�F]����[����G�Ր�����[��JV��Pme�)$�/�QW�A�t��/��hpY,z������u������9o�?G�OS�1�C"�ehEѦ	�����L�F�{��U�㱲���HzGd)4��-�n�c>U���3�k��zI��Je��O����לf�Q墌7�� �,�����@���zg0�~��Ŷ��2�0��-ߒ�}8�	�ō�8]�ΝL���%ѼE�-Un۲�K��]�fLZ���)B}C��h0Ȱ]w�q�۴+�p���� 4ox�&��Ե��+%�o�]�sF�/�o��S�{ط�Fbm]t��k��t/Ub)��Tli�Қ���&��^Q�z>��K/Gι)d��9Z��q�����
[�a����;��k�D2Z1P�xEKȐe7��|��̋P�n��}>!�0�@�F1G{P��/�^�Ѧq�Z��q��2߸�$W� ��sa��ԷC
�D��[���`	���s��z*�(�$NW[�d���&�*�90���{�ь����|���)`ȭ�����2���
|�۹"M�]B�#x_fu��s|گC�ؠHcg�;Ujz�D.ċX��}�d��/1��B�i�fO��>=-։�Kˊ��Rޯ������l�6��?���Cm����ޫ�ǯa��U!��܇qK���.��GNM�[�b��>�	B���3\2˃
=r��G���4�sN{I+��п:0���O���u�+�&,�|C�*�s#r��F0wcnf�N�@�]��$5�gnV�
��#p$[��vq=Y��Z��94_��+k ?_��f�p��-s�j$v�e�yHq@���t�c>=��K5at\�'� 8�\�i�G'�/�.�֍�,��0KM��B�㘇��c�!�2,0��sMU!�T0� ��.=��c���m���cy�]h��B�h2$r�=d�,%ҵ���"�{-:^��7�<.!tY��tS/;㌱��OE).������c�8�PY�a`�$ZX�!�Dk�'�Za����E�����	��Q�1�7�;jV��+G[��-�e��ћ.���>�4%7O�o�"&�/�hJ�vC���p/�9	H��!�={�~�DI�����'��;��aÁQ���x�v��鯂XIp��lYf��d��fA�w_�%�(Rf�%�?��p_7 �FҮ��v�,���i��R�����H����È��id|X�)��^j8!��A��:t7�>&��U� C��^R�dXÌ�/�^���r3�Ņ%ǌ���W� �S�+���x��������z��²�������p�E5��>"�0;og�Ue֛U��9���\Д����Hfg���S��i��8��+z��DY�GgV�z�ef���� ,4�s<I '���j��O���/(�1�� ԩ��� h�.���:��?����7�䏅�����`�9�vqO4��i�����X�F��� ׏'s~Dif#��ԱC ��'_����.�s�����s7V�Bf�1�"����l���B"�^�u�)������!��Ȱ!��g�)����$y���P�����7o�!�(��3��f]��^��fƸ������̨o��dn�ZA2�_}(��.�!��8f��&��VۇU�f��1���0<D�Z!��b�t"iх �� �-�h�\�[C�I�t:��N�qZ��B�p�\�N���&�Z���>"���6��м)D��	=l5�E6��$1x��̇�(;c����� Q	TB�IP%�Tm@��AAMx�� ByRn�������&_��n�hJ
�-A�J-����6��ݪpf���!����d�Q��wU����蕽pb_]줍���ZCB6}[���uK�F|��u��.!��0��@�/-V��ޥQ���4����=s��O5�DV9��^��!1��+�E���Y�i�ت�0�;��)�6���3���Mp���^E��N\�
�_�@��a�����`����j(3�;�4w%��P%gC�<]#�$=7gy�o�B�cuY���55'��>;����P����ƃD�Q������0���!�%Ͳ�|b���*�,,���j���l���	'�f�ψw;"�����P�g��y��N.����v-9B��YE�
���)��)|IܾU�dİr/���w�s]���-/�<�D4s��+�v��h�g䅏`�>о��9�N=06�@��?p�I�<�BTr���yX"�?u@(��b��Ut�A!6&����i�B�jH$[�d��U2b�A���o�;���X�[�m�&X�tzt���}�T4�)a/��gu%��G>�5Isw�ЋE��=j�֢�}��؁?�M�ůp�<&z@~aL)�O�#��ה@q�*ߟ�R��S5�-���K)��C"x���|س
�)���l�W��m�)1t�i˄P��:�,^C�;��9>
�i�-��F<�q���3�_Zgc�lD7B(W [��9\W��Ff�m�O��7ّDQ�%�yTK�y��.�pq��D���ٴ^>����>4S�w��T�Be���$�,�TEW�T�nk3S��B�}�\�%b]"�d��A'Ah�M�2jA��}�^�P(�C��n=���;/T�8&��,�Tla�?	��W�����[�m��b�ZȰZg �O�ԛ�r�cKv�^2��:���jI�{�k�dF��Ǯ1"���L�]��\�dT㭏�|vF��_�}_�mfM�qܧ%Ē \�?Cq�J��Q�P�D���
.hC�mr홦F�u���v��w��/�Ԧ:,���rՃ	+o{6' �^`��S��~��<��`�c� Dj�7�ul0���#���XĒ?Ƨ���������O��瞹�����Z��6�v:�k�<�_�A��z��T��u �f}��B���ҿ�ϖ���$|4���Y(Z��[�'4���T!ݳ��Cū�q �>�iy,O2�X?*T��$)��ĭ��)��0;�r&wiy֕��A��
����z���#ʀ�=�#�����	����,���G�鉽כ�´���Z���K�)�/�����{k�ꥀ��á|��S޶ƿ�H���Jߵ��7�
̥5�}w kg��Ǚ�"�E�̔neڵ�F�,���r�v����xԋ]��.X���a�Ƥ�E�� d�@R{+&+wƉkސ�@�p��PO�iۥ7R�q���{kF	
��Ynĸ*�࠸�|���_���t����У�rK�@��CJ��2�y�I��b�$�x�$N6D��-��G��
��-��s��gP���
f�!���� I���ػI�񀔌u������ys��I�Ox��AԀ�+�b���t�u�ɬl�%j̰q�-)���؜�7�0��b�-�|j�-F�Qxl�5Ŭ�0��Bp��{\w�S��}�Br\�61�q�7��հ!�ؗ2��=Q=���m�aP�$E_��tU�68��XS�}6z���.L@�u���/?�xD���-~M�xĶ�[z�����4��D��GOzQ�6�D��]�OgF���$~	߆u.�PQ>�THS�Q���t���A�����l�/�s�7�s��cdE�v{����_4|�1�Qy����)�7�f��8kh?�פx]�l��X���w4�#�eA�7Pg�J�������v,P�0:�Ǩ f�d��-$��sI�2n)2J�˟ύ��:Q�nx�P){H�B؍�'���нɻڳkv�� �]�&���|�I��YB�i�����S�\��N`n8�mg�������9=`��;�S��a;f��64}�����U��~׭��N��g6"��i�0#Q�E��(1�?wӓ�+elc�c�k�3�W��Ai�)���4?� eSP�ò˝s��V��!��ZKt/��U�S�����R�+�#������o� �i�ӹ���əBUς<�X�T������R�y�0/8G�5��Zc�s�X�>��N%����b�[��Y�!.�&m�������	;� s3�bWY�=t��%ަ�ȏ�X�j!z2��yJ�SM�PY�y�I��J�k�w�"��܊����Ө*V�}���9�]Ҷk_�ߓ��E�E�-U�P?��Sm�5�RhHߢ��|�����,�e�tR�
�m�����+S�*cb,� 6|�X4[��U:`�a�c�.�>mC{��{E����:d�֝a9�0>%��V�H��h9C$��[�+9mb�6`a��ʟ�l&��h�D�~�D���+Ɗ�Jp0q,�ߚF�E�tZz��Tv5�8�y�]f��w���]߰����Z$h�z�D�h"�^혘V�`]�)⮶�26���xoۍ>
 �xH������x 
uY`�2 9@fh����#LeK�Y����3:.ּC�Sn�.؊�n)��y� m��N�>����uvW?��{{(�ګ�W���4_���~�� ekE���{H[{��L�1��b�/)��/N�E���)���i׾�U�?	a�H��i�'�lϦݿK�v{w�m��P�It���z��8d?�QS/�,����r(����s6ʀ��i'#P�HFޟ����:)�ބC��QX���.faY�0����L�F�><��>���|qH1��r�����=Y��s4�*��/՘��(�xʘ�4!M�z�C��׿�^'S�V�Hޓر�8� �0�"gNy��_Tµ!̚�0�*8�flf:v��T��R�|��̓�B�����؋�M@�3���Q��.K\@	i5������a�!�4��w�r�C�m���v���?IzZ��0[���5�X|����R" *Ҹہ�g/E7c����AE�1I�yZ�W�6ݺN�A=6�r�\y=�1�s��<X�{k���jWxt�b���gQ���c�08N� ���C�e�Jb�#Y��������T1	W��
7��{w���v ����e�0EK��O�ӕ-pp��. N�3FIJ2���b�W����]7�O�kV� �?�/���R8U:҆�~p���/�Q���&�䓽�y[���}�A�#�(3����N��C���<�������@���7^���?şؽ�`����QW��֨�i��y��g�%��ٛ�lT�DC��}U�=g��0ٓ��:6q^�`�w?���L�E��?�Av����&���b^����l)X�6��c͍�VDUd���6ش�����1!9 �������B���#m!�O�����݆�ks�o3v0��fz�d!i�P��ߔ�>MKof�(	�.).�3�1C�:�i��� �m��I`4�J4E��|=1�r�8�[�`��w�� �k�λX��Ơ�_�П������-K�!��Q��}��t����l�u)u�݄X�����jS|�c���3�dv%uq��O�g�5��aF���h�5(��[QP��Ic,��&�����P��E]�������(,8'�Od@������l<lrM��A�i��\����C4�?JO�%5;O� ./��X.��C�@���1z�p���mk>(��h`����2�6���^�	�GG�\=]i9�� ���ߤ����dF"d'3�8�+8`Us!�������R�����ֽ̝����J��sjD�/��G��{A��(L��n�t��MH���\����!(��c��¶t���ѳ���w���2����-�됇�nĒ ��b�ϗhS� ��|l����S�!��3B����#��OS�D,�I>q�h��T慻|8�7@̠ٙQc���@�+�r�!���&��q�Mm���P/�P9z\bK�j�F� �՟r�\�!����V�P�סguZ�4a"?�4p�oT�r'�D��c3��ז��aa��p�#���п	&O�����	���ZXa�Pn=^�@������� �1\�1B�Ѽ9����� �p��B�G��7GJi�Ғ?�<�y�~ӆV7"� p/��O�
�z�%��lV'%����M���b�AE��q�@V`��Uo0ҬJl濍���/�>��@^ag�`��h�!��#��n���E*)����\M5�yM����cEL����Vݿ��)�UjÞ,�
�(�.	���W�`b���[�o��b#���ab�	[�x7��k308�k͛�}�X��B�o�L�].��X�e���y��6�����Ά3��3ˆ�g�=<')��K�(���W?��w��jD݃�Ϭ�\��u��W�Y�q"D����0b����b!����q	�����*�� A�4U�u5�BS���W�~��b'%K���H�`��F�Ⱋ|��Fd�fuq��B+Ebau���Yy`�-��
�=��'��E�ZP�
D +w~�D��&����4��+%�W�ar��B�[g����]�i��l]px��*��ʫ-�&T,�����Xp>�1'�j���ji��֝:�����)����t��M}زk]d��Z�>T2����������l�I2$�iFb,���'ol4���1�����	at�x�;
Ҵ��O�+g�v���������V2F�}�b*$9(4�h�~Qќ�^_8�P U��^$�����^������j�>�]��6*�0Yך	��_&꫽�U�<���-��S)�D�w6TfR����z�Z9R���� ��fs@��gp>N��ֶv�I-�l�z�@Rp�����+�n�ӳ�Uh�g�FwZQ:��߀p~�>*�̨�ʆ���xQW_�,��HI��������A ���h�$g]�m�M�l-WyS�ZZ�.���G���s�3�7_��BY���9H� �R��ܾ�} \�8���R�
��ܒ����� [U� �����C�i�!��;G}�u?xv��T�Q^V%�B�Z�X�SB5fU�4�յA�#�9��3�W�]r��}�<4�{/��oɂ�`�ن\��94���W��W(�����Fϻ�4�.ך&'f�U2�󛪜�^/��$����<SK�
:MI��i�h^�ܽ�B�1�z��cH���c���s����z��.��>�ڭ�
�Z
�0o/e�� 9�y���t��?�8ͺ�S�\a��ǯ퉿j�U�2E��;��o����b~"8T+fN(�=�@\_!X�D������ʋ�	����_��Q��
�>�uK�/L��-7sᚻγ�cs!���lTeOR燰�ŋ��%s�łٓ2�4�}����
�_�ȅ���Ǵ��81%�e7�c 7���[��X������Fu1t������&`�J��$I��+h"A�|I��|�jaD�?�O�+ⷔ�I���p���7{�~�Q�1�*�w%�?��i87�O�h��d'�>sx���G=�ʞ /M;ai��y�X�o���@ٲ��@eU��{�(;�]8$0(��Z47�P�pd�A��Ե�L�K�	�Pڵ���b�[C�����lnr�ǻ��}h����a��=A�f�6���RA^"h���F�����~�2[��b�3�~�vz\J�ow�l��(�KHL]D �����A����>���M>��>���@��JAnG�#Ej�^Br�,�j^=�)��љ�l?6�z�����(�V��_M�6Q����҃�W�����	�E�~u�������Y��oe
lV�l�&M��&wq��l�N� �9����Ӫ�Ƀhx��F+Q�AT` �&���;:]Q~V�o(`bj������S���#u�[� ��U^�ٵX"6�}��1����g/��
�ڴ\�	��s@*֞Fbc��S!�4�P�̷�o�x(׋2a�����8�){� �&׵di�G���A�rn<F6�R�d�!5�.1$�a�+υ�9��xp|g����\�\%��#�"�s0� ���:L�],:��;�Vi#$�
���ʱx��Òo� jΊn������<�t�>J3�ɮ�(F�v!g}�6��l(Y�:�����P����՗�����j�>�W:���-���gT�����;}�Ŗ�S���D�01�MF�9�ت�@��xW2�8�U�wb�`v�rK��UL{��yٽ��+����H�q�rgz���f8=�¸���E>3%�p�5=G�j9Oʷ�%K��:KN��g��7"Hxd{?�FRx�h9��ۂ�V����m��C:)�L��-�Z�h����>$�����DWm�23(�k�	@�bw�����J�ڰ�B3Z�M5z5��v6z8l�\ɧ%V�_sf���|?W�o���	�pB�_�ܞ��;F����&}>R���#/s��ӂN��P`N�ɂ`��Y��st�*�1�b��g����[B���5N���FMX}�gƬ����W���CZU#�f�v��6n��W��\�ba��L��.�_��_�����~�|�� �jcj��O���{`!�,i�?}����˵n��q���ߔyWF&�(������B��D���Cс'�[`x�u�#��2��̥�2ʲ�O��#���"h�����ײ�����zZ��_V1?�Ф�d-)3��>���ÇP�l�3���A�!��tE��	6�$6��c�	�^:���ye�%�>��J'N�Nq��>Es&����~ݥ��B�<l�Td|��G% ~�w�-��2��	P,���\��OxJ8U[�.��D���ʼID8�T*о�iEsjp-i?�ƥ�O����c�8���
�^�T��I�2��x+u���; �[�s���+3���b��P%��5R��}�:�&m��!h2�#�z��ҳ��g�Z���l�5�\�#,�����Ȓf�c��X�xw��)�`�At[���Sa�[��ų�u�D��)a�c�u�1��$����&"�ʂt��!�)�X��{����TA_���ŗ��2G?U�U�4������U76���l��nA�ޅ�p��D��Q�g}�,]���67%�����7�>e��b��c�寘E_�r��T_�mHҳ��j�,�oή�kQ����*N������y��5���Ҏ��u������ 5u TS
�)N$��&��(� ��:�:�g�]@��dj�9�iӗ��465=���0Y�6]�6j'�o^#6��nE���=_������ �#�sܧΠ�mt2�k5�,MD2�7n$�Y����AG7�:Ӷ_��-V�5B9[�����S�+�`>z]~�ɪ#Uփ�Nbo@Gw/S��1��~��������Fً��e*a�ӳ'V�����>�vL��cU�> E���Q�1��^�eӦ�Z�Y�q;б�I#�٩a�V/J��{9o��zٴU�y�����-��O d?(c�m����Gmt�������H�Uam�LH��=sA�
U ����Z��W��Ϲ�.��$N�Z|ө��aw,f����o�|��_�vv��C�	e�o8���ǣAߏ)J���&M�DmbB��Y�-�tîg��ɕ �Ȳ^�%�q��5)��Џ���
Kࣦ��)�ie�>�Z�ڔ�Tg/+k�D-�"bs:Mgx�)��>����o�4��a�U4tR/�!<H$�`� Zw(2���O�	������M�n�Nd��N�J:���o��t�K�g�C����#�x�@�b��!�𹃖p�]��Ņ\��I�ѽ(�!�S�^N{h�܃%�c5��MJ�m1����[�bAr�thU�V�zi��Hh��d��?<�;r�Y�÷��*�Q�/����~�ܘ�-|sW��-��.}�̴��)�.���a�@\��_Ү`6�KU$�*��$���Aŏu �:l�O��xcك>h/������o�⬿�H"gp�W����(PIa�XSg��K�>``}�WO�HHRw���z�2��)���|	��2\��	�W����g�RI�n=�~�ۚ�΀�4*��h��,U��ݸf1y$Z��q�,���lh�7G3Q�}p�Ŭ���έMT���Y��F�07VI�
i���t��w *�u��E50��l�~��YIy�U���rk��+������>�A���i;�>�T�H�+꿞��"�Ù��E�}*��;�K���o&���x�
n*���N�)@�	��2Lv����A�ͦ���7�
�n-Ӧ��'!/�pQ��p٣)q
�fT�w�W�p���B�E�k�#^Bn�RV��a���"2V�}?ҎƹgV�|�(���OY�Ǹztb6ü��xH+�9;�W���P=��!�OG�٩�G�s��L�*i�kO(z4�W�g�U
�z�p��C��o�w"/��6C]�"ٺ�'(���S��d�!���P�X�otk�� *蜎�?���$i�!��G���������׉֓�"���'�f������h%�ݧE�����O�*�d���g���C�E���şy5H1��R�?�A��83�@+�o��V7����fߒ��h���!C[%���W5f��֚��fE�z8J���{�E�n�n�f�Z�k��9�S���Ӝ�Sz�y\�D�	����6��j�r�һg�A�k�(c��"SN̘f��*r{g0���z w��ٝ!�Tۅ(�19᜙�8_e|�C~���>�����Ҿd��wj����z��?㼻���y���^�K�Y�%��������t���L��\����Σ�'S1S� 1(p���N#��C��Ĝ���5��ف+g����k�<�["F�ߜ�|O��<�����z�S;����E����N^�37�Q���	�̫'6�;SN�*
!�vQ�0*L����x�JrjO�^Ҙ/ˑ���������(��T-5����\�����qCD�?d�H�E�t^՗%��'��[�p�I�sS�)�4���\v��N���D)�?�𙞺�����K+
��</����S�\g/,����(�/�=8�b|{\Û����j����I��ǌ��U�z���ԁC�G�31f�Iy�?�	$��S��!�����Z�z�mE/��,�f�������^Q"�fa	W��K�*�[�^��Gy�b<���v��W�:o
i�זH/����F�kh�YY�&�q��pV���0�:�����r�v����N�Ew�e�I�>-/W�.8;�M\� �?n������xI��k�(��j���ہH��D�/=��5�T�?���V)��rKeݳ����W��E���˃/�W�k�{���0�u�G��%$���Z�0�%�i=i�Z�~�G�5 ��4o�.���NU��"�~�H��鿫ŧWKքpHC�{�^H6Q�Ko�
�vy�0A��۶��	�ci�K�,��͓ţ7U��m>����*�(�~��*���ig�1��y��{��RǼ�pBA;��+I��e���R6��0K���Ifz�8CD��F�%@&��w��\����5H�M��
hьB����Tr�X������1�vTCH�r1 �.I���j��
wph8����t�is]&]�Ė�ޫ�=�n�臨>�O����K�_��Fp�Vch\}�6V�Δ���0;lm9���/HVB?IW��U�7���~��]���֝��W��[1�to\I`��9V��t.m֛�-jD~����:)${�1Cm�x����R ���58���g����,�l��QhK
?Ŏ6Z��Z���Ezv����@/�V`�i����[s���ܠ]w/5%��T �!BP�_���ﺂ|<��?atܜV�ȿ����@omH�@�[k��g�o����*o^�W� �UD�k(!���Ydh��w�A���)���E�MSܽ]$kuOP6p{Ÿ��O��]�aI�;\��Z����x��˄!��g�[���~�5I���`hn�a�vێ�G=�Q�'����~&��*�b��Y��$c��]� :7�´=d���U�m)��������,�1H��*��?��)��ͷ��hH�.ŶD�4tL�@��r�g��7�3�q���J��_�+�Ȍ�:��m|�>���k6��)��Q['BCNH�3�?�p�	B�1��rӠ��ϩ�v}Z���:��D6}\�����G��*ڌg�j���r䩜������Y��nJZ��c��.}���WQ�kCHg3R��BzZ[=���l�m���(�������슐��4p��L)W�'�@a�%B��}�i+~Y�R���h��+t��� F?�{�4�'b<�)B0�V���c��&���@�%R�1��IcDMlO~t���,.Z����$��E�π��->�@��႙�yظjpdF�6���#���6̩�N��+����ؽ��N+����X�C�z !Fw�� g�栜Q̅��յ'�k'���ں�&�'�4�#����R��<5�l��w9�@�\?��O��/�`��u�9sy����=�Qk�t7*�-_ݓ2�r\�v3%��̵Z㔶7uH�M�SqOy��ۣ��L�lL�V74�޶�Q5<�o�\J7ݏŘ���� �ǽ�t�}"�Y�i�͔"��y�"m�m1���M�x����j"F�Sؚ�t��Ayo8�F(�t)ޗ��	�F���xG���]�n���u�9��AV���
������` Z���L`���P�E'F�����c�v�y����̥��3���.�H,�_MHC����o��;q�[����Ka /�
x���I�Y;��Ek>G���� k��P�!t,�t�P�^����H �JL����s'�>�bd���w'䟵F�5�5��^�m� �a��_�CY�t��;髨A�F���r}!cf���v��Z���4��?'u�Ԏ����b�uJ!:����c6VN�`.��Vp��z���0��u�02�
�_;X1O�W}L��_/F���p<�A�R�#��C�-)1+e��3k�?�D=�O��}�m��QSz�C½�$�GM O0�0� ���Uh�ƕ:Sg�vhr
њ�_�	�Ghyвx�B8��}��fJU��clm��ݗ.�U��7�J�AR�(��H�潸k%?n2ఐ9ږ!�C��8��m�*�o�,&��u�Y^�S�? �;/�WR�p}��p��P`�
�~�E������	d�������%a�T�H�$�U��]�g/:�|�GHC���\�/�L�����*#'y,@(I����/�	t
�pȼt���ޤ��/�c�b��m�ٮ��xkCy������]⇷�)S(�6��&Q�\ہ!t���bp�T��rh#a��k��&gE��4��\p�{	�$זСx��JZ)�)8�:�|��}O�֜��uHqTX.Ă��Y<��e�UZE����_��m�Ci��mY�F��e�۞勞�{UV�m��Ν!���Ow��C�r��x�EPз��Pi��FrYM��$D7Q��8L��)��:*��f�� 
uJ��*|ˢ�$��*G��G��.����6�'�o�G�LV�5K����i��}Ǒ�c�9��Q`A�OJ�{����Biţ�	hK� mQ��)Wu�`�Wv s�)dyEcm(W���p�~��˧����$:un�������^>��V	���O@I�q���vT��27�ͬP�.P�t��#�G�����j;��y��fn� G*��u�7�������/�u�T��;xm{hx���E�u4-��Y�a��TU�Si���H��jF���K�1�e%�
�)1Pj���b����B`���
�9U����B�Ƒ�noǋDu���P��Zg��Zɶ}�&0��	+��aVM�=�#2�[�#u�q14��v~�����DiP#m?�����}�S;cn�j�����9)�zQ��c�X:�ƚ�<� qr%�a��2,�kS�

����M���zH�ѯ&���w���ބc�O����^4ɹ(~�L�^�k������q9�N��Zę�Ԛ��LB�ǁ�_%d��Q�����UӒ�+����i��:�z��'����~l���:���0a7<3��ꁖ�����HZhIgKm@�O���~B��������(-|�pD����M��(���<Iƥ6�4�Kf��V�9��K��e�D��+���9WӮ(���͂-�Ј��ӽ�e��t��Xt<��S�LD%D���V��s��g)��bߘ�pE��	���x�(SV��g��e%��Q|=��?��e�=�<�v��97�l��[���E:��NC��D.d@���ծ3b��s�l��^�3g�\f"��Oƈ��s1`#����xf���%�>܍e�Q�y�7��8�t�'Ҫ��U��Ǣ�ᭀ��7�˿.�5�����~_u�p�Ҍt��h��`�{b�Id��������\s���Ǌ��=4-����ց�bB�jI*"�������h�a���,/r�/�^�gD��K,�v|�Pk����f��1Q�������$�8����,�����	���쎿�w�A����ܨz�e�k�V�;Umn�
��ō�q�%h�t��Թ:i��)>�u��R�y]p�u+1?�[ٗ�ۏ\n�~�dI�hD�P���/>�e~B��~Ȉf�,�Q�eǴQ�k)���%s�S-C�8�4��7�鯱��Ag�T��,��ڕ�FU�w��� �V�$q��r��XS�5��c7��]�E�����X��t����`�f��X���b/]PF�y�5��]o}1�h�v.��p(�(�X�gG���8�Z�{�Զ|�)�UA��)�h��;6Ƽ��B��FQ'Gh�;��Q���jq.h�YjK��%�#AF�w�k�����W EQP�x�HFE��З����|������xB����λ�#[A@��Ӧ~)�L��b�s2�{�׏�=�+@����y戨Gm�՘�Wt��v��*7�T���j�m�Z�1�?�1����%�kz��_��;F�HE%��A��x@����QL�����_0"ؒ���K�߈�\H�C�Zd0��J�]�����F%��d`�N��� lp�Ec��H�o���ؘ�Ƀ����;Y��{��1&�;鳪����.LN�@�A19�l;�3q��������;-,�=,Ȓe��Yh���v��p4Yvɓ��ʚ� z�,��(4 	9<jy^hM__6o��W�
Zo�H��&�`�iZ�4�ш�lv��kl)sk�[=�u��9�I��_�O�N�>��D����:27�������t�5�N$���а�-.����ئ��
��C��Ӯح�G�XP:䵶M�=M[��kqo�s1�M�y�ǄB�GD�FGc�/�	I���܏C�W�K%�-��g���}��~��K�����b�Њ�U���֕��S�����v�S��|<�Y���SIz�� l/����%��'��PT!��_��xӗ��L����P1��EYx/�<�_���S�1����t�
֖N����]���+�q�#}
���L� ��� ��*0o�j8���6x��?��m�^�>��u���!�̙��♖il��IXb��9J�:��$֕��W�,Q��b�Z���՟�R�0�v9o�6�)<���e����0H�j} 햃�����y��j}�k�9��{�g����9^�/�|	�'�E��T���Kd�	i��w����x	RU��&���S���l{�\
�ho]}��c�����,�c�*��Ο�C�v2爁<4'�	c���oM�+�8Z���ڙ�Ojʊ���w׉j�ؚ�Њ�`�&�Ee�W��?׊EJ�-b>[������x�����M��Zd����ֻ,uNQ�hO�Q���_����⣲�0�����?1�[A���ĉ߉�%�xJ���T�7;�#���h�=`^���%'aO8;�8�1o?��aVE�#� �KN_^�L���Ix����6���~_�/3[Eq]Gpz����Mߐ��ުMe2c�j���>��w��ϻ�L�E[�H!���1N�����M�~w_MS��(���ePJB�,e>��5��Q�����4����*
E��?��'M�f��W(��۾»�[6����H%E�eܙ��W�K��^���h�t1#�$�ܖ���)v�[@)��gn|l�����T#??8?n�Qa�qZ�TJًF�O�؋���5	��]Er3�2!	�e'�+9YU��e7�F�����QF	A���)�&qA��~��(��U��Ӟv`c��$	H�cz�ޙƝ�-(�x�6	ⳡec��-���k*NEш�4�N-x�~�[�1��f�";4���E;�iD��� n���Wt�uay����Y����M��#P\�1��J�X����Ӥ"�?���-��O{3ya#��\L���<E(�s�H����a��s�?��[�=�{�9vr($�@X��F�~4>l �I�f�s��ܟ��6�|zjn侃U��7�I�E����Ź�"=֙����!|�V,}� �z���M��7�Ǌ�����s|#%Q� 4ȼڧ��A7�� �V���'�$�-G4��#���1��n߅w[�s���,Y��b#��{-�W"p��-��$�mk�P�$�F%Ԓ��:_ j_�|!���Af+��|]a�6%��$)�l��]��%���aRx�c��lPTX10�\�e����?JH�.���|�F!��+g~�vЕ�uA����Y�*�X�Fs�4�,$dޖp5֜4��Z�5����TD�jD^e*�hx������@;��_ԟ36����Y�w,�H��$�L��L�͚:��߮^�7�"�!��Y��<�t2���N,-ba��RAV������BŦ�x��=X��2����Ug�������j'��«6lm;�&�����9.���W��v�1�o���F�&.���!�l��8E��V%MA�hO�<E{��z+=و�9����+$��KG�l�7k�sܖ[�u����Q���=�y?-yA�Q:�h� �q[85{�e6��P����N�D�d٤[E�/e�����Vq B_�[�T�2���m���H���N�Z�@�jS7U�3�� ����!	���-�a}%u�!� X4�h�G��`)�9�k��+�V��+4����|�O��.u��9<ͅ��	�c�)�P��
��ݜa��2幚�A<e����-���y�l��z#�[QyOw��L��x��~�#��`y`:H��I���kX�n;���'0wj�,!]�K�vS��T���F�D�z3s��z� ��3 ���H��a-qd�3D7�W�O1�e�r�Q��~S'-�|��m:]eW$�̕�=JN2�Iڑ�1�x@r��3�^K��g̀
Rv5ʾuAB%u�^�������Gts��G���
�\%z��ݽI��e�Ԑ���Q=t�r���~���	#���o/n�9��-����e8ru>��uy�$��9�n@ľ��R$v�bI�y��Z�� �y(����F����������aJ�@�:�Ƈj�k�`Z�KUM�m���vP>��ـ�.�>8A`�0jV��WUU]������7�	��R�/������Or!��D�"4�`'�i���Grz�tx����#��� �1{��]�a`�A��鐐0�Z�oi���+;�G"tA�����]?4��4*��S�����*���٠�\*Q�;�>S�$��mךY���w���[���F��9�f���'??��!�.���דDڛbg�-��5�� 羿�}�_蕨�EhE{��Us�-[��rv�q�\$I�^�:#>w_w����^Q������~Қq�f����/��N�P����Em�[�����RCʖ���r���q�h8,3j��&s%0qu�Q.Y�/���ֱ��
�J7ҍ�)r'�nui�:so��t�7�s8|47שy%�w��D��%�p����)��N#�]������&�&�������OBGM"V�K�g`��`���V�<�����/��*MXB�_������� ��k3`���sJs1^���u�APSR�N�f(����j���Z6DA$�)��lko�9N�ս�@�����]��^�\m���A�1!�y��qĀ^-.���y��-p
�t�U �罍.['qV�M�v���x�p����/��y�����UHY�=��*#9�ֈ��I`��ATHH|�M�YĲ@l�${�d:����D(�u������O��)�]j��9�1��~��v��*���N�����<���;��Lٰ�� @���[����֭Y�[��p�?HC���O��Ny��J�'�Vm�o�I.�E�]SfO�_���nT[LV�t��̟�u�v"�z�Gh�4�Ղ(T�rꇰ����Y�Y���S��hѠ�w~�b�1���aa�$iT3z�&DpG��Ǝ��C�����U�[�D��=Z�~v0���M�ާ0�C"�؞;�qz�F}��֙�㎔^�T}�����^��!k�-�Qk�x(���Aif\gy���EH9@����@�!. )�8��±@w'�D�v�mEL4�`Zv����P���nJv	���8&��8�M�xH+��a�rX2A]kk5rB�t��x�xbר.eU���^gh�`2�HX!u��1;Q��gS�r(�"HWQ���[���vb;��/�Jz���(o=�E�����D���7�jY�.��G�)CH��?2���ew�w����k�X�W��vAM6��%��Gi](�e_t�5%���v]M�}K���� ��Bk��8��:��+����&;`�:�Ӟ߄�.��~�����h�Z�
�Wm
&Ͽ�Ge��D��8�\��2Fs�Y� �������S�/[�鵻,6m��=0�y$���)�ɶFu>N��bg�>p�0y��T�H3j�Eg���_2��{V}~+��I5L%�����4i٪�&峳�R�������e3���d���;e(3Hu�F�V���Q��j/�k$?j�l�o�df�݊�O��"�^�ģe;��5B;�ߦ=���$ �Q��Z��O�҈D �z��[�tn�|��E ��ϕ?&/��dX����ѳ_[h�DwKR�) ^�M|��I��|wk�K��� ���E�Z-mK��R^ˬ���!� ]��܅�>���V��Y�pNد���!YM|�Rӳ%���F��}��Sm�L庶�ܖsʕ�+b��R��-��0<�������� D��n��"�3?��������Ʉ`�?�,�������(8n�S�Cx��9s�a��GvC_9&�`+����)b!ۢ��a�O����C�'X�,j](�0�#��B��@�md���@�"AȤ:����������r#���u�CZJ�Z)Α��݋��d��>�1��K�x�O���
� v/��><�������*�x۪�/;�����爓�Q�K2+)#���+�Am���9K�	�{�s�D�:2�Z�ϑmx��C�Y�Y���&n��|4�ք�К��@f0#'��eAi�,�ą���_�_&D��^����i����v�u�1ݲ�t|[G��ѱevd]c%	t�k����r�@k��D(η��̻H�H(�4Rs@�5����N?$�Ʌ)~��&D�k��.��%��K~�B�)/�Ǆ�"8&�;%�n����2p8ȷ�['l��N;����R�����J�]ϔ�8����̨Ӝ�e��t�	D̆Gp[�Y/w;G�dݵ�!:9|π��r�)M;��o׳i��L�Ь��Ͷ��fn{ſ�4Ӿ�B�`P�WJ��Q��\��K�vlͮ�kT��K ݒ���v�+8��W�)r�O��L�����!��	������#� Ӗ;���k%�n�*�R�ޖa���	�]��A�S&�<q�WC6����A�_�k�.��%�urQ��7�� ��J����"��"�#�]�I_�h�=dK6`R���������� ���^��2���@hJ,��L��j�[���g7W�b��N�\^嵉 E���� �I���V��x��k-��x�\����x�!�(.��A��ċ-�ަp0X>���J��(����-���de���ǖU:+ �C+�����o����x��ϥe8�z>��N�C�p����Qԙ�Hh��Rm!��A@ev?����y��l��!7���c�nF�[�G�b���S�@�}����e��u� �۬Q�y�2��r�G=� �����J�8ߐ�]�f���ǚ�?���ؿ��AZ5���~�2���]�0z&�H@�d���:d�A�($��<�Q����d�S���$�2Y����%Qd�|տ�s�O����&��Q���r��=r��G�So��ǹM�)t���O��0� ,��g���x�X?��n^���6��Z)��h��.mDK2]!�� \�>��+�H���
+���.��4�v�8"P���{v+�g�L{/�lی���en�.�2{h�h�H��d` �ik�	�l��֖pDc%z��նWKvd VD	�d��>c�r��P[��^��X��ta�z 4������	S�xb�x�ݬ"�\/��)ZC��D��������W}4��Ǚ*"��������P�y���?C��H 5�2T���4[8S�g��vPO�n��➭[O��%��l��
K�vQ��'�iI�����i�n���V�Y��s̚@'wj!/to�����VN��3����}�����L��&�S6�&�&}��}a���.�>"?�Ή/�����^�&�a'ae���ſ?�[�R~�jB�.W�� :���u�J�E=X�y�vϱ�� ��#���w�*���c�}p8q%�����ɸ�,q�ws���A��$��.)N��|�_ý_ ʟ7�¨��0�b��71-LYB�d���^#8c	]����O���F_�P�ŉ��o9�PZݴd�,��%�g@K!�	V�l$��5���&=nl�Ȣ=��<8%��$Gy���>?�J��\>����W�2Z�i�n�l?D���~dP��r�qn ��F�#Q&��@�CPhsg���:�Tc�U��@i�|��]l���`8����(���J�ɼ&���(��]�܌��W撒@eS���X�^�éufjAi�C����M�3d��	S�Λ��:V��R�p���f��0P��a��_�+�\ �!��>P�{[/��8ѐ����>�'Oj�Bt 3�ŰP��6؋-?�����/��K�/�'-¼����i�K������ahJN�&���̯U|���X˲|6! Y)3]U�MDa���c!�7T2�i�*Ŀ�/z����/�����µ���R�M�>��77�aX��}�j���!Whm����M����Vh"	�]c�eX���xnj��'�Ro�y��G����ȸ�VM��;_��X�Q�Y�8O2�$�t��*�Fר�O�I��ߪ��'BM;ϝ��N�+�AMpj��N^.�R�Yj���xttׂ��)�V���$8)���]8��ť�N�������}�9���[�9�~��Z�Y��A�]p�!m�ޟGh�FԀ�Oq�%/5��+I.NU�ĸ�p�$�i\�p�m!��K�4ʑd�.���8��,I[	5��%"���q$N�üA $����K�>>\
?�f����V�J�JB>e���X�y�O5�獮��˫��/��� ʓM�?$�����E]jZ+���w���%�s/���X�_�#���S�E��ψ�`�Iؾ�mOXr���qS�%NĴ-��Ղ"��`!�V��A�cw�B�|��ͭmn=VL|h��>����4{j���r "~��y"�p�)բ�� .����T�T�у��{�'��z�HW̦ݬ�(�V�&�� ���+���h9�ߠ��6ۋ%?ұY�멤�B�_��n����>ܶ^ɧ*��\��vz�c(:e����z?�o��cݪ�ʊ36�	j1��an�c5�e֮��J"�]v����K�Χ$<E6t��؃<��Qo��S�K3yh$���A���sI�{2�e�c���g�X��� � 0d�l�����@ֱ=��VS����~
�Fc�"i�t�pm�g��]=}���d
Ѹ��
�%󄷘9��AE��*>���(3;U�D�����L+��{kԚ�����L�19E�"G'8�r����]��֪�]���I2�n��nɠ�g��0�e�I>�g��p�7!;M0�%{���5�x=p�ã���\VK�.�N��[qN����M���	#s4͏YXc���y#�L@Gr�*4�|��2�E�a `�	B�..)X�s�yGs�)i�\�U�} H!�wRg�#�+8��.tƄ��\���M�^<VXr}Q(�����V�C�ޡ��2�-�������f�ST���k������S��b���];y� ���/U��ï$�2�F�w�.�p��5A�4��Ů���{��V2�O���#إy�����˼X�z"~�g�����%���S.X�����j�^~��S��':R�+k�S���U.1�bz�S�5b�cf���	� �_A�erM�7����Am������઼�iu��;�;Y?J޽�ъ�riMK������2��l��+ҳ���ǘ����vn���Cz���9�`�E9!>�N�ֿԂ��$z�~C����}sfƄ*Y[<�u�yz�ђ�s�v��e���Y���#	��)H����fߜ��S����Y/h㹔i-ݻ{�wwyW��(��O��z�wu�ϳ�e8jcֻs����b���hp�"π*.˵�="�ČZب�혆,eXf��r�_�?@>�"�  XYxӞ!l��W�|� ?>�#0�i�x�t�$`�-8����Op�"��+u�Hdo�P�7I�Ke�H��ص������q�-k���2��vJ�H���y�k}�	vc�_�9-���l�Y���n��h8��S�?�Z���Ψ��0��G�����O��
b�ft�Z��MX:���gTU����]�d�EU�֖��荏R����P�A��1�p)Ϛ�u��L�Xɱ>�5��w����m�F��xJl/N3�uRwO�]�/���͜�	 \Է�	#5��=�*������n,�)�b�0��i��7D�aXf���\�����-�Nfz�9��1ėo{�D�]a�W8�p��z�Ѳ��m�V��F�J��n5̓#��xd������t�tf�q'��
����lr&�c�+��:�3D~���Fp��
7���q����IT+L.�E�U�>ҡYQ:��K�J�@��{��/y��x4��0M�=$�i>;����[<�f��&4$w�ZM�h��t"}%���kg����Sq4(q�i���Ż��G
(
/����g7e����|�����]�e,���vq��v�!��mA�����je���	Ѩ��x�k~dx2G�X�=���;�&U��)x��F�*��K���B�Ҙ\�J&�,)�J=檔�I��d��*t�TRz��7�Ů����`,B��̼�)�V�j��q �oz]�.���4�y������4�>��q3̕pz��e���y|�(w� �$_�ء?o9`M�=ʬo�"�4ޖ�� Nh~�$���"&LR^����Dy��<B{�IT��Xf�I-j�n�=u����/U3)��B�R�ċtx���B;f�/y�<�1���ĉ�PY�O��+�e���}���G�R��H:��>N���W�|A|�1i�_���(w�)���9�Og{��w�L�<���P�9�cYS��E�\͋RL�h
��K�� �	}ɍSf�eLa��ŵ�F��m�D��yJ��t�NB��y�	X���Ɇ2��cz�V�룣ti@\�h��_�#�� ���1T��6Y��rQ��V�k�5��8���Q�n ��S�(j��[	{a/E���!W�!%*b���
�F;�;s�G3��^��s8#�;��a���d܏��n���E/��pDV���Js�����"^K ��ry�2 }�^z��}�R�Yg��'l�+0�1�{Ξ��ۅ�E�T���&��#���v�A����t����s�����\��sA��"�P"ҳ7�HR���T�6�cA��m2��"���1>o=��+p?�m#7޹_��U��-_�Ze(��&DYf<lTk��=O��D��d��#l)�Y�::���@���_G�s����Sv�~�ds�٨��02i�#d�%�6�KQ����N�+�pD�:ꖇ�1&��DCG���nRT<�d`)��w�g������7=�$�
6O�|� �NE�z���������3�w�����K(ӳe���o������	�[��}��)S?W|����*|{z�$� .�?�+��u=s�O��@W��5n����R�?�B�&�k3�#H��X�y2��*����I�ѥ��`�o{a��@��6ز9�s��}Z]��>�j�N�̔�;����U��ƥt�^�
�<EB j饜Z�p�D��$>HX��X���(��:;�&�:��^y:�"�1$%H>������J&���k�a����~s�*D��R0��0$�q���R��c��`ޅ��y40sΨ�1��j�~��Y����p��ڻGFi-���ᨽ�G������Z"-���ՇƠ������g��U|����#/�X�K��T4 @�eX}�%��~B_�փ�Dq�/����)v��r��O���(�K02K�A2OE�zI�.�ƃ���;ܼ�1���6����@��u�O��x��j�,e�>˱"�b�Aѭ��=��a�$ue���
d?��
CMH�]��9x
�o�Z7� Mo�,j�7����?���Śq�}X�r����Æ����O5%9rN�)��Ӽ^�:.e�\��˪�fx(�Ոɘ	�\���J��`]+8e�x�x���w Wb�H+k�"��#�f]]�dP���u#���n�M5��t�a�)H�5��=���þH���oD6�A$<�;)�hKփ�(�	�y��6����ކ�iot��3��24�p([}f�蓽ԦD��"� B���{^��~�р3fC x�B�f��V�|7���yL�x��a���6��pJ�G<�8@۸�C��;�<�}Ҵ� �OYˉ��bA,�g�
0Ǌ���x&*�Ju-rv�y��{�� K(q�U�i�pf�
�
�K��֔�Q��Μ�!�TSn��ɥ'u�s`Zg�� Fj,_�e�[�Sj�׽D�aՆ���>PCM�m8f٩/���9B���q��F%�OS�F�� y��tb��T�Ӓ�S6��+�c@���VaEQߌ�W��J�2��Su��#�E��a�缵d�j�5˼>��C|�g�� ]��71V~�=<Fb���6C���|�(-::��w���T?�\���-H|���KRT��"D�f��2��.��]�G�
E��-���zqk�Y'�S+�-��v�x�[�)\��� z�P0L���~f�0���c���(�0���ׁ�0ȥ�2�=5b1��Ou_�D�0X��o� y����O��n�ŵ�%>�����@L?�7	�K�r��)@=U�U>��q����UTH�#���uw:H��u��bz\8�,k��\X(���~��^�[H�-�0s�E;��$�0��6�w�!(54uH���EpC2A3��x�&�,~+@���Z�M�:�))e,�nOb[��kbU2RvkJ����)�fa�;O2/�a����.�RBPVWϽ�:��l����A���{�'� ���<�Ko\��ak �휚�=��9ogS�+�LvM(�C�G�g�*��f�@@�]>� H�����]�4%&?\^^��R�Y�Ҫ5��#j�Ų��&��f�Du���#(�h�k>o0�K	U�N&yr+�L\gu�YmD[i��E�W�s?]=.�l��*���zdޕ^L��V�Wh�l�!$9@�_��yi}k�l������A7(0�
fD�Q��˶G���mV
�FJ���:`���a1-���ŕ��&�5;�&Q���s�}2��O8Z1å�"ܩa�AE� K����px5a@��-���{s,�����ޜ.�
�ڐ�_���\5j�\1}����>�>��W'	Q�	h���|~g@(Ϫ��N{Ϭ:G�D���j�!���SvI�aW.�6O�<��Қ��
�����Z}�0�z�~�p>��K�SN�P�1��X}hiZ����h�	,�W�k��-��#�b��z�h��1���0�.�N3�J?�*x	3�(�C�ڂN�xg�Fm^��l�\�t�X�&(��4�]�����o0"	���dh�F�B/�T�o�_]�}i�D��@_8=B�y�;Me����r���Ĝ[�3�M����l�,�8���.�}a7��������l{�vB�a92����f�kC�Y:����.�1z�����6�^�O�Аl?����J��r��d��6�V�F�»􃡅"`!���\�2��+�0����	�,�߉��u�7š��w���BN�N���H\�6|��8�[�-�?=Gj����"r��Ɣ7Qh�����Z��(�"�:3��

6��(�%�D2.�N}@о;�ƶd������ߧ.��	yG'+��'���eЪƘ;JZ|$UcJ��fU�� �JŸ���g��Pr�h�.�[ �q��-R�mV*�]c1�ud��b��l)���M�oN|:�2�3�����7��L,�<2�-��~�2�����J��x�w�q��%�2 F�F= *55 �u�1n��P�M�|m �QTW�ۅ�����t��8�ѫI�e�_Ö�s�� �fi�� ��@��E�(��`ٿӱ3jޝWe����^�w9��Wm�\�]Y^���9�`��2����=�b��ә�^G����8_���#nNA���Ø^sms��j���F]wa��Ѽ�����O����c�� �n3�Jǂ�C�\��/��[�w3��C�x+�p�x����cp+�w�����e�
��NP#���Cq�r`@:�9_b��
Ux������h���'�+�<1�����lE��g��C��P�u=��B ��P���f��u4&��ͳ�s˪�A"��בþ�j\BјȜ҂P���T?�����L�|�S]A;����)��9h�X�B�5�͑1���(B�e����Q:n����2��#[����b�ghz��"���4�Uf�j�N��]�sT�Mq��c�渟 �9Z	f��3��X����;6�C��0��$�g�6�8*��$ӂ���D������2יP�P��V���Ǭ�Eo��8��6�
N�l���s�.&�_�..W;�_���ϝ�E݄��,"Tm:Z�J4m^àӜ0�%N�d�B_�yh�]e&j�	�迭��t��q�E�������^�[r�FYf�hU����!�þ�Y��/��쬇o��
Ԟ>+�_�[&g2=i]N0	��魹0�]^77�,/'�t����yg(�آlg'e�����!���/beR���W|հ�A]��z�M�u[E�`��ͦ�^�&��F�1��ݛfp�l�����4)K*
�!���+W�w̵|~MwΞ� q �&�+߼K�A� e�gj�AK��G~L���_t@茒�-s1��F�FA�V��{�a�S�Ȗ�|�N>oD�8�f{�`�ݏ��lgH�4��h�O�#�z�A>AYNꭐzA`�#�oIyyJ��-�Eɍ=��%���2�1�_>�L��/ZǙ�nW6��Y�ʭL�t���6w��Z��s�>7R��EAL�};[ɹ� S����@�b��j*^��u�f
���}������:{�&6r&s�����c��冡��J�ĪK��h�z���|����`�sHv����M�\��; ��!m��Z��`��)Q;!c ~'X���mӜj�@�&�r��b�tV�=���,g�X�d��0[E7c絽�
�eJ��U~3��ovqIQ�T��$&4 x��Mr��0�ҿ8Ӯ��� ��#^l�_?h>DUG	����ϕtR:]Ҙ�	�-��q�8��{�1G���܍�;Ñ�h0�|�ĭ�л�
K{<���!y�7����J�Ԟ�(e}�����?p�EM���ga�x�iRa��^��jH�����Ȳ(�(�M��_�,��L4����1��Ǌ��J��(c�I&L,\���0�Mb����p�]�����2p�"q�Y6k�>����a����v畡���Ö�����G�Rm�)�$�F2v��f
FH6�i"9{��"����"�N%Q�}"�ύ�Ħ�i����W��|���0��Q
RY|_�E��o�7��4$si���t����t���c�Śp����Ig%�i��]�ALK?�L(-n��>�"��F�
�O�K~�.�}�C}X8%�h1҅.����j�K�;@��
RCjx�;y|���)���NIs��Na[��8�0xCm����_ 6�IV)3�T�8�dabF~q67̑�%9`FN������*����{�+ȧ�`�o5	Ja�	����Y⸍9��u�w��DG?��9=�}Z��ki��R��G�GצR��)�B�x�+=1���N�^�e����<=�+u`��p�f�
�R ����|3�aB��U-T�v���p�֙wڿ�;��#�.y�j�`a�u�;��#�Mtf֨⟜������·9l��*��>I����[�t�Q+�O�n&Xl�MM������UĒ{l�V��G�f��~�O[Rp\�7���~�6JQ���Q�;��b[��0��?���u+���5��1��!P�0�
�k���e@���5�<C� �S`��'�0�#c����1�R�^��A���?�2c�}�ye(��ҕ����*�P���#M�m�8�壢.	��G�H��4�Z�C�p��-ڱ�`W�����*�����ҒGXvI�O`�P�{�7<?B_���Oa7�$;�6�S�LK�/@#�H^*�i����5ޙ2�p
*{1��6��}D+\yX�1����.�ɠی�M�9�H�Z�Kp���u9�Iok2�r4��#��L�,P��9��wA���%�G�̗Z�e�E#s�v���R��k΄YFqaw^<j�/���8�7�A�������'�D�0P�5��sJ��6��%��wOvd��3+A�1l%.�W��f�:���=z_%���!�\͍���tm
E3��TN�5u�ۮ� �Eb��Iz��)��M���k�p�K�uM:Y@�����~��gxV↹�5�k{G?��ff������$�:�	+p�?��N�	5��(��3â�N�-b�4�`n���	:����j��>��	ɏ�,Yu�	����vƺV�Jxy�Q�y���u(�H®�-v����V��55����9d�V�S"�ο(���Ҹf;���f�|2�v5:M��au��d�8�+��	�D�J$��8�f�|��	��u�����+�x��7��2��i��bެlQqh��/�W�F��[�W����HL�H��ժ1I c�EFi��͝y�N�]rS~&9e#�w" ڇ�.h�O|����PtITם�o�>ͪ�vb��\��Wv�
�h+�bY�P�ٽ?|�y%@\3��<΍��*[�|��->Cn>-T�y�d�U�I{�s9�i�#h�����\e���t���8�-U��$�dP�^AwR��%�)y�6���c�eF"�tv�v�1ૣ �2	Ӷ|�s�8\��y���e�9��){aK�F���%��)���'*
;���s�ݶT�L��xV3Ԍ\F���ȯ����m���^+�H��T�P�4#)�p�Ud 9Y��X@ݪ�����)�{"Ʉ����=����d�5��d:Z�z��iwZ�pxB#��Ȋ�I�IH8�����x8u��98��}����f���Y�>Q����ua���`.��L�*FęV��/
*�D�����`	���_�^T���԰c<2�j[�С�Z�f� ����
=f�:3V���[�|dS �j����%�%;�ڙN�]�X�f33���YVG2���8���1A��d w|�!�����ڌ<I���0�
+=b7�w��?�q6�Ń�Z��yॏ�/��h�1_F�^���2�Ք7���&�N�ⅱX��(t@�f��O�7������75\�p�i�{qw� �0���O{CN�W�8U),�!��Da���Zݳ�W#FtEuP��s�%�a�7��{3��)�y��YEQ���l���#��=��O�첌kOl��&��8D|l����I�x[���'7���Ƙ�bES���3Ԇ�1�[�E߈��G�L�ph��En�0B�Ϲ�B��K�enZV�bW��L�w�ܞA���J�SƏ[�_���@ ��P�j��g��;Ӹ!D"��M7P��ɰk(��~�һ�7��}-��/��Q�?��2u�J���^~~ �VlÏT�]�cJ�
�
���V<s��C ������|��_z�=))
u�����U�R����_���J�ޚSZP�)�jcr��q��{�C���Y��`+����s�v>ս�`>%/���lﯚ���@�a�bOlv���=����ݒ�t���=υ���R�t-�g�%H$,e���]�L��� �N��N[{*�߁�\�l�!�G�d��[8}E%�4ߵ+`F�s(@ҁ���&TԎ���~�߫l0���P�H�
�8�������n5�Pe
�x`+c��1y��5T+�s�Ñ�6�Ћ�q�U���מ]Xe���N�����~�9�ߞ���.��iF�Ќ�E��k��ܖՋutON��z�c�Hq̀s��Lg�9��kp�K��t=j
�0_m�;_���&�fJI��G�
W*����w9��5qr��j���U�`r��x]�r�	�Q�r�6�s�a��QO7��;��t�'����Ǘl���rsDHWX�2���B����Q*��	�@���gȒ�A�h+!�YG
��/H^o�H2O:�>�eVA��YyY��8�� ��"Q���D#O%�f:��v���p,�.��7�Z�A<&���G\3��*��`KG���o�l�AN(T��Hd��RnfC�k�v��G�-��p��Kv�t�B��)W��58 �V��'�s� �e���)wx��P��eVg8)�N�u4���r	*��n�+�2���+q��E������0�A�͡�R6����̈ρ��KA�K���2�US�;8!R��#잽��6�s;�?�������T��EV1��e��r@��Th��*c.�{^�A�cbD�;���U߰�����.��Be&��[ۯ���=��~��^�.5�� ��{N��~0ΦDH��;S�^��ޗ����Ɏ�S�f���⦜�����)��4=��]]���-�JT��m����*�����6'��&j�����>��2E����Ayn6�6k��cE,.Yιjd�
��ﱌ�#�ؖX�%�x{�Wg
@���v�G �}��?2��[In����#�C�E*�s�1���"K���D�h-T���#�ǐ�ֵ�`�r�q�o���( 	d�+3��]>X|L�Q��<���TW����x�7�
�2��J���n/G r��	r��+���O�8،F �ԙ;9�M+�Û��L@�_�/:GDF�1[��rg��ɨ�'��Χa`�}���t�̓b8���w+T�jv/�4"��8����}���6g���w�?��le1�ŗᲀ�CO�ޛ�_�ld�y����d�;�D܆({HOP�w��B8�ݜol�"ꔀa���`S�I�uЙ���$L����j��V3����U�^_��k����k��[+�@��D�YԲ������>���'�P�]h@���?��o�y��m����掍����KA���-�z{�g�b���]5L��Z'z�}�@"�'Z~o��[Aa�]��Lz�i�)��gW����6�tx���R�*�G�k���zy�A���:yNX��N�Q4d����:9�f;�>�L�Ow��#񧁻?	���lR���`�o���2�q�����tp8�8b|OQ���Jh�%�^�|�������`��Z\�RZW�,���Ʃ`�v��,��O���/y�i#�p�Dt�m�RQ�����J��1s�Δ���
���õ��m�3w9"/�߲�K������K9���j�'��?ܡg�U�G��v�m����V?h�ڜ?�>�á���S�U?��3�G��Ƴ�0��c(7m�\h�c�k�Lr ~T�'M���#����^�t$plz�@��4��f0�%�&H6O:�N�6,Ƭ������֯i�}��E7���L�7e����s���k�������U�D!ȃ��A�����䙓������f�y��2��	R�NDa��6�g��{��o�8�׵��8��Δ+K��a��!�=�d�p{��TU�@�/�3����N�e*wT@F՞��[���g�7�X���d����Xܖ�{Uw��_*�Q��x'U��ؐ�����$fwtA����Rޚ���q�g�X�m�:I��V�
�^k ��;�����.y~��>#an>��"]����u������CJ�6pE~�����=���A��N�F�oo�uJ7����Ӡ�,0�}��;�Z�i!�Ѕ�"�ӯy[��.c�r�Qs*�OX��P�bٶ�~up�����	��k�l�4�P~P �6���(x��.Jx^��ʑ0�ǈFT�C�MI�<�\
+��1ȣ�\<�_����@ߏ��`�=�/��@Yn�G]�fѢTk�rZ�DH�*÷ɭ��º;�r��4�v��������,j@�mW��h\DK����<��d��'�ˠ����ME���E���.Z@��N��JS�Ci�������7�t�Y��Vwb��F�+R�JU!��ִ���0�H����+�^Gw���,Lh.�1���8o����|��=��~X�*j�M���܊(b�r�&\B�N���@ @?N��5��4��C���Y3��g��Ȃ�Mګ�-�1�s�P���6w�+��UF�D�	b8��4F���V����b���+24F��wq�B�<5��C�����+@����Ś�~�L��#�F�� �A�mR�]=���!1����(4�+ԍ��ά<��x�b�Zt�-�զ��J*�ح�83�.;��F�������=�%��ސ�=��Kzcbn5%�b�ۓ���Ax���i�c:Ĉ'!�l���|� p�=h*��z����`{)HZ|%!8���=:w",Nqt��q��s�V���#��(��tz��Ò����ʗ��R����.��p3���,�4�t5M�cz#�+2��KwFV鯟����JY���g�/#����Y���LTC@��A�vG�<C��D?�QL�F+y�������]c�Ac��d
����b���x/\@ɯ�y�n^�89�B��T�����Ol<�tĆ@[P'C]L���&K���<-�R�y�c�ȝl]�*��/�F�DlQ�P?�^Չ�)9u0���2��-l.xO���56'�)�F�
0E��\�dF��7�c; ���p���I��6+�� #	(�zi~��H���Is7D�ٚZ]-�~ƃ�Xl� 0�'���4hQ%%t�?�a!�|^m������5��>+5�>"�D�3F_Ld��Ao��y�4w�U��;
WF.5a�s����� u Q���������͵\�h>R�C^�]s��/����̨�1S� y9��j��cʹ-���}�I8F���)Tx����?�l���i�
�ت5������^H:!���G�����U�<�5���]�J@���y�~��Or�l���!7��8{��4�ƱN�4kȱ��"�]!�,5�1�M	H��i�縢y�kZ��q���������6�T��G����2��N���(��I��>�i����vQx�G���d3��rTP���#M��U���� T�V6Ăq��į�^2N%�k��6�-4�\�Ζ*�L���䑴4p3����E��ըA���B!),Ĉ�˓(\�0��!(}Pm`-���[�
Σ�n ��ʷɓS�k��iU��#��oAl�9&�����0U�
���S5�O'�I�]��r�?uE�<xċօ6.L�(fa̩H#��`R�0,�JVF_�!�Z���mU������(Ãm�� ��1+���sb�:��J��a/XMe׿���!���fx-�<'�GlȀ��xE@,m9z�&�EZ��e� i�b�tjlk�L�y�kn�k {�(A�m�*�������3iJ���lM�h
p������]ڙx��Ii��>Q>�]���pDAk�o��I��7��O�/~͝;�H]4�{����Qq�~���a�i7v���.���փ��~٪&�n��m�]�q�g�?b.3"�iL�� yh�
e�\��'1w�3��E��no���L`{�	�x�����h�`�b�u���?��j3H�Ic��]S�'X%@�r:���db9� yb�Tt�z}H�K�E|��?�R/�5SC���)�OX�ߦ��CU����o�";k0 �'�$���<���lA00G:�If��~��;�x���B�UwrPM�K_(Ȱ�5"84؅� ��$�D�c���Y��;G_�ԛƌ}��O0�t��R�"vwc�;# /�`�r߂�,��b��l�>O�`",����1�0>x�IB�1[�ǩ��Ò�%o}���nhŁI+��|p�����I�������!Vi�� �tћ�w���E$Y�.p͜�u��ӗ�X-(�Ǳ��-"a���*�Dܲ�1&>0�Ё2Hl�������2�)�\�=yc�ql�lgl���d�w}ʖi�m��;�'3ԯ<��k�����h����R�fK_�z7	�gZn[	��	vӷ�b��b�n'�� 8p��ls�]FF3J�q��=���E�m��l���RM��WӔ�m1�~��y�4)z�g%n~�Qu`U�R�8(Ne��8R o� wq�cy���D��C˶��`&��c�}$[�85�`
 �ї�L�U	�(oa���[��g�ָD������N&.1���n���-�5���YD�!�	j��J�f̭��yVͯ#�VMtA5��X\P0f״*f��Er���������Y��]HSK��0Nf�v:jR��AO���x*ul��P����:DzU?�#O�D,�j�Rj*$��A�Ќ�?�*;�+���<�8NɆh:U�0&`��{xCu�ˬ2�����l�A���_8�pNӎ�އ�'�9Dm�=M�����F��������c�f���n&g̒ݞ���i�B�����+�<�~��������^��`�1���S��� ?�kr���<�R"�s.��R���\i�,��s-�};]�8�x�v
��N����:�'Ą���%3�D#K9�a܅6��r�\7[�U=��*3�ؾD~|����I�`�4�P�wY�#G��m�p"N�Y<��4k��l�~�@�V��#��G��������E7;���S�0%m0Ȗ)�/�!�t-W8F.7o��s��P�@�
�`_��̢��f��QZ�!����ƽb�@��9<\�4Kn�� �G�%!d8��,O�����!������y�M�a�@|k<�.6�"d��
��$E{��t�C��l](������9e�����}���d({�m����8��u�^���.�!/���u'*��P)?��%�Z�&��t�a�׫�o=J
��|o�[�^����,��j_�K�3	|��[��H���o�nD8�?�m ���g1í�8�/q��e�!}� %eAH]�p/o��]r拯�@����3��y� 4�%�����9�Pc�}(0�ɏ��x�#t���������t��"��/�j��0Zp����6�'���6*6BX�}SDd��v���n?�7��p��{VѴ+��^�Ϯ�Oϊ4�m"SyuJѧ�="i�LB�R��)tĆ}f�I.#�\X�r>H�����B��)�p=yt6��"3�(\��9���v#Qs��U�?���H�?�����a�xB�-@�n,�����5�6��p-�5�"Xv�CJ�<X�O�Ͼ�mb��B���<>��?:���j��V:�|���v�Y�"�O���op� .��F9���߿$y�6�_��<^�?L�M����
��3��ǘZ������;�;#������tt�󬮩�������tc�ۛ�L�x��g/�2f�Y���5C����E��t8� q����8et��-�MZ��?�B=+A[^��_i1�9M��ots;�Ɔ��lWR�Mw�R��6�Z�Z�a��~�^�YX?�~A����Z���L�X�1 �9�cD�J��;O��+e��D����ˈ���V�rWT�A��W�t���:��2)�00Pt}a���.�q�`�c��T���Om#��z��(;�p�!���e�8	�"¼�
M�;s��ʙ���B�����Y�ä��0������%DH ,n$5P�h�e���y֙����̙ڃ���� yS����c�W/9kk�\���¦���\t#�m[�=�X�j$��IPI�WS=r��%n�M�	yU�5�xs�]��x���N`ӗ�T�Iv]~����u1�P���W��I��nʈ�e@��}w��iԑFb�sD�_5���z�C�����}��-Z���JCt��[�X_�ߜ�&�]8/V̥���x���\�Y^2H��\��izK}�<"D�,`���:\���6z'+�H��əQ��Lh�1��~����V�3 NdG���]���R���c�v���yKe/W��\���8�,Ђ4^��yBx��Hee�H���}�8�L�E#A�jC�7W�ʃ r]��L��Fq�����Rܨ�p݌\��1q�W�n�]`��
��x��c�w@��2�T�I�	��&�����D,�I�mg5���W�����Y�3 �n��N�\  ���p�����D\S��?;�(��*��T��}���OH����<���9�
;]��>Kb�y1�j��6����e����R�h�+�`@[�`�^Z�Q�F�k�!��Q��*�Y���)FSp��Jn���������0���CPg�ѭŗ�ۢ���?;�J���g4Z�#��{Ym ʹWz�Zg�'��&��t5 ���Mj;�qɜ��h���y��'�0���wn�+��>鱂��J�D�*�t�L�ž���V��
q�8��sh��Φ T<�G�=X�A�t���
�s��&A̾4;a����[G�5��j�~p}wM�$��o�����k��"������LLzԬ�����1,T�d�[�pZ��B� �f:��߳���5���
��(Ko�	���ó�� 	'k�)�-=�[h��wՕ�ݺ��G<7������ł��v�]ߵ�Ő����F��4�B����>���B��XZ�X�ӚG��-�����A�&`��ѵ!d�6���!�b�(��I�;��XA�g,�+TE~�+����id=]~4KZ�"�K��3F�m��e�B����#w���Xe���̓�ˎ �$�.
k/%�c���^����	�����"�>������);�Q�$��`���=����h���.? I�8��`���͋�Nm���8��l�q�Uz�4lE��T�:+]�qm�b[tf�J��`gl��v�w`��v6��7�95��k$?%>�ſO#+�`�?wo�;��]A�%f�"�����\��3{C�Z�F���d����9�*�s
�)��q��})��;ƾ����Lu�'�
�5��Ϝ�w���XF��V���9{V���_b&�1������8�������ZGlCu)�n[�#R-�g�9��[�\a�':Y�'�:���=��`j&��K#��z��zoP�սD2@	<؝�"���<k������a��z��B�@AJ��x��0��I� ��^�퍇��(�L2{	���޶�<X#�*h�9���k<�c;�W:E����jQ�v��ә��Y��.�Nx��X"d8���8s��"�#;x��l�-����uv� ����j��*��Ny@䲟�G+r��DOX2���?��~����	E��+��`z�\�5�I�4�C�h��k^��ՏX*����$�@Wy%�B�'Z^����v���QN�&�l!��&s�x�Fv�?C&=���w�����h�R Y�����PUH8}��0Ƀs#=� ��0Ր%;��=�K�vN����u�.s%��~qQ�Q����%D���?���5���+�Ǆ�
�){�-E��'��i���H�+j^�&���&JM��	��n��9#�##M��Fٟ��n�e�N��F�-!d�"Ў��D�*!j��ڀ<���xf�7A�����َ�f�8��H�O~��������
v�Τ��ZUοIp�`����l����t�����������T��X=*4?����0���l�<!��hTK,q-{�)�9`��X��������=1x"T&O)�{�k��!u�#Vj�	�_�Ш�ÃV�1ږۊe\e�9��HR��b}��z�e��Z��Ct!�6����u��vƉ���y�ו}T[.Xнw��]j���
^�)`&�����x��!�K3�{W�k���{�Q�����v�6Sױ��w�.�~t�~6q��� J���U_5�e,��1c��ǡ��K��=�^���`����x',���?�.��SIU��}�9{f������(�����!� �{[��h],�� �2�
���3�-�#����?鿾�Rw�h�9�
WX��x|�e?��\>��5
�s������fv&��XG�����tO��|]��24��r���5k��#� /�6�2���ǃ���r*̺��f�?.z�J�B_�=�Ϫ�y��u�p�n����-�*�N����	��4��l�FX~�����c���oػ�܆�jŎ>d[AGh����`vo/�) {9�`u����w��~>�%g��`������~6Z"�3�<�#�TEZT��J�$��,�:��p.��^K]�Mfg��� �@��������T��f>Vw��0��7�]o��}O�Q]�'�_�.$���?�ܞr�l��r2��5�c�䬄������yz�j�9�뻆�/�N�A�k�Id��q���CpU���v��y�PM�c=+Ơ,jせ�|��yi��Vs��&wRs�8���T���@^�����<��Y*���z��+�מbI��fV����b�J��9V6��L6�6�bNL�y��������rP�7���Xf��>�����%z�a,����G��k5�>��W맗� y˩GP�Ba�M�m�N,Vf��莓`c�s�+6ҫ��p���_m��v�������M��7:�`-���m��\mҞd����q���2�g+X����7!�^���6��AEC�V���MQEq*�Z�I�'v�*㢙U\�Ŭ�!��w��'��{U+u�҅�����Z���J3�0f��1S#��
��2Xa�\����/W�\ӠX�)�M�}UnA¯&�M�S����l� ~����[G �t���_��Ijb1����y�!e֦�Xq�B�n͠΃��=C; \1������~�m��)�X���pC��G12̜��d���i�u�r�L  ��;�?r��[��kK_�r�J q4|XTZ ^�X��Kp�ƴ�����;�z跰�{X8J��� �x���"��״�킋��$�i����$�Wx,$�K�����j��±��,=�v)�Z��X�M)����z㖴�O��0WxE��^͋�G��_�´	�fN���i�ͦptxpﰓ5�CA��q[�c��aW�v� �Ë�a#���m�?L�**�*�s�'J-<8�T�3�w���r�X�m`+=��e��x���rs*��bg����5UF�i����w��,D���-ߛG��f��Lgg��3�P���j=c��+�ؾ6�vqL^���*ϒ� ��J~K��E�T��-��~8�e>�D�ŽHq�ƻ��z�̊���uE}iuP�U.�l:j��J�b���X���v7�D�l��'n�g;E`���Uj�P@,4�c983���u���
6��~�0�G�KG���ա�rG��a~�1l��ߚ��I�C[�X��d��DJ;��(�O�
$Vl��/ ���������z��<1k�s*����L��a��.�jp�Z�a3�����ŘB�y�[3-������(��B���y%�1��x�<dW2Šeg,�m�����iT��.h�R�͗>^���~��(Lۢ�tum�
Eۆ�~�5.](�]�Y?�P�]Ltw��죀�jҲ��y'���6N������ƀ�bi���X�,�b��*�䶳�W�t�y�4���T"&5�

�!b��!9K���0��W��g,�7R� ������@n�Qݾ��l���ڷ�(15iZ�C�G��m��`�j���b��Gn+x
i`E���ƹ��BeGg���:����f�q�q��.����d�1z��>�}����&>��h5�u�$�f[�OMe�#m+_�ģ=����Q+�ވ�"/����'==L蟄y/�u�����?����w���je�o���^�#�������{��e�K�ܜ��X�k������[����F:��j�~��X|6�"&��J:w3�_�QzJY�]D|F��良�N�w,(b�HC�3�r��!���.:�JA��r��AV�pm��4}~�l�S��Cäo7Q�[�J��ۡ���e,2I��V��NLL��$�ᩗ!	��v���-k0wX���'C}E}��w�_z�AbmQ>Wqɺ�4���@��$05l�+ �R�	$
����C��{j���T]�w�V4YKt��t,��-���U_^�Z�>�DFV> ���-N��� �cP�u8f�r�E�Q�.Y%7ZK�U�f�z�Yx�T���YC�|e���~A�u�	t�"��k��bD���a�������0�&�RR��ե��V%����	�|q+�bj ߨ��{o��J��-��dt��0Dh�B�)�k}�O� lU�!l�M`7����	�x$��M�#�]&�P�4{��)~ ��1���g>/��r$>�����T�ęy�t?�Q��;����c�0��1r�0۽E!��x�q[�DNo6�1�u"v\��\���҂��|���5��'t�i @�ho)pب���&_�#t+�3�$J�5�\NST�u31 �P�&_a��N�h5�T�b��S}4�ƣ��HI$�vjf�tą*�I4�~(z�w"�1q �N�:,w���ҁ�QV�P�-ǿl��')��u�J��zG}���bi���(�ȼ�@����q&Z�����ڎA��J�6 ~)�z�V֖[+;��dk�x"�����+S��Q4����&�����`j�m%�&��<R���,�ˌE��ӻz��uiҒ,ĤL�g@�A~���%X#D���/M�l�4=JĀ�H��
Os��99�����D��?N��fRwo1Ь��J{�V�mY6D�*&V�\_9�OF��r���p�b`鋞%�B�ױ W͍�x��#]	�^��hw���·�@,���ɗ�\Q�eח�:��]}O��,�V�H���^��L��i�ǋf�O�xtd�I>X�\�6̐f|0K��N-��3��OBռ��j����R&�d�Enf٧�:��u���̌q�+vf�M�7�慊Ė�K��F���B1��p����[�ۅ�4���R�.ģ��@�����5�X�\��5��T���g��?��7~BD[�^I ��Eԇ}��T�B���U��6B��{5���N0'��'��0E���
2h�k2��Je,M6��vj~��O.l�m�7ӡqTQ,inG��+^.̨�f`�җ��D��J��i�iu3���,N�5�j �Oo�3�#mOwmBKWv#z��&2m����:'4���@���a��;V �d�Q�RP�H�S���a���2�t���xBjZD�_$��}�2��豄��s�p
Em
�q&*Oz��)��`z�fUx�;]�-�e�z��M����E	�_�Y����w�nЅ����>Ɵ�����]�N�Gk\*tFhn��Q��L@%�m�0�C�%��b�\J��)�E�J'f��2��UFO����$M$��Z]�d�}GRm����+K*�Bjm�}+i����w�#:!qI賊�-��l������~\�l0= �=K`Q:߭�%
39{\�yw������������I�Ϝt1����v�cZ�h��KZ���馏�Y(~��L�hl[dD�c�q�v7��_Oκv���ֱ0�$�����i��s��Q�%��a�^���=p�XY�������G��yDfXB�1�f_�Z�����V+;��N=�89����C�K���j��)�ɞ����7{�̌#�T�#i;���P�������]��T#���3^����`��N}VQ�Ic�OO|�'uz��^Ud[ײ\�0뉒�MwΘ5*�I��Q�=�o|�j���h��?�/�@�"�����=��-���9^s����&�T��ׯ芟�gk�,Ї!���U�[	B��/�⃬��Q�W����� �P�Z*O�E"�F�;�o��U�,���ᛞ:h����-��K'�6��P ���&�-�/�ܮ5K��Í�2c_��g �X��$���d��P���8q���Z���Q�Β/��},uA��/�>bB� ��(hF��C0��ov�9�4|�ū�k��xAS�Y6�����4�}�!�Q�:-���C�s��d��'���V$��[<��Yڥ��/oW�:�ߓ���0�Z O�9E�K���f�Lc��&fӸVvd�nlm�Y��TK\w����C���ܜ*V�8���׃m��Q�#c>��ld��W�!��S3]F��[�ڞԲPR��Fk���^�d%� �9^�ڞ�-¿���y5�b�1����A��D�]_8����Y�gψ���qLpE;��]��&���p�9*DC�E$�m7A,L&]x�[�4&���Bx����'�'c� �>y޸� �y�˥�c����>`Z@��{��삾\�m��s�`k�QRjC�@�&"���f���?����5�_�$*$�G��?�`��Om�$���hd��6�b m� �DF�k�l�);�V����S"�0��p�4��'����.nK�9�h/�ָ� ���a�ө�HmUc�o��-k� (��A�K�_u3��ܮ?9�a�L�q�;Xۭ��od�L:�^6��ZB���7w`u�+��m��{}��K��K"wHk<TJ��*���TPd掆�]�j�Z��NhC�\��:	4J�q��fk-�o�x��xO��y�EU�,t�PG�'Ӽh�n�9���{/B]��;M��s(&絲���F�?l�U8�p�c��gȜMNbe�ߣ�_ۚ�n�*�}��'��٨8֑|��G�@�=�`]��:��-��C��}-ʫx	YL7�z��a�5K�&|׍F���M#���f'�����xy�`����j�c��q��i�̷N�<�Ձ�RX���f%ȳq���u���l8�Ў=hB���}����\�\���_Kfmp 8�-����:.�&��w8��L�p��Z1˕~�����;�u/e�.k7��H��s�
$sy����򽿐�yק��h4?+���/�a8�y�b o�����!y�]�{��R�I�eLl���WxqK��3��!1��;d�uĔ|�L$j�����$�6g[�vab���
�1����ǭ�̆��n_2��~�__�R8���+-$�Ʀ��e�_2@^�TwT7�-�(���ޅ�t۽�=}�t����aѰ!�@nu�`K���GP8jփ;�C� �Jߣ:d\ݰ���0�I�N�I��:v�)y�.t���ݩ����|T��F�$ZR37!�$��3xh�Q&q����(%���;2�:��Mw��r�6B8�}��/��,d9��n���{�c�z6��|�����D�b�g(�Bu1p
�e��,/��jZY2P1�M�L��`9� ��7���b�2��j���4)�Z�~q5!w�z�_�P�e�=3��/������~��+q�$�P�Y�L���{�-�y��S�G��6 ��O�ZAe���nO������K�f��e�is�D��"z�fs���A���/N
Xc��.����t�������d�y�[��l�G_/qł�U[�*ʗ>^B��yUݹ���U��ܿy� xe��!��v�la�A�x��Z�t��9�H٪�۾-�:J 7��(v�a�U����e�J��5������I=Re��y�8E�prDrĿ�瘼�2k��5 ��7j���,�b�
���|�t��F�Aza�b,G�lʴ&|z���'/�+d�#%�L���X̠ȽLV��{�.[��f�7 闂�R�����-a$�_�S�=��{p�,�/L̩�G�a��k�WHi92�c�������$�do.9�,5z�������.�8����^��Y��5�VI=a�~E���Z�W������M��PZ7�<f��V��N4��/K�&�Q�٣�����:��P Γ
u�$ż��0B)Ҽu�=�?�����Ե�i�}��ݜȬ�@pq��z��6Y�b�#�uyJ�&v�є�r��,SKw�-�Q��5Y��s�*�;ר�k�I��M�Ϳ�:(�x���"py����N|���(�Dv��o.ws����z���Oe���]z���5�"��D�%pd݊)��\]-�Y�!�#���S���Rkko!��<���-��xG�b<��ױ���4�儜M��eܣ>���0���e������%���%JҾ�a��?��nC���q�ɪ�n9�]��-�ƖmF��|���РzG�z����So��F7��� jF��B��qP�x���q���f��2�"���/@c!�`�|�/���&�Է������ѵ<O��8�X�C��5�����E�s>U�O����Cq��� ��+�!�q�od��+�B�#<���3� U6D��9�CF�+O��a 7~f!�b`��"�xbŕ��r�&�r[�4�q?BI����R]Z�KNQio�mZx�|�sʡ�~S ;��b�c��]���.�ny�Rn�A�	q��&\��ƀ)�A2Y�ސ%Un2��K���k��buM�"`��ֶ�Tٞ����[�5a�������	%�F�e�� ����)�}��yD��Z���d:ʤjg�K\+��ϰ\W��T�2��������8�_$q(�ȇ��'�jC��Y.M�}
^3Iqf�,1���H_���(@""��W ���ۮ"Q07!/�Sx�e�hK|m��(>����{O��PVb�z��:�.2o��^4�)����䣠ӱ���yzeP+�x��E�������4< �W��_�6s+o�J&�Q�1m��3/;��&�ϜuCL+*}����K��&�gY��b1��V�a������>�^:(�jfg����ܒ�IW`5��L>|[mqF��ϒW�����$Y�G����rQ36�D���	��;��a�/6�C��Cܢ�u< ^;�{ʹ�o���:�+�5�U���,������*�ͺW���?T	B��9.�"��ݲo��ߗ�y�oC�����d��{�b<�������SWs������ޚ���¶����A�@�/�B߫#WϪ�U�ڱ�u9�@v����f�f�J�#'�$fA�*�V���3de>��'���6S�Ǘ|��¶��Yur�Z	��^��c��-k�A%x�6_S��8�T�]�/�d$���BQN٘�l�S0g��-l����X�(�O�9�(��r~	ѭG��XBf��)ҹ�GF�M7�r��y������6���`A>��?<�}��R�-_���� �ٜO;��$C��X���Ó���c���OQ�� v�D��Fd�^��~,��Jk��=��a]b�՚��H"A-�9ږ�5=٦�퐡-x^B�0x�G[���=Rԑ~�el��ĸ游����Ut��$`�#�y�\5���)�I<"~*Y��D.$���`z��ӷ�/p�����<G�����aK����(�I<�eoN���]5z�\b�l��ӯo�8���uE&�v����u۬�v�bpp5�,���ƒ�Έ�W�h]��²���ۓjO�O�K˘���_��')���2G�9~q���,7�+��p�6B�NL��س����BUA�f~ZpF:!��O�PV���N�'����R��*h��z�j䈶�£���@�r�V��;���k���H[���H��f��й��(p�Q�N���)S�{w�2���xl��،�pv�`~B���SO�&���1?�����am�,�w�b�X���u��.�T���p-�t����ʱ6���k�Y����yr��?�b\����(>� ��R7�1>bҗ+��[�G`k�J�Gp�1��������G�¦�O�ͭ�Ry��\�����<��K��6��1�&�9�U����K�P�Y�R���,�-)������di��`��<�Yl��,�����,����)���Ν2̀ wJ�дj��s-V�>�:w3��d
�v��Pn��y�k�}�M��1���L�c?�����8t���c2�񮷓���ي�GqK
����-z;���j�w����]>!)���8�hn1��V�JĀ5��b>�os>�a8�>�!�;i�OK�T�8�B�N�46����w$D~X��N�K5�c���
CL���!���`�k��>}�5K3���ŬQs"|�Q��8�e�k,m�r��/z�[������D����q�A�Xc:>(�t�����'��Q�Z3n��:t@��ݹ� Զ*��Ձ�A���H7��o�iw���R�:�/�oz�	;F��y�5��v�D�jh��8����޿�N[�>�HU�x��	4#^�1O?��wy�{
X'eQD�E�<�c��P]�+�l�ךD;vI.P����"�8A��פs��?`�d%Y�!E(1�)+%?
����q�Z�V�w�Toq�@��Tl��o��e�U	������Ei�^r��~��=�ዒue�B�3>2v�Ux��[v���v[��7���i_s��oc�->1l--�,]�&�~*���T�r��\�G$���2�u޴��+p8pi�P�p�����fNo��=>ǑK�כߔ�E|����R?�ID� �.5���%ْ�c0���w�ܢJ��(�"8�56!+7t#tw}�t�
rm1�$2;�(��ȥ�8��X��Z����-�L�>����7�A�nZ�1��Ɔ�^�Z�aHV9K��<�����6B 5&�Y?��`�?N-��̔+��)&k�,�nų1�(�[f=F�v�ZUcmM⧠'�~��L,sX��wJ����{�[�K+I�qY�ۆI�elN��%]3��ӑn�݈R��A#��ˬbٵ��6z��x��U�IuG�-���V�"���DIg��&&Ǌ= �c#p�@���b�"@K5<Y���{��aQ�g�� �OFZ�Li��,.�nBk���w�H�C5�������궁�M$?�gD��k��?հ����F���>>�;o+t@oL���3`���i���ɤY,�!�G��7 �>�Z�l��W���D��8�)r�H!/�e�A�9��������&�N,�C*�1cAa� [.�ܔ���w�}�>�9D�jnïW�UR#o�����A��\~f/и�[ń�o<�,O9 G�@���&͋�"Ź-l�\�$Ao���PGC3���U҃l}��Ы�u�3%,�����?ls�
����=��f� �nEύ75���ۯ�/�<�l��6�a�;&Ӱ`>9����#8?K��L�ٌ����S$̟+a�Dz��y��������UJ0��`v[Z��!�,�j� �x!�h��P��:��?T`82�6t"�k�Ӻ�^R�+Q,�U���ދ��.B{3��s�B�-N��s��ۛEiV@�?��ݒ��Ǵ�Y�5;�&(�P��'!y)�H-1-�����=�S,TL����ծkZf��T���z��!&�����rX�M��VMC�ҳ���ֆO��3�>�H��j'v^7�ձ�N)/��T��3�\�����v�E��^OK`��L�A��m���Id�f�7l
�3V ;������ �#T�8��`v�/����[�y� ��8�����v��^�.�A��=/Xז��[���O��xT��)�gQ��P���d�^��l��ִǙ nb��$�Û1���j���B���B<��6�tvu��b��j��!�e/��zԥ�Հ�é�ә�6C�u�"M��yq�T�u�#��j)W��bI�,�F�^�S�Őb���C���D�P���y�]f��pn�H�{�힆�'1t��x�!�(B���9�臟[	nV�C��^�G-�AZ�_
��+�0���^��S�P"HL�k(Z�÷;ERz�@��7gt���e����T9��n���@x��d/7>�D���4;�5שH��C�@Aݥ�n��m��H3����I1�\y�ql�aJ�n߳Ś�Z�)�G�B��Y<��y�+&UIzE,h�������K��T�k�ο�� ���C����6��z��(�v�*�?�Cߓj�T>ǯ�g���&�
�)���N��:�)!�Wů�
{�f��w
Z�hn���{Qw�<P�T?�b�%���<=�"���Ӌ�O��3@g���ԃ���,`�^�[�>fxķg��I���oqz �r����_ya�\el�����2�5?;O��U�w̭�e�l��ꄬ�`��P�.DG��ա�1Q|<3<@�'�\�/,�Y1�to\x�e�΃�0�o��uv7�&{�1�<��D�]:�%����aմ[�/Rw�7y&L�}.����f�&�p����_,���%�j�"4�&��M�f�.7��~Wf1����9-ym��Ȯ�3C����q���}�����w[$�.����z6
�!�Ѭj*Yko��k졖�3ǘ��7�t.k۾?Te�I-����/"ßS(?��u��;�S�x\�V��Q�R8��Uî�*�V��t��*\�l��)�*�%�?�����DG=�� �_�6/S�)،�s�JW>�,�;��ۙ���kX�5��D�k����4of���F-o��G�AQ�~�j��|�ȟ��!��*�	0�Y�z@�P���d1R�R����$�`syD��2���`g��6{������lD�5+�y�8���HLW��~G��%�XU,�&�I�,�sOg:�C1�B4���y�P�J@B��߽�%ok��7����Ԓ�S��\��{J�i_x��(��Gva��A��AM�V,�/�G��Zf���	��A�X'�ӮH�S#��Ma��s�ן�4Z%�^(�j@��G��o�X�w�vLLկ��_�;&���T#��������cNu�3~'r��{��h+����Ĥ^�4g`�9�e��}k�V�p��-�П����-��%F&��'Ms�ό�!��V�&iR��Q^�z�y�ד p2�Ra���0�����P��R���Xa(�D�z�S���h��gZk��`H��+�v��w���2Q&��=���)_b���n�[(qDC\|�R�:t�	}�@�R�ᵮ��X��:|,�;~6k52�#��[�k��1����R�� z�֞+����Ȗ�y��/~zDI��XL�����z����+��W .�T�x8�6��k�?�pk3s��2uJ팲�V'n������w��U��=ԖE���nm�i�%�H�#�����`i�;9G5+��C��WWQ�JKtU��^1@�#A)��Q-.�Ț�]�����<u��}��aڄk?Nb5}��kl�"Ƀ�FC��<�m��3	��X�c;�Qեv~B|����m@�5�n�@\}!%s7uT3��%�:0@���ͨ�~��	���Iƈ��vK�V�#���ŃP'�h3�T1����>�r�U��B��w-��J	 ��P����8k�o��w�;���E��aȞ�@=��ec5w���@t!���@�)\�]�w���z��]EѾr^�.Jr0�Kz�-�,P��֝�o]�C���PhKE5�ѽ��&���A�Z��G��ۖ>T�B�y���꣥uC���^V�>hd^�:Cc} p��"ksy��+���Td���";�i�H�cMn��`����f\�u��1�!z�N�'BDM�.�n��V4��iE�g�er�qt�Olz �7�|Y���$A�=�����K�hz>� 8����)}?��~rj�'���Py$j�KL���^뺘���x�&u@�1�?{�;ݯ2�>{��f* ���e�c�H��I��:�H�n�D*�d�-ψk�i�!�k�@&Ad@�xP-���h� xõ�����^gz<z�o)O[u�h��ђ��p��Z��ù�᪗�<�^JK�O����g�p�'�bҺ?*..��ϰ�{��A����%�	Dd�q��儕Cb�f��F)��ʀX��X踴8��B\C�V�\�a��?�A�)ɻ:Z) ����#���l��l��;f�B �ɍ��I�;{�|�7唸� �RS^����V�%��2�[W�"Į�}콷_X)�n�tF���~Q���8�v�O��� ��v�sL���^�*2�uej��1�܍{Ǎ���hg����l+�2Ӏ��K�~�3,F��c5(�5q�JXN11�dC#�zq�ǉ%1�8U��Oj��[уC�d%v�.�U�R^��eD����B�}ؚ���y�Q��Qď�<2�0.�Q��b4��d6/��`w�L@���	]� n۸�ݧG|�nFvcl������S��&|���<��u�V4��� u�7�;���U����n�K��$���t�Tn��4�TP�x0%�_y��5�݈H%B�,˦>�+��w��`�|�E�Ř�(�h�����B�n�_�B�a���5n&��xDહ�h�P]����tه�q�d��{���:��y����5ȼ�[
�rr�p���*�ji�ν���r��[���%�O?���-��e�M{Wh�2����`F�	�Qѳk9�r�p��#9�����u� ��\��Y��\:�P�ﶄ�,E�T�m����G7eTʦy��)r���3y�� ?�뺕TnrJ᎐�`�i���Adz�6v��J��-����U�AH��+�F�#���S�2�߁UX��;7P��N{���G�������|Ҭyں�4�)t����l���ğG�p��
�L��N��)T�	t�/�ϧ�s�㙜����4։A�wݑBA���J:��]��4礙c���J2�f�)"aR'��q����R,��o�Ps�]C����ͧH�:N�֌B���w��yy�M)���p93� ���%w��t��Y���_c">9q��s����X⪇�$)��^�3R4��8����,O��^Pk�Fo%Pu���K}J�w�Z��¸q`BaJ�����3�21�5ք���钟Ꮃy�/���h疈��Y�q��<Y�O�_3{��O���22��6����)<l��"��s��E¿�,y��	�v�Y��\�H7'܇ҵ�m���1��|���2���t&z�KޏR�,c�'�(���ک��Fý���D�8���jb/?ߐ�n�?[�������q�&���BVލ��EqA��tY��8C!��� ,���}�Ig�Ϲժ��k'�F��dw��|%;���dҩ�Z�S�)�m�?J�~�2��T?*�>r��;~��!9����Z'���W�����K���$��+!�f��Qb��ޠ!}����\��+g�2�y�Qb{�֖��OQTrb�#��p�	WJr��B���[~��rDt�#�����w��{Au����O�N��^�ɋ�'0�G�/q{����MOu�J�<~z�Yg�MG�+�C$}�2���H��ѡ;k��gp��W�+�ï�������W+Y$�[&�7�3]�߭]l��5�j�J��{ͦf
����#?kc|�r��~�z�@}�kCU������(��L����� �#�����4��9V^�@�|�����qD˴�f9�c4�l�A���kӽB�E ��/�/�Q0D���'����z������׿`8:�,��C�c����ɓD���I�0Vj1+�}�	,��ڙ�z9c� T���/��c��[��!_�>u�?��R�Z��i��ՄX��d��$��c+��v����'+�ܷ��D��oJA��(�@��U��%�w��c��������UsC����檒X]�}m�!m��'/�,/?$��x0��a\�����F:Yeo��~��X�����R��ꦣ���z@�]M=w��aԻӫ�>j��:��c�0"�`�RA�V=�s� Y��l�r/�A�)��q���l. ��ufQe�YgG��_���8�B]n���6=�5�9S��}�]��k�W��)\9��a}��gA)"Q��ȹ^�O��\��뵯��\��C�h0�:r6}�;�i��o�@�A&�s����O�p�d%�)��#s�C:�}AB[���\���#�F6y���nG��kۻ������C��	"o>�Tl��x��!y�nL��QSg;/c�s%L'�U�������d%'^��LkN�l���Q"�W#�4W
^.�|�C-5�I��N���:���q�N�j}@��<�� g��������4�N}�"a��^�#�l���Wjl����T�u�v�5�|Lh���S�j?��98qBB��n����T��6�������gn�a�|�ќ�&l�7?0���h�/Y ��:[.��rq�s�S�	�ޖ^%�څ���kqv�Y���Q Wy?:.��Q΃�
(yt~Vs��<��.4����HՆ��s�{��\�C�-},��Bæ�2����M_�%�����P����OM��8�&m�����x�1J���TI������;ݤ!ù�p�ĽW{tr���޿
A�*!��j͚g��=���dj�G���`�x�iX
7��6o���%��+�6#^�|k%�ʳ���ï_�)	Ԡ���R�"+x�z<h���{�&t��X�.Xqہ�H0��-�'O}���uy|�����0�ͥ諕��=Z���2�/�~L�6&�g |�h_TK'$�_R�%$Ƥc�AE��?4L$�/�%�G�:��]��d�_h�;}�Ĥz��tK
����#ՂN�"�)�����X�U5�jز�D6�6�P�)jJ6r���Bp0]@8�teu���cK����4����m��g�?��T�!�l3}���erje=��\�u}洝�@�-\Y�]�1TjYPilՏ��c��]�bcU��{���ꌞvk5�Z�)�,� �0���̫���HA�ܽ������;�5��@ݦ>[���A�N p[�5Sb�;��<���n��k�T��	����U�ƛ��Y���+��i����O��ϼ9��;�6��3y:[\Y���L���6bm$�]�]��H��4��;���w��M=!13nJ%�5ծ��q-��6�ݳ���^3����0����Jzp7�EM;����e3�\�_=���.�XR(cK�şIE-�����K���s���:h�1`�i2� �3�2T��ufs��'r����a����ů�-m��я=������'U�W�v9L��bރ�aU\�����<Șx�RFO�\Vn�9*U'�D߿�53/�t��Oj�Z���H *�L� 'J�w={�g����Rg��%��&�%����F�����?P̄�j�{ǳ͕#\ lr�l<,�A���0̟ML����QQ�h���)��,�}� ��M��<�r��U8R����z�ԏ��ǐU�+�uDF$��
Q�{�& �]Wt��(z�N�+��`����F�6�XA���jX��_��u�*���BHD 4H
���Xh�fY'|y��Ɂ6wC���e�D�t�
��t<r�s��ݧ�[n��-��ln�-����0[�d� ğcS����s�e���X�$��*��C!�uUqR���LMU bd鉿�vwθJ���]o�䭹�M��2ʣ�p~��r+�veJ������M� �Й[.XZ��XO���\�ќExz�)-1䗵	�O&Y"�U��H|l *z�+:0�j^\X���-�o���T�.B�y�L��fI�kCJ��8��POt8�fx%��\��7W������+�]׬	x�ՌSJ'���o�/���O%�|Q�"=?�۷��G_��S�>�o�[�h{��X��d%r����W��6��M��<���r�n�[�������Ε�>*྇�͉�f�5Z�+i~�3^� k��>�$�9!�*���A����!0�"n�䧼�>�GRa=�;�J����5��'&�������~owy�Ґ�j���C;�P���ψ�iNEn��el_^��Z��q���>�؂+b��D��<��!h�f��Ba�����z�s��}�S�²�]w6���<���\�pk�N-���g]���os�x��c%J
�ܫs�f��/9uo�����Rq��h��Ӑ����{�6�o�#�}��&��s4y�+�����%�>���e��R�Z?h�� 5�!	.�ei5,X�	��c{���?��+xG<3抖>�"2��X-�y��x8�����_Pz�ֳe��;��R���?-��䪝+&��R��l�5Q���$k
U�J��_��И���F3��(��Z���f�5�9�Q�7���6J�W���o�'�>W�ƅQ�ꆲ:����iU���@�X?Ln��5_M�E�.Z,6�~��<2р��oH�Lex�d,t�I)�b�f���c�E�e��̊(b�&���?���O����o ��<��?��!��F������AW��8�ݱX�CCkVQ��)��;�e���?�ԲeP���䅇fu{ځ�g`��\�F �r������-Pc���j7��V��+��zQ��fkaպ���_J��)��$w}�8{��Ge��΋�?�Z����fb�䶤"����:�ǎ��+)]*�-���"��B��ɼ��W�[u3�X]g�O�u9�_��6�5z1�(����x^~�%tJ�z#m�Ь6��;��n�G�r��\�1A/��W��b;m�R��u�$ZH"��Ś�u���j�l��+��Ʋ{�Ӆ�t	|��f����B�2�
���c�#�J���-�v~��ަ�/Y#	w���΃������-�*m2���=��e�	5��ç������L��q��*Sɪ0�vV��|��so��m��\�Df�,V�W=v�+�ͬ?��i����Aս��-u�=P��u�7x�N�2 ��joݽ�P%���q����U��M0Hr����Nۃ��(Qƽxe�������ɮ:�ъ�dT^�#ɔ7��6}g�L�_f\���6v��I�vpT��`��6�r�Q�4�?L�=���9p���1B�������ۤ��q7�d��X?�j��	��x���_��T) �'Ȃ�S=�����`��@����i�T��)�K�,�r���FVd�b����4����9��~�6�Ɗ��(%V��͎�	����Ȯk�E赺S��Uձܞ��O�x���b#�9���-|�C{,���Cv�N�d��j�F��n@��'|>;fߋ�G/�1�v�ד��s�g���ֹ�_~ �.��r�A�l.ͧ�zͥ�(}��ܙ��YQ��6�x��@�Q�.�|&��*��0S4���.~}O�hz����΋*:"P��G(��E'�Kܓm������W���n�I�� N�?Z���4AL��>��1�ڸ�(,n���P�
��qo0F�����I��'<h@OV|^�4c%�%&����Q7�jn������2����ɐ�-�6�n��map�g�Oa�і�A^hnB��ขZ� R��IW:q�&�I�Q�����V�t�V|k0�sb6K��th�h�m���N�� Ko���uH (�ny��Ps�\���� ��S'�5K�����}���A �R���6��ɔ�:�� \⃬R��]>ҎR��q�k�Ý��@2�1.��������'��[QK<�|hc�L}>��v��@���b�+�MB=ۤ��$���2���{e�E�o2������]n�f���o�B���颀�V�y�q�Ֆ��3BiU���;n���*mI�'@�>A��exO��Ϧ���/ ߂j��␱�<���"��r b_�> B��v!hքs���'���&D�R��/�
�HР��e҉��s%�+u�y�o�0�!^�Ne�U<8W��D�&�QD����1�Ge��̮5���ޟ���e/��ORc2B����f�n���Gh[X��+�_uS�����ؔFP���S2Q&�R�����|(]��p��de���I�k��{���נ�)d͜���!��w~�)�`a]�;jC�;�w-S>��s`����'n�#�w��]|Qr@n�,����9mr�t���i��}ȓZ^�/w���U"�A��#��Ǔ!L�#��1Ra��g`�ϻ�x��u��N�pr$����e;Y�>��D�y�Q;�s���	�_>����W�H^,��������~K��(�$5*�H���R�|��&������\}�u ��t�-�B�y���@"�j�\�~����F�'���A|�!�䝰����ڂ̷� �D�
J�R��005�Ļq��ߖ�V��#�3��>v-;���.�U�����W�&Y�g�����W���C�LrY�z��9�Y���U��Z��5��_\��މ��4-k��JDQ��y�Fjس�����Y�o���I�ഁ���؃ًA�c�m1S�����V�ȉ�G�e'�':q���$��UT�<��~�6��D|�w1�-�9�F����8Fm�d2~tDZC�߇!�Ж"[�����\�B��/��5I$	K�a0�H.R���D�*U'���ʋ&NB�Դt�S#=^�}E�]��;�/�ї�H�����P�Bπ.1��U3��J�1��z��PTN�K�w��kQì��#��������k�9bƢ��"�"[���[X�%��� �����v_f�cȗv�k�=7*jՂ5*KF�zbAm�#Ᏸ6�������Aƀ�y�㤡�+Y~��X��1�3��k�$p��S�/B���{���jO���`0ύ)?�^0%�r�D��te��ɤj��bYyĦ$�t.��s����W[�1��h7q}ү�h�	�e$!%b��ژ��0G`��#�*��m%E4aݿ��Y۾=H79psc ���E%t��k��͊��4C�rt�>�d��5'ڵ4�X�Yu�x�x,�>����Ϥ��t�*��h*x��k���9�a�9v��ʄ@`�<L���V(�=ѩ|�G���`�Bo<1�l�r�N2��)��1��5lyߍ5!�n4�6-�w_�~�5�b�F��*��t�5��JB�Y>�Tr�'�*�a
�H��(��:c�;�g:�Ѓ��1��~�d�(�;"T�	��������p��>y��Dx�X��ڞ����X~�"�å
P�d ��V����pEE��,�y����$���ف�՝�/JL�.A�)���������x}����;�w�)�(eֹ� #0k�@�xW�Fqy�?=���g�=-)/W,@�������{����s�Mּ� ��*"Hj�uo1�[+�A�6�O�@Q{L���� ��#� ��Q�&]Wf��Q�2(��re��$��  A��D�Y�U��>��ˠ6RG���P�ҽ9wLu�����w��������ɮ4����ʒЧ1B��L�2�T�Nv�f��j�4-B8j�-�/�9��@�0�����y��=sSՈ2$�>���6;#_�R�6%T�<{�����n�����S��h][>C��3��Ti��hI�@������;¸h��_�i ��y�@�&^� ��++�U|݊t�]�Nw>9��2_ۆ��x�E��[�����9"�%�$�o���e��������1ժ�4כEc	W�����)�� /<�!��{������,�^*h�S��U��{�Θ�]t�v;�wA�_7Z1J�4����<�J~�^�zQ�uxd��20p��p�N���A�j�ܶE��?0[�I�r3���u?�������G)5�6�9d^�W�B?���3��~���"�ǻ[a��qD"g7Q��3�?%��������$J)R�%�`۠&328%����g�5w�,���2;k�ecJѴ�2�n���J0N_X����F�Ugy�g�^r"�e�}M�En}g��1����g�M���,��ȭ����6m�����`>  i�绱�|�E%・�:����&Ng2���(���
hjib��
-������K#V�y��~uߑt���&���#��|H�^C�"[o2�}�r�x���#k�	k�R��m�5�����A	�
RS��7f�=X%,;ظ�� X�;{�/�2!��n�$x4��)� +���ݶ����~^PV�[�m���D����8�
�X�"_C�'0��Ɨ+�.����9~�Z�k&9^z�����#�嫜a#�l�73�8�<3��&Lni�N�;�@W(�t������̳D�e�u��q�����aK(�ѣ�$0��� �\=��:�C%\homf2;���Ih�El�r `!�oW�i�'�Fe�� ӮUv��>��;;���"s�$��y#��	 ���K��l�t�/x݇��d��qd��H1Q�&o�He��L�(Sm.���,~���w�[�q�/�x$��ͳ�+A���O��)��	�kǽYS����d��r���<-}�,Lj䄑A�.ͩuHd���Ԍ�S�
j�cr��{-�J����$i�e*���|6��uAU8�(�� 鬵*�H2�}2��p�[�Y�X�Og9�0�@ tk���5+���R��s����?I�3Is.�!@����Y�X=��4��ʠ.�qsގ����p��%*��/ď>��������J=�����T2��۾%U�����g9|3�L�B���ս��������*��P��U�=�J�Emd�[�?;��1�.�ꗨתM,D���Zq׺SjU��e6��\�0Ef 땪ì�\��eH��)c�B�)��E�� �0�HW����Ae�c�%�,��w1|���@�Qʣƺ(�z���r���%����Z�hQ<ǒ#4�~�$[a�"�&=Կ4z�O�/����v`O�^R42�q�n���Wb,�`�"�����ՙ�=�0i�Vp�7��E�O;���;���Ɲ�܌����u�������E�FT�Z��U�u<?��bJT��z�{����T7網Y���][ն�#��q���`��,�nuXi�Vq�ʹ	Љ@ڣ&��5�D�\����`�Y�}�1�����z�{���'��~w$��Zz1����gO�����)�߳wR����U���iԘ��"��Eq�2���V0���r Љ!Rʋ���!̊Z�_�g�!�'�	�'�gx�j��������39�@JF��
>0֬ʔ��Qd_���%=TPp,g%��{GT��	�BEՒY|�q����b���\���������H�++�X	�Z���Gw�i��굜i1���Ku�[�譲�1�V���\sBxEEw��afD�RT�`�[[�<O�9ycj.
���K�8�ncrP�B �,�����\��2_�H�o���,  �d �/����1pP�Cø�Mvu:��!%.�B��n#}/�_ٗ�t�lq/�+�����F�΢^"ڳ��>�WG�l����<C�<~?6�ao&[N�C�*a����B,�K�ჱ���w����ʦf��߇��R��*נ��s3�C�*����P����ҨP�����f�(�
���c�L��+ȍ����,*E��}��ƙ�01�����0��V�'M;^0+0���s��)9HQp��W�H��!�y�q��Q�*�"%���^+�=�i|�>+�?��4�C�:�n������T}��H'��5L��������];��[NP��Ap{.�9�ɛ� �tK�1nG	�������u���3(���e�>lv��Y�����K���P�Y9���:�����
�I=�����A`����0��&w�$j9�Ý�
G՝�-|B���B�5��Za���ܩ���|��9�M��X���^�+�ɻ�Ǖ�����0��t�n2@6LX�����@s9����CV�4j0H#�l�!P��TMn�M�	�0r��[��9׮d�7w�<X�]�j���Q/�|�ۉ��6ׁv�����L������I�&����F�RB���ws&L!Ds�RȓלOu�������am�f (�";@�e���1��3��<�h�ׂe��G۬g��>'���Fon�@��U�;�aI�fgc����-�* �Kx �'�댶Ь�A/��%�}�q8�6�]o�5Z�X/�g���YE�n3��xuL����!�����I!E2?����-�^�����w���B�s����I�I�nY%�#�)|�Ώ�J���dlR9���{�҄�%p����ݫ j�j�І����K�hHah[��01`n�q�sΐg��wsHAa�D�����Z63�`ޓ`E��U���_G��e���kR����fa�ZxW����Y_��G{�g��j_6�$`�n{��x�B듡#��2��	�����H����C*jky ��]O|~��!�j�8�DR�y�����%����TdGI�ĩe�l�o��k}~�g]��9bn+�Xz~��q�N��n��b�9$4mwοC:)��\�4������ΧSgɨ�o�&��nۯ���ԉ�s�P��q~o��O"θ����%��ܥI��I�uRz��.�z5�"�1��aP��W�^�R��~6����%5�ݷ8{��ߵՀ�����iX�	z���>Ҋ����>a��H�[]j����e��y6�G�J�%���^2h`�5a�����%km�
�T�:� j}dE<R��^h�}ap������ې(�����`� �'E��J�ՙ`�����./��� ����y�$����y�B���q��n�L3�C�N�S��zBkYY��a�'+������J7�������J��.-�,�ϴ�5(���rX���7?�xմ?��)x�g�^k�Gs�+PS|%sQ��ѽ�ޭ�3ӗ����&��4�C	 ���xҬ�я�S�0��x�C����_�����]��r���x���T���J*�i�i�?��T`1l]u�#�Q�oX��j.�:�3]�87CO�)��{�>[`���?'�Mc2���x=�z����t�0�ZcS]�Q��mK����֖d���ݍ��Ka��|��|�ɢu����vo�P�X��O���gǌ�\9&q�k_�,���d�}��X{$�c��B�5�����D��c�ܔ���Hû֙� �ݜd��XAA��.�P�%4�����+D.*�_�lo[��*�/�)���l�e6	�8})�a��o��YLG����d�:]P�-�ܨ�����e�?c�an�����e=1Ԭ�C�It�'�>���l���{�;�I7(��a.��$<��;jݭ]Y(��<�^K$ay����'e�����8ץ�v���;�����ZC!?�걭�Nl/�s/O��y�$�Dk���c71E6��t��Y�ܹSɮHIۇe�y�<���[8*g�*�O��%2;QO��wd�%�Y�MBXj:;�wp��V�yr�(�y�)�Aq�E���8��5j���1Ƿp8���!�dZ���'7��_(C����"�D~��h����kӘ���(�g���zؚ�h4�t|{\&K����$������o��� ��6`�ͼ�:r��_nk�� �Xf�2K���k�@�.��k?��M���Z4��N�؈PU����t�}�3�z4�8���N�?���AN�ɶ��F�gXa�dD�;���&��I�BUF���<����M�$�#>�mM���یrp<d�w�s�V�����IEg%AN��8�>}��T��*&g��ER�.�@���Ij�\��֑'Dzm����_�%���p�٨īRd�jC�_OB�;�6�~��_��A��/�j:M�\��0=W�!�oLv�w�(�	�Y�B!&=`�K���kwh�3(��Om����[���%Hud�`�Ό�3����͚"*h(u�}o��d�������[�s�R���Yj
�ӄ��\O��1+�[ �jݨ���o'�5���Y��thB[�C�U�ѷ��~+v>Kp �a&���-�gl�8����.G��ݕ��ld�&����&I��8�:�ֻ�9�^��@�XwQ����T�@��y+M��~l)��>	\�;��Z~�Á$]]�E�ݹې��e���g����4M�oF��j7���A��
�l�*��v�z5L *o��˔
Rq`�,1/if:��w��zQ�y|�I$�ɴF�����/w4�Q��Fá�-��0�|n����x� /,J},�y+���is����+�ۖ��q\u��jT>hC\~���`��7PA}l�x�I�'��
ZӖ]cx��urVs'e��0Β-Z�m���$"�Sۇm�O�;rd���w��W)�$2M@�a��u���0���Г�t&�M�_-�&I3�3epY�ˈ��Q#�醴y�Q��l�X˫�Qf�P�Z<�xB�J�`$�O!���H!��rH}��@�>}z::6��g�<���[�i��/�=���3��O�[���&��v=�ߡd���8M�����i�>�lg�|�ָjW ��+g��DgD��ׂ��?DQ�����j+�Q�P!��o;��׀dA�D}�l�]IC��=u��]��>��XW�^E,����7;W�������m��7z��G���[��U�I�F����� &'`����[�b�4�h|t����o�PFO���|�Y[��׊��7Ye�œ�|D�����0��� 3u�_��D��*�>��0��h�����D��X���m)@�i����T3�h��-G����5�0p� �i<Mɲ����}H��-�_O�
^��z2֚^����Rf�i�B���]��=���9�o{g8����|E����s7���]7����aF���^��Aց��T[��[��_.z��i��3cBVa)����o��Ř"#�8�����a�Gj((��~���)�%ύ�AU���LAZ:C�p.�l*�{v�;�W��pKE~퇍�Ȼ��<�T�_��3/uꔈ�OV�D��$��8��=t)�6y�mP(�e�cЫq1�^��nZ��8\��ʲn=fo#����#K�1B�ᚏ��:��N��&�̈́�Q�UE,*�L�������IA%��ĺ�<��*�쾐����p.���j�18�F?%d����d�Z� �vW�V^@ 5<���3J=��h��Ur����[��a6Y�c���F���X��"���S2�V�ΝrE<�_�[�b���$���NґQ�.�Q�^"�o.3��>J�p�V��cTU�ۇ��5Z�	)ƨӴj*�l�S@���0���2�뀥n�2o~i���s�|�'H���X�a��Opx��dfL�i���Z�W��/�q��9qr��%:>��}���
�m��1!���Ƣ�m�ޙ���.C�6�Zb��:S"�2�D�T��:�clS6=%���gn�`}�pxH(��c���)�~���l���d�3�cV�"Q�~Ԕ��Uʿx��Z�4Ί�3��K:@��C:�7���ߒ���?t%���0����^���.5���ꢿ��;.Z�İ`�_��m���!qJ8Դ��	�/~��%Bz��$��T��,�ƺ��ϼ����aa��{X�U��?����Ψ�\Q��W8��:�(%^��ܤ����x�7������<�*ΰ�����=�"JP�w[�Ӌ����(n)���W���j2@B�ȶ=
���}�/@���*a�ݽg�w�bY��*�R�Z���xܣ���U������t�g{�s�	���5i�F�%��Q��.Mx�b��Er׳7����� �w�q����"�Bk��>����l��*4(��ۄ��x�0m�c�VRk���3�fk]Xf�y" h��mZx���H���<Tn��p��?����)����^�3V_Ӝ�H�=[�"J��#�n%�/��u���E�٘�������3B*�Y�5t}.�ip1l�|�_�i�t�����W�Z�V>1?�����JO���\��H�V�����8X��l�$-�{���Gco�"�"�v��؜j�G��R��E/����$�l�Ə�Tr��ʡ6��K[�@ߧi��o�S�K� E3�z^s*4c���6�%�������w�rsYU6��̭d	���f��qvj�bJ��_ɕ~�mR���<��}�)@]A�uk����A3Vy�&�n������^21���)U
%R��{�4?A�kƸ���@�w�`!_�T��s�>.����=�ʒ�lG������d�����8�y�7z|�V�ЭD��G_)�W�p����f�dUܬ&iU�I
�;�wl@���|<�n�|��KQ���/'�s��޿kK;ӱ�L2X�Za��d³���s�3�W}��W\����Xߧ��غ���RBY�1MC�(�q����vV��I8�'�t�9g�̫Fb���(� ���a/_O$�M\8�D$�L��Y
�4�g�N��J��B�����x�o��ץ)�w����is�vG���XD�KAN/F����n�T���B�=�{�P5"ﾮU�R��!uL��¦���)KN�N�60�e��üKE���C��^��U�8 �ҡM�8/��.���&�X�;�����P�A ��氱����n츰�j���rS�Ah���S���.�߁��x��f�fOz�!�P�vk�t�[y@7��S{;(��J�������&�����ܜs�e^a�� !����,6؝�,k���}��U�H͸bB�;�����`Vh�I|���5.Cn��Z*��m�+�[,v�R�"����}��3���'zC�ys�����8�ME'mEdz��paݘ>��/m�����&dϾ���6M���o�=�sC�;�#�>b5rk�i>P�
�e�|�����)�dp��]���B��� �k�!v�} ��\-�DA�����ԡ:55)��\�}x��¸ך��@�m~C>��n�q���˾b��-���xKWug�%���X�y@Z%.��Ă�!�s�8��TB��0ců쁮���\��^�m�N�@����QH�dK���zBLZ8QW�3�ͪ��Q.w���;=�iV���֙7�b���V�����Spr!`~��D�ڭ�-���|HV�v��Ea��֠��iB�Q�D��Ճ��s?#bi[�g	I�1�{w�&��ghwx�)���6>xW���w���`�O˕���M���B��ΦZ[^K!��`J����E���{�9c�ޡ�ƊZ�;��`��_�?X|�a���]� XM8�����۩�*�eB�w�f�F�ʚb�̸"��n��A������e�!�ft���~Q1_�1�^܂nYhL'<��>H�"��
X��1�ٙHHo��G�֜������ų�L�*�����`�޳����EwJRbv|NC���0�-����K�s�v�����o�'}��V[:\_�@��	?5��d�բl!�`(5�7	�ꃸ�lH����ͳ������|���^�&��>nNTuVgv �]�n�rP�(N��ɗ�du�K�j��2	x�2Q.��k~
b0�TS6D;�^�=��o	�� %Ʒ'�q ��Ɍ��:���.�Ř�`@涍H~�.���.�\�9�Zt&��* W$m���Ơt���7�4�x4Ke�z�ވ�kka�ZPA�K�e���F^�DK�_������-�!�lx?�j�)��ݭ�2��M�	l3��4L�ͳM9&{1Z޴Op����63_D!�:���M��_�9lLn���MZO='l�����(�0Jl������!UTƒ|�KE���6�����"*�2���7 353Pb��ҡ�#��������Ua���0�Ȑ�˷k�+8��;�s;v���cQ�/����������VB5$p�AWsb~=Jo!9_��k&��bSk]�����C����'�R�wq
52�"�>���q n��!�f)/bsҥa�gֹc���.�KR|F��ix��f���$�����]-9�x �vW}�M����h�O�u�v��>��f2�h���o�y��i�ɖ1g�e'�uL	TkN����ū�����M���a]4�u"�v��˦���wH|Y�֟r�/I
�4�w�&�)�#y�T�۞(��<L�{Y#����C����۰�SixE3�?cp��<	�� �R�zyV��,T�!���WQ�t�c�\ \T�GGZ�7�!:�Ks��^�d���G`����'�~��
��[���k[��p�J�����K���s��>Y�'a� ��h����1���F5��gy�2��`�R"Y"�8�E�x���Ӹ�y�Y4����[�B�ZJ^�<�\�z/�FFoSx20��PJ��۰�v{5�7���ܽV�����c�����M���9�`����֜C�d9[f� R+�rK�T���p�c@w��1��O#$�ϳn�o�Sοl�[�^��;�K���kA���"0��P�rz�J[3l����Tø�C}{+��lZ�?�A=���~��g3�������IwG⠬h�)K �i3�j���yV-s|)�++R>VZ�o�b�5�0_�'�@���[Eȳȱ)����� ���k�myؘv��E|}��GX��4כϠ��pL#���Y��t,�b��3@?Rf@
E��Ǎk��[G����y�!�D�� t.ߜh��B�9��p^W�T�x���Z�_X�2�h���V8(s�d�j	^RyH	���+N�X���R�X�P�0c�i���p�Ģ�~Yn(a�>��9ڋ��+Q#gW��c㛶����&�	���#D�`p:`Dx �����.0��\�sp�_��vH_�ø��b�&�F��W/��3v��P�a_�@��-Q����������U!�����]tF
b��=�%9!�Q�Q;�\�Ӓ�8��}��b�O�Una56���]4��e76$�b`P�Z���ѝ���5��]Q��Q�Ý���<�w�,-�m��NȶyU���ج��M	Y����l�s,���ޗ��	� ��L���q
�Bn��_0V��,A���R�*:i��ۭ@�W���5�ɛr��1n���"B�u�X�1"�$��sn�Z�T<��	��[K_xLbX��E�Gz��rB�}�T�]	mU���cN�଀�b����$��(Q�W=��r��ݮS=6�y#�\1���z���Yh�(A��?�Q��Q�N٫�տ ��J�MR�)ӿ��*^�\�~�@?؞	����*:�TX����]B����n�r������Yً+H�V#ҟ��E�y��u��H�fȿ6_¨�FY�f!�J�)->�ҚP+V6���J��iyrQ?�~����򥽠u{��Ǌc�;�AU��y�i����U �Q�0J��(�P�*�Q)�W�sr�3=�U%�Y�k����O�Dt�ձt�ڨ�����)�)N�i��0���%`R�)�d�PtM�"";pM�h=���Z�=�r}����?u�m��)�I����mJ�f3�z�>��k����f��;�m����#Փ4!�v�o�I������Ӝ�<�}R���cb]p��F-���2iL�v&���~�?I���3��y��@���M@bII�����9�� ��=u#P���
�1�
د.�3 Bza.�p�1����M,MU�j��P^u�����ʴ'���� X�`�:�Z4��1'Ny�:�maY�K�	�^F��C�����dJ+4"K��c^	�6���9�!�D�R��]/֣y8/3�ڻݓP_��Jtc�]�\�93[�j�*"�R~/<��������'����=��3bM�
 ;J��כ`_�@r�Z�U�m�8y�m4��զ���V8�s.�P�n9�:�W=c$cL�i�4����<�y�%��FW*���!H��ⓄKJ��?v��[y���\׻��<>^���8�ڏL�f�Du��<ґ9����z����J����L�� ��ԃ���j�Ad��~��6�7˒��Э�ZQaPm@5?�5 ���>��e������HSB�4r $"R�u1�N�36�cK!�O�����{Yi�r6�zq�"\�Eg�&��1Y
_ԀWJ�`;���̪<��������yaZ�C�N5�9L���c���)T��E:>��9%���+�6�A��%M��[;x�����,3m�s�{�Mѝ��BM+��Yen�]�b�����v��0v�������� ��������2���`/��� ��pGb7g���lQ8�j��[D;`Z~
��@j:-� ��`	#����>l󸠖^�~W�]}{�m�]ه/ީ@C�-2o�W�l*ĥ�^��t�K �ǆ~]ܯ�H&�֒�TC*���	�ґ\�w�/ܺ��p�J#���z�M�${i�����UC| ��Լ<d����4�����iښmP"w$@���C�ٳW2T<�#8#L��:Ѓ!3���[�)p��]�[�Ϋ�|�8_��r�����1m�3h�M)��h���a��f��x�ƥG0ֱ�D�)�:�뺚j}i�����W��X��Xձ��DW��8QA�:���ߓ�/P�dIɕS�iV�>�J�Ip�J�dUt��.��W?��1��C�!mz�V��HRW�G6u�)*�8��AP�	�����?f���@�k�6Hk�6�l��Ph��Oxٛ��,{Fɨ?��Ӌb���S�?�`�g�l�����=]�"'�
���:\�������e���O�ݥ��������q�b@F<j.e�dhH�!��p�dk9�C����d�{�fT��T�gcX�+nñ�$�/�=�*� 8�O-�^���iC�&�C� B�9�7
�rp�3s$>�l��9?� ]�B��|��2{���U�ݾ����<�-�;B;Uk�h����q�<0��&��&
��d< �����n 1@�]@)�44A�$��{hԃ"��8i�@}�'ғ6>=,MN�B��a�_e��L{硵�3�|����{�D���T���i�%
���66nU�8E�<ȁJ����@��:�A��EVG�d^c�E:�f��R����6�j�BT���8���[�[��ꑉ���������@qe�]��r�=���ACUL���Q'v'�N�N�\4�Y:,�]��$4qd)	OR����iw�J������1��6�i���T��y/*�t�=Skg��|~�� �!����L#�;�S��\n.�I4@D��w��~>��{L�{�K4��X�
���{�i����,2e�#���m+��n��!DS9��:m�������^
����巍;�v0*�2%u��Y>r�t�	:,ݗE�ʂD{Ƭ���#�c�M��t[
�l�j��� �Pn���X��!י�,���>D��  6p�E<�s�=���0��M��^QRd�Z�i�䨴h�)�����K�*�7���J�X@�m\��y�4���.4�1���0�B)���F-X��9CTG�o���Z��㿇v!/9ꖾf

֠�=�Q�߶��٧�d����[T�b�-4��ϗO���+���Ql��^ @R�
��DoXȆ/�����r'�p6�����kM9��]�b=� �8�P~�k��2������G��* 5��tO]�]������Q���Ѯ@T��Bj���a�d���b��䌵�D�]����F���J�>�(�A��rP�2ӫ��Ɂ6$'	tL�H리^���F N���(���p�`�	�����{��I"�Ւ�d�"�Z-�dj��dUM#CΎnwn�C}���ہ�J�� ����·�E�����>�k�ͯѿ���>N�p�P��7�C�*�S�.gm����;	���L;��΂&U��{�2Y�ũ-64,!��0�9� ѷ��>�1 {��ݐX���U˾��g.��ͱ�_��%	t�h��x!����$$��C�.}�TeA�ˌѱ�/�����G�O���6MGZS�������
i#��;�qZ�L�K��4�,>я�C�9�b�nب_��c0̘��0�Q�L�yt���?��l;�n�c��0[E���g�}��~��:Q�����F�Gc#�����DXiO�5�y�J�^|�)�cG�V��]����>��2 �0�~�Y� `m��^K�sM�C�x�8�c�����mWq�a�G P�"h�����.8�I�g��>fX�g�����QI҄�$U�V+.'g.D����DL1�TɐB|����~[Y���`x|���_�Wk���+R-��m>S�J�e*o������-~�M�Q� ~[R�D�o���� ah��d����8�c>eP�-��m#aD�#����j�I��X&�&;��_>�8���Yl��C�.� �ߵ����L�Y��#����9�"ة���|��)B��|o��#Q˒(3�@ JXK���r����?���ؾ��������2i��� �����'Av1R	I��Mo'��z���|x� ��wHn�$r�O���m�����'ċ�y���c��A�2�,��,/���7^e���i*������*15��@E��Y�:��آ>AeSS5�d���9�s�3����j�;�'�)'�V�sAj� ��Fj�^�y�_�lQÂ��{Ȃ�:�P��*.��X$ǝt5a�1�B����G	���[�������Ili�Ⱥ��6ޝ�:��� �vnL6]�]�Y��jÏRGi&�D+�����K}��oJ�������h���Z�����~��3�A�1��8*���//Gw����tG�P`%r�ZH�>�Ʒ��U�z�;��D|"��Z��F7/	�,�>CR���ƫH�s�Q�I��ZQ|��,2rM{Vu8��4x�'�y5�+k���كg��V76�1kpND{�: :4+������BL�%v�!�1~o|�J$N�k�Vd�P�a���0��e�t	�����<{T�#�~��5�\r�t6޽JC�,� �x����^F�u����Ҝ��(z��/�B;q������gu�շd� ��U�M��_�F��_�_��\�a\�ٱ���/�i1�^^7��4]#�J+��|�-�<QQe-����N�hsp9��V��Q@V�Gʵ5Jŷ�H�>�+�����G�:�6�Pr�>^��%���5����M�&�qQ<Y��� �dV �S!�<}3�?�Iڈ\������g4֤�J� ��4b#�:�rc�D�7Ӷ�f�"E"�������Pְ*Kyhx�5l��n-���#��%O��Q^����VM��:�Y;ʫ���$�'�^��.�}��gwP��2��.����Ea*U	�6�^�ߙW��䘧o��[!\�S�0;�I�nz�=H�t�g��}9 leB����%�Y�@��>�Ngd|2�g�����%���r�6���q}M�$âINV�h�)�1W��"x�!��-�$v����_ܨ�Q�9y�"!�4G2�l��35#�kj|�؁w�����y[E�6�k�-_��_~a$��2��K�z*�t/S ^q�D����WS�"�H0�@�����l�fx�&�	�G��[_�b��B>��UX�4��z=�X�DhBP�'й*@��T}5嵀�L�/R����9�#��7k��X���j����kj�=��WE��\OGT�.��M�� �ɾ@,v�!��z���dPl�O��o�]+��Э�5zO��
|5��t1� =jq�Կ�D�Ӥ����6�I��_�va���C�d��.�~T�~��~�9G��t�pf� ��%�DZ�G��(����q�T����'��H�;��:�P�dQl�M7Ķ���Q3L2�q+e%�+��SG5��7�@	�L�@���P-vnq�mZ������7&�6XK�� %hdq��y~0���c
Q��&�Mf�K%X)�2��?����@'�c9/��<�J?�$Aڰ~��9��Bޘߠ��!��,�1}��=�e����J�����D�Vx=~'�s[y��kH�g"��/�	����G����1����)S��֘�=֙&�Gv���l���6��SqC���h,b��H �Cu��礆9��w��}�ǤB��oz�s�ג�	�pzd��
}w5��OK��M�$�.������Fp��V�w�*eŤz/*DʌqR�*���u�<�,��m-�G�r<�q>",�}��c�D�}{0Q�,d-	R�.�󙥡Q��"Ւ~U�昵��+AM��Cd��;�ȡ�E��\ �_�$L�$�'�n. ��c�`X9O�`'l�T<)�Fq�#A&�~:.)�6���Te�GN�09�	�[�^7���9@��%��7�Ӹ�Hŀ��2/ĒZ�y�{@�$���f˗lcܞQ!�T�h����M���%q� ep#I��K�[nO�wn����~V*+���E�!#u�|io�C+}2:���ꃣN��
lj��Z�س�p�~s�����y���=d�D�NjKk��$Y�&��*?��>��2:�=�R�^��T�w�[������|(N��Y�x��V7fȣ���M�S�xc�(����΋'#w��O��^aX�x��j����Et4"8df�������Q���m4��( �}=�5' �!���|=y����\���["!l�re��#ݾ�� �P�m��hE�"i���e���i�a�sl���j�.�=$P�?�Lm�d��H
���<׿S�ڳ�Uhj�ۛa؅��c@s~WJ�uE����i)Z�������u�F�]y�7�"9ҩ�å>�^����bV��"�5�]Dk�/)!�]/d��e~ҿ��0Zᷞ~������ù��]w�6�:���0\,� ����^:m�q^_1���5
� &�&j�?H�.�4N*�>�����k��7��r�E��� �jʭ�#rg�9t8�R��N��f[E�/�\�H�`5�o����
e{ �(�З7���@f�Hb7���-�p��	�7oq��u�f�<�[(��恿���ԑDvӸ���p�Ao:�d�1�o�L���Y��
�,3�]�Y�-�)�i��T� X4����ȳ���B���΄��}����(����vɑ\�j��B���n�Y��]����,�_�;��6��E�%3S�;�S3?�Si�AR��D�1�Z?u�+�Ÿ M]���Y;H�Lk�S�vvI��|����9\�v���>ւ�"��EE?��^t��\0 ~';������
XWLG��4�� ��JO��'���_�Z-%����3irpi�>��AY����X���eS�,5��f��sŤ�'"l����o������D�q�A�%zQ����"����� 2�|�W��Ƶ�$��:'ڜG�������X���v�&>G��M_���!J8�� Þ����D���H�C��Њz���O����$ Xa�K&�|�㭌�0��I��{�i�82?��T`�f��@��F�٫���+<��SI�vtve�5�-[6u�({{���ɷҹ�f�Q&b'�>$�� ���&2�����~�DH��]t;Bз�g�˂�T�ê�u�m�Q�[���z��]d�j1r�sͧ���6��&�nU�j';Le?#��i��X3�:�ңDzd��#����N7���ޙ���	K	�؍Ý7A�Vh�E�Xhc��~�'iHX� �w���3����O��~2�<�b��N�C���5�o��C6�;�g����<=Z�J�����M������l�vY9�"I�뭜D��/������71r�;�N���c����4酁k�*�D��y�K�~X��d�/G��!�}�/���ջ�nݔ���R�%��C���*����UpG��2*rm�������}��Q^ҍ�<�9~hJ(����P%��:��b`�E�a�x� ׁ�D��MS�JǬ�ӢsP�^��0�/�����cݹ�}<l�?��iY�j�A�De��$�B�`��<�������*����]�8�'�;�_ފ��ѭ�RP��)��*\u�����M�uh 
�BT>`y�Ŷ�Ч�X3��s�x7t���L�
k��A��D�I�ZG�ԃN��xԍ"ix%R�͈�{|#��J0�QWJ����N7�[�?I���<���l�iňt	�5a�~"��3�J=����*g�Z��Y�1X�~/�ۋ7\�Si4:�#��${��d�E���?bpO�L��]f�x A�^�M���-}.��\�fZ�2p���&�����<m<.���̣�q.k�H N*k�e��64&��S�ʑsH��4�v?>�L��Y7b�ϳ�ep4p�o�b`�$�&�F�&�$8fތK
:�n���l��f�J��4�M������[�[U��kq=v���I\)�N�S	r��u�����5��EW�h�T��(v�G�0����-���rà�M��fE���Tq�����ЋWk?��\M�m���Wޅ+ ĎEr*�������l�`U�W$6��s)8gV���U�%q����K
"t;P�ɞ�����@:�-��UG��Mx�����e��6Z�if[��+�㑮����]͵g)��u�V�kt�u{5����p�e�an�j��o���-���7��"@�sZ�+�m���%��Ԧ��o��~)I��=tns&<��%�E?Gw?��X���i�-n��~�)�x���^te�9�z���~wI���	@�N"^�&�(l4H5SLk��n6\����6o�MB�[|d�TW����u���
7���$+>�,ց;�O���r��V�U`m�~�OH��"�85�x�D+,�~O�����`Gb����eRĠ�� |!~cl2�ϊď�d���V�5�4&d�`c��r^�BQnBASeŒC2���qD���|�F&�DDL-�丅������N�,��������mϻ���oHm�ڽ߮#�P�ς7I�2ҕ�戾�&��Y���ډ`��- ��9Qu5����ə��[���y#F�#WŐ�<�j�	m��lAS�f����qI"$݂��=�1�Y���Ҕ��~�_Oo����p�;�HH��5�r~l�w�q11���m�owߜ����!b�p�� %�l�	��d�й�(��09�	���j2�KL3�����F쪲,�z��ږ/x��j������$/�X�H�,v�Y=b7�a��©�VF�V/�ّ�k:w�L|�(ƚ���"�YS�ay���iބ�T��&O�r�'�eP�s#>�P�
o���}�mB��\�'{�V���o�(�ҧ�Q�s}����,H�9��j��b��zK�u�!\P3�>Ɨo�� 	&bR��1���C�b|�F�c��]"_�ɒrd	fͤ�Mɒ�"�y�T��)P*��kNc�/Z�W~c� fE�6˔ī�6:jM�(KS�~hL��X��$}$�0�p4�y�p�фq4*a�}:�WŠ��T���2��Ekn�U���ݎa�-�T������p���z� �{��z���۬u�^��WО��͠��*q9�፴vb���x��VӢm�m�vu#r$�[����IAI2[t��V+ ��]���\s��ߒ.��5-�:��a�,Pۥޒ��:���J�8�C-X�	��b�S�y;�q��z"�Kr�����ؠ��e D����=@�b��FX4\;�Z�y��P�9��Cj��&�N�1�]�;���B�m}���Q"-͗��:ka���X��G��i-��}A������,)�C���<�U�������=���KH�����!�nS���8��D>rn�{kQ�ޮ(����K !�R�1<�NY�䚎�A.���0�c����Ġ�b_�d\WC%�o�Q�+��L�x�-�4��-mW�X�T��Q����
��G�uy�X��*M�5�;�]	� jտ��zl��S���E��`�o�gɈ���!�燸=�9Hq;k��l�d.<�����mWYZ��5C~�)�]�5��/�	Oq�z��@3�oq!M�i�Ke^P�=Y�E�%|/�U�4	G�1Iο�\�����V���Op?�Д�<��F%�zl��"��4@�W[>k�t톮^��w�`�N߼ ����B��vt����>��������A�\��؆�[R�@���,7߳m黡���$]����́52�kD:<���,�hv�-*:����c�W�ΰ�����d=��i��hwA�_B�7;};���G���ө砢�� �n0`�ǹ��(���hQ�SWS6��7�u+	u���7���:S/��h�^v����9����f���2dNu�ӹ�r��a�6���;7kl:�����6�
<rq�D[��-�<� ��塁A���7P!UQ��1-JRo{ɱx.�`������M"�!�����{���v���(�ZrU�B0k�.���R�?1��V��Z���/9������L�(��f�[u�G�84���g��
X9��2K�:�D@�, �#���!Ǆۏ���.�Z(W$���g��T��n��fE��tyGhGڿ$T������y�چj@z���ۧ?�������͢DsZb����ff13�V<}]ʢ^r6�uL������9d�y$�{6h.�'��߉En�l	܋5c�q�'���!�{;�^��Z���F	��r�����"���HcuB��-t@<�e��� ��s��$T�C.l�"L�Ț΄w��U|�F�Agб�q��!��2b1��-HO.�1��b1��vv[|%���ğLt�;��AP���*�tq�Ţ����F���>Z������.�ɥ6O�F���V��7ԗ挥���h��I�G�wV��X�1L� ����V?*5��bUz䉐G���'O�f�����〒����i��u*!f�E�m5�j���dD�������_�q��2���cMl��16$�}+_V���N�NNo@~ʂ$��=ݲ���t�Q�+3��!�K�V���m`]��DX�k���������N��k�
�5/��Rt�K���VgE>�Z!��!�M����D*�����=��v~�y�g�r������?�>����B�cL{�z�0�]��u��⢲Y1�t�L�!�8����dC0C��������˺�3�,f��;��d��@h=�
�ۘ�d�lې����֗m�*�2�*��(�T��E�;�\ԩ��`y!�-]�|-�@_�7&���ZNh���RN�P-v2�5�NK����k�V��X��W �āԎ5
`ڴa�<`�~��+D���,1��3;��E��ٝ�a�ǩ'u8��*�G��}~7nN^�g��Lsc����Z48��}j����~=FM�j���h$�Sp1��
�3ǥ��\ٌ<Yo[L��JD3�X'����Xb�J�l�6�x�~�l�3�ќ�
���@z�a����4+c�r��"��1W��u�Ui4Ŧ��%����g�L��s]���yld\��̥�l�|#d&��F��F�vHT9tã����8j�j?��G��R��秆W�Ѣ�?�ܚ�}Y|����)��p*snb�-�$!\���3iI%^C��Ԡa �o���DD�����X^��w���v�ӟ�K �=W�+F���C�E�ؤ��{M��Q�>W�}���d��#!k�֗�;�dbZ�h7 0ͷ�m�u� @"�}j���N�!əz7wN������f���C�h�H#G���(M�MWQh�	�/.V&?� U^_��0ҮL�Ԥ஠+̏��A*O��s'?Ll؎ 2�W�"���q� �$��^��W���=�����p&<g�����"�[��ւگ}ɂ	��.e�Ți��EB��B�y���2�q~W�P���yk���^�Ԛmq� �*Kc{�e�<`AB��- ̼�x�X��Ȋ�i���sn<�^UJV�G��8���.��Cy�[�8�~m���J�:������SQ��%MQg�A�[=u	�����.��0�mѴ'�N��ThĞ9eެ����:�������RA(�~���uxb�3��1�Õ>��V��B�Z�zt���8Z��A5��iQoY턨C0}i!�	�o�>����?G�N!�Wk�T��l��ƟnBU�	�.���,�~m���P6��l�N1jw=�_&���(0�H-2x`3��Nc��vT,.������.�~u��P�f-�(u;�Ѥᢻy�}Y�bMD���0rdk[�E|����D6��Β^��_��V�;���/��F�!���Z�;l|ovK|K98>Gˑ�"��#l������k*�Vd�8�M!����m�C׍�W>i��o�z���Ů#�7q,�O��E-�ؐ�*��<l���>Z������+	�ּ̊#�P�r�\�Ɠa����~󩜵�i���3��!���3�D�š�'���<uP��1<b68�׭�E3�]�ѰP����8jS��w��mw���<
h%�j���=���	|D['!b���{@J�<���^i]k6Q�e���!��*
�{^�#/�G<~@ܔ���,8�l9��&��+�)#��>������Uk�+�#%O��y�
J�k9*Pa�]Q&tx�^Ą=������q����Y@c���=]�u�T]J>q�Y�Y�l����R�����U�"5�#�L�ޏ�̣� ��@+o��H��X�I8&>2H�oh���s>����5��Od�"o�1�Ŷ���Q�C��+˳@��W�wO�r��ťp��H��d���`F\Ֆ�ɸ� 7�[Tym�����!.�d�Kԥã��DJ[����W��dE£#Ȟ�|�9�5N`�"nl۹o�q��g��w�飲Hg�	���T����DJ�[�����c-C�x��I(��������=�>7[?
k��4��-�K%d��HV�^�����Ka�"2y >x	�հ�$�ކG#%\*�lDm�#�j��}~�3 ��fp���T{F�>���ᾂ
�(GF>Zo��먀�����؄��W V����Ww`�f�}��K/K������#b/2���g�Z������"K�?2W���8��ˊ��=���G���T�?�=��R����:5w�^;ao�S�d�a��S|��WćAi ��_�e\�5�\W��m��{t��w���g}u�g$����o���}!T}}�>\�+sG'-M�m��>lº���cU6�VE�i�R*9|f<,�\�s_i�I-�#��'�9��.^�D���,)�Hè���=��i�&�Eb��C7P��X�����>Ϡ�F��h��fd�|�V������y�h�����D�ԇ��x�.�/�#��s?H�yy��le��8u�(���.?AޅP�.��_(��|˧���� ��q�ǻvƛR(s�C3`H�q�؎��cZ��Cj[�)��v9��>3`f}�T幝̋���q��3�.6}�r������CC��vRyo�P�*T���|!�b3�l���06ω�F\VΏr�Y�
�p���m8x5�zB�y�<�~���WJt��`�*fcQ��c-\; ����U�'1��P|��A�dY��g��n~�S{���dqK�s�a �r���l�Y��4�������F��6}�vX��¥S�]�I�b�=���q�r�/���un����so� ՛O�.ú_�R{���Z�a��+�RK��y1������X�[�q�@�qilɮ���-`h�c�^}|ݤ��ҼF��!����T�/:�^;��M�Q���G|x���� {_�*l�
�v�2�W�����ąM��U �FeEF��@L��z:�z��QBF�-������O	m!�|��� 0%W?����Sz��i'���{Nʭ�π���l���Є�ߔ^��#�-��/���Q�2�w�Od������<-�Yq��|���Cuvb;�ΠR�4ʁ';���?2/�����Ǐ�y0дCF}������O2^�a���)�������7� ߫R�1�;4��]�:�4�H���ڇ�x��<Y�D�;cÜUa�����=� ZX��i���?��J�#�2��� {�#�[,�?#xm,��^2�R!@Kާ�o/�ި2��'���1��I���;��A��g7�n,����-�Xad�����)�p�h��(�
Ӓ�lY9w��V���XQ;N��a�m��vL��J925�ͷ�(�m�4Y��m�"��+A��`N�* ��u}��o�`xJ1&��P�Kֿvg��H܇�@7J~`[�/>�Y'�<�2�pC�}Uh��u�0����RK}��#�\s��7;�T!�##�i�0N?rz�Z�xw��L����ϔ� N�Q�F�G �N����?ų�M�dv�*�!���m[�����S��y?]}���
O?�6����1��_&S5۶EE��[��ȴ�`K�|?��}Ē���z�xmY����L���,m3d�i���f<�b��w�β��u�z	�������Vї�5�`5nlf�Q��|�n]�1L�CA�ˤ������߳ I�ts�q�~<=�s����z�,O��+1C�;����i#1zV�>�T�+A{/T�&*�3��A'I{�]TZ�P:�������|�Uݟ3�ú����j��O���Ȗ��X{���;
^ƛ�G�{��`�9�Į�K^����H�����@�H۽D���V ^ g �k����ȭ�Gᮝ����C�Y�����E�$���x���)��7Y ��z����e�.Y��(Y��^���� ��W��dЊ83�ߓ��|�Տ�1Ib��:�gG��&geC?�C_i�������6�k���GY\�_&_�K����Z����{�1Z|(�ڐ��I�}�nn0����Һ?�����+s��܄[�<���Ґ��p�g9����"|��	���_�z��NQ:}&�\0�x%l���V.�:7��	��&����}.ޢQ[o�9��<�S̒%4��~
�w &�݉�U������(��Ꙩp�)9)5)��б�:� T�N3�S��zۦ��߹��MxMH�#�� �� �C�������d.w/�qf�h���U���4�d<ηyٖ� ?nE�������H��Ĵ�"X�Yz���Tl�6�F�w�rA��a����%��X���U��<|<`��oA����#��¸j��q�U$��޼=�:MV�J_~GPQv�8��\'Cc��]��%2�����t}�J1�^͚"���\����}/DE�^�Lע2��V�5�R�d��f��! �.���/3�zY��C�����!^�/J�1�D�b���WoG�������c�描J%>Ba����:o��7� n�*��E��}-y9���ÿ���DT�$t� ���D��R���8�Z�.8�tL�e�]�(���j�Y�*���	�gv����o�����boL���&-�/K�3zR�*no���Ɗm#���%zʒq��a����9"rk�	pW`6v!rZ����Mи�e9�_�S��}x��>��	�y�B{��1w�0 ?ޤP���
�<�$��ʛ[���r�,��*c�g�E'����-D?l_YG�C���`��=�,��2.l��^���1�#s���q�9P���� ��f�1|#�+�8�S�����
�^�
k͡�ҏ�6�2&�b4��1P�|=mYɜ���Z/�F�Gw8�<�p-��~� $s;O�S��Uqտ4 �/��-T�46���Q˸��C.���p�.W�B ����Dk���2�q�]qU����E��
�m;E�[[����Ic�i�>x�u���%GЍEV�F(�𕃛�*������j���]S4��G+�B�gq����V�~�3l�ש*~QcN?b�K$]�c@-�ڼ�@G�G�.!���^
�@��)��d����<#=����N��7�̀ɼ���k(�XC�ɦQsծNLb/;i
�~��WR���EA��5r,�oC4>Pf�4����$���ߖLX:q,�@�Z�3A���M��P9�ΎrT��(|r�lPB��e7%l*|�%dG���R����8�����y�,�G� :��(��n�ۡ�
�0���ؘ	ɥP9L�k����螈��D��U������0\V�ղ�ZƼ: ���k��uVz	�Vco��$ĳ�3����2
-#�q@�: �$����Y0��?M�G��}YpY����|�����G�GO�������i������׵ԎV��*��C�
R�U�:�L���*Y��f�2��w��c��)qML��"��A��1�y�����c�������q[�o�(#��U�/`C���闖'�T�Z7��(B���A�F�ևݰ\�d2�|Z��ƻ�<V�O##c����#�Yg� ������2yJ$�7��1v�U���,*�慳[s������D<���^��1��L�}�nF���X��<�uV��9@M��(��1�������_�QS�/��(0�.��o���*�H�JN+�?���
_�`R;6�`a>_�� d���śL���m��{��	p�TM��۩�Ǧ��q�1�o�~��`�c�"}ۄ��`�)�C��S���6��S/�`�7�o�w�v�h��lR��xdJ>| (Ȣ�p9>���ɗ:�ҍ�g4��J��O7���-Oܕ0ӷ4a�^�&lKo���)��
S3�"��n����8�[��b�X_	���i�#}(\���	��&��(z-.AT�o3�!B%������zJ��ӈ 7��e��I<ST�� �ܫm�G�>�p���<?�YȚ���F�5�3�u8^���w7�5�����)�6Sk�|���c_N���E2���S�
�x┅�!�C�w�D�y27^S奁�|�n��7��
���>�0	�v�`��<2�W��� 7����o�@���>ҒWQ�Y��S����m%|h��C�b*gP��S��g���b��&y�>t
�i������:�J������̷��n>��x��|��K�	%Ku{���:eW_�e@���j�K~|f�>4�W��h�O9w�f�A� ?jEʷ���-2؟eY�F��c�M?���v��E?F��/`�A�%�=��<�C#^��\R�0#Lm�ce)z#sx'�4F��^�S��ڶ4Z���?ڽ�#͡G)��;�I.��r�[��tޒ��-�N��j!��t�ڙ�(P�����X�2'�C:��A�;w�I��a�"X��zx�a��}��j
��"D�v������A��y7�h4�ԍ�t/�M���l�y����a'�/`97}y܅$×��}�t8}�乊Mpz{T\HЗbb�O�	�w���[2�t� W~���帲�D|�ƣԁ�uX�H�\�1I�-��<º�W�}�!Ii�x�� �&DGw��q bC`�W���3��.���7�΃vOM9�����i�A�q������)�Q�] %��}���ot���-_q�x����Rx6�j�� -��;ۀOU�w�j7CrEK�{�����ֻMMQ�١�)|3� �3zB �����^}<i w�/���:��h\�R����g��	8	���=x��F�� ��(&���Q��^���ps���.�W�w~���� ;ʀZ,����%H��z
�ՉQ�+�.M�؝D��oO�Ek\�!��v���"&�(�D{b(���ۥ�1�r�V��vIX�wc�S?�I&��	F�Ev�x�4V4_�Jf�/������p����E��7i2�o[m�&:A��_L*y�?�/��ȕ>�A��ςn����@51`���)�ix'�tGZ�m�u$�8�M��A���!���kF��P�>f����*�^��T����"��f�b��ތ�����|��A���'�y�#�b�Y� r���K[5=�>�OC� ��>RY^�1��GA�L]VA*���|qjF�ޒ�oPx��'2����w���
�J���S�T[�@�>J���(�'F�}��C��AԄ��^��^�;�x�p�]�V��]ݤ�R�5N/��"�6������`�k�*�ŭ�yi�>[�<F�)TS�<m(O/���������
������N���Ϻ�1\���g�Xw�I���RTq��R�XSpʣ��bR?H��K�p��nY�f����x%�֢I�P6ޓ���a�Սz���+�*{����1d`��d���{�NV��Ї\+=�'�2d���b�D,dT�erj�> r�?R�ß���(CL���})t�I�n�9<aBt�8�/v�'x��P����5hhO�,���!��zn�C�6ג��k�:��>�7St�7�?�����!��@�GB�b�ց���Z���{Tʟ�����=��&�XM�q��2d}�zYMʌ�{F^����,@�e�br��A���<o�((�_/�� 5L4�As37��S��h�S�s����,\��ܤ8R���x/<4&|��G~Q0X�n Mm�n�� )5D<>����k\�D��>A������1W��H!�� ��?����[���i�ep�ڄJ@+f�92ؿ
�J�����f�$� ��S{��bO/��2�J�0	�]���6���G[@�E�a���e+��(��D�,OWmp|���=A��xv/��{�� �ނ3�c�ݍ��<1bZ�XjϬ��ϔw��ܷw�5
`���r�ԩv��پqF�	�Qχ.�t$D ,�K&�bF�Y�,��j`t��[Cz��̚�E7y�q�TSiN�_�
�Ftu||�0�����_q	�q�?�-���r�c��2/�e�sY�t���(�1^���ǟ����|�W���xp��[=R����m���C��j~P��;r��Q�oS����������51���T1K�����u�1+-�A�"05�
��z]AAb�:f[w�;i��Un�
B���a��M��� -�s��Y�Ҋ\9��~�C�$�"�)V���5�>uW1�s+J/��!�#P��I��I7/��LAk1g�5��W,�х��bft_�����_o����5��l��c��!�TAm�`dGC��}ߙ�w�@�Z�^s���$���� Y'�,"ꋪ�n<��rУ�)������Ԓa(F� �����
Zmn�Ȱ����ȗfpW2a"s�Dq�bFH��	Mb�������Tb�jJ�'�+�p)�m��xޙ�i��	{LU� �姻*�h�#�Uw{�T1�YpF��1���n1]�1��)���/DN�an�Щ
�1e��j��t0(��*����$G9�|u6�Y�ȴ"m5v��G��-�h�]�A�7��{�v�.��n���6`�7<ڇa��H�;�45!���R<�q�P"Z���ִ��l�e����oF�U#�R�#	h��c� a<I����è�7������0�r۾Z�,��W�F�ɛ�A��\�o�z�)�B�[�n&�W�d��8T�N�
<k��|q�(p�2��&��o��J�q�Fz;���)���5�6Z�S-� �S\4�>�q�ցЅ����
�����g���]�7W�Ƃ[�V�'����Wj�n#s���#߆��tUÞ<����p����5K�lܘȾ���1�����wL�L8@q+3VK�$Mxz�7�,*g��J�l�;��|i+����!z�LUUv1R�V�����b�]6�4���u(��;��U�ORx�y$y ���~{6u �NGs�%�?�M/��qE��_u"k�რ�>*t:���q|*��2W��wVi,OD��,���3�;��8��`w|���8$η����H����k|�*%�ģ�ڭ����(�[�M���_�`�'�ďn��ݗ��͙�R5��b�>�YX�BZ4
7O&��\�8�9�8��s�u&��;��oo���d{�rS$s�>(Nm#B�6*>�-���)�<fȟ�����T�;�oh��};@pp��PX�8f�6A �qS:cLӔ�t�縓U�[ՆZ}+���h|�_1�<A�z�+8qC�chтf�_ݸ��4G��u�|҉l>�|���V�L�͂vw��~����jX�x>�d���X@`����_T����sI� �����c�/3)ۦU`�\`�3�Np-Ʃ��F4S̑���d�ם���߱6-���/�."nt����-_[rö����J<�A"?��m�ҙ,V����Y���DF�����|
)���v��dx�g����5@n�k�I����*v뽭�j��ʟ�����r�݀L�FҨ��:��(Fs�M�z|R�;	�C֭��\����1�E�S���׹�V9NRC$u!��c !��yiS���1<`��J"�o*��r���7h�ސ,��%*� ��WCw�'���wB���LX^W}0���0��@y�S�Nm^z�A|�D� idt����;m�&��Nnj�_K���̟D2��$ƇaL�&�����<kO(9u����^�(�A�'a�����¢-+�<[y�S�u˪���߷b�HN{��m��a���:��Z:F��`΃�bp�Ml}���4�+[&�pN;�����	��,J��a���M�ur�SHQ���0zD���~#G��S+�l�}��n���Aڒָ
h�'%���$a�����@hƗf/@�Π�kr~Z�/(�P�띁y����f�����T��?�pOF�S�dy�ٗ�Ć	�@/n�+�h֏�С��՜�rK�l��"��P��x톰I`���ġ��L����(+���Ѯ�N��Dc/�H]N��W������ȫϪ	�:Eh�F#
�~Ӈ�UȰ��"L�KT�ߑ'�⯝�Ч��߽�{;!wп� ��!����騢ED��y�<�9�\Nx��PX�Lu�s`U�l����H��[1�������~X�Δ5��*�@1���i���aM�j깕�{�x�/<B�s�f3�����`�^����b
@hc��&��@%x;`��5=�������lI	�����@;�{wd�63�wp�z�ڜ(g�3	Q&�;�;w���_V�a��?7	�)"3 �ڂ *S|�Ք��B�Q��X�5N\���"^�%T�T�(���|_׊�*��0�D��I5[�9�����i��Έ2�u� �㇙qO-����� �$E_��<P5����ؑ������NT�����}�$�05-�r�ľx{��vl��7�^4���.y-���N�����q-�0q��iv����ᵏ�2���M�N]�R@7?P���m�ǚo���J9�	�8�Zt
9�V���+x+� �1u� �!��Uާ�Z�~��|����8�L�_��!$�l��a0=�	f��+�V�����g�!)�Z�f6�����ʲ��I3�Ո/�w'Php���C1ؠ8S���d�g=~c��X�'�S�-��.c��%�����.SY����G���]�{�@7��g4/qp����L�Ö�:$�4T�*�00���c�lr-��Řa1q��� `���0���@���E���}8��s���"H�oq����Y�O�Ȱ�e%�T ��eƳ�=��LO:C���etŅ���]�B�	�e�D9c��F����(�X�7	�T}���de��0� q�v��$!�%ʭ�α�n/��SY�M�B��m�z��X���}S��:�R/���0r�ە���CS6t{���x�I���[S��;U�V�nhO<J,LY4>
;cGǼϺ]q���.���n.	x$\J �~xZ��J��S8˻���(��1����&�b-�ڎ�5D+��i☒�\/�=^�W���?`rB
77�δ�fRâ���s'���90� ?}���=���Bo5�¨�4* �K��釣�LM�D�}��N)~�$#D��K$��A�Q�!�d{�'������D{-U&24Ā�,S$��8��t�o�C~�ʸL��r.Rպ�=�No 7�LgC1��o+Kj�ɳ�g��4 ���sX��ئ!h+��4�}_=��$Ҝ28��Un섄e37K�_iZ��g����,<�x9M��b�
��&��E�"��,TNA��:h�܏�8h9C���tK
�`=��h�C�N�t�Uf毢�Iq�,�C��zQ����-��%���E� L?&�?���K��ɘ{����	k4;�5���8�pp,B>���.��\��G�\F��~��:_-ѫ���IE�,!=��kdm	�6��щ��r����ilM���'
mk!�]�el�w���eQ��x��d���~���Ȗ�����e�ПA��`��.�ߴ����l�K��3/nz3]�.yߔWy��$��OS��_�`�\q��O�O��-eg�!���'{��x��b�S!��*u��)1��@9���n�c~�I�r���1s��$�P��{%��gξ[~wM-�i��iW�컶���� ��CI	��Mr${� !��^���N�K0m���ờ�t�33y��9���~9�^ 
ƄI�������o�%4ު@���/<�v�Թp1#*%��Z亷�Y�WQwJ
T��D+0�65pu���_w/����e��0���{�dL�oi��	���������A���8K���q��nf4��-=��a-�	��j�{ƙ�]�v��@:��R��G�pk����^a�5
��4�u(�K�.7�b8E����:r댫���Iϓa��K�$5ܺq����!B���7�}2�;7e$��g��%�N�Mqr$v��l�u��h�C�}�N.S�`t��A�O�p|�v䮔�6�Pm�c���G�bHSS!�wk��3��:�ǃ����[N�TM�oh��қ��՚�~��DSsZ�n����|wtB�cmir�t�_
��ðHe4�z'1�$�5�m��MO��K��r�ڗp��e������},�ZG����l��o糬�ߞ��@;����@S�<]3�\&��D*�.��=OP��w�yě�hWw&�x8g��Cu�Y������@5qQ���C�PW�G]��] [koQ<��Tt��@���bl�T0�nV�8k��0S���,l��K���ɺ!��;Wzⷺ@ t�����J��Tr:��G�t�~�o��5@7O�jJ�ŘT�"��FDQ�7���F��LpcJ�� ?����������e��C�:�9U��~�u���s�V�����c8�ľ4_Q�"��ڱo<o�����wJ�a��Y�0v��zz���BZ$K����;��oC(��ӑHZ��h>�k�@վ	4���*����{���pg��l*%w��?��aC��6?`�*��5���I%��y�м�Q	��R"��yQ?��<�'���Zo� ;h� e�CO@-���	|L1v���E��	i�R1���!<��^Y���L�nK��k!(>Wy�::V>dqϴ��d����Y� `�(����#M8����P��^�cIǚ�ί�Q���B�q�d����<Yk8������(!�L�����Y�;1��J�$o��c�|*�y�nB�g[�a�	���3o�WmIF<�Պ�����$�������v�����8\_XY+d����;E*�-%��im��Vh�I�X���v�Y�49��+�`��K &,�4������g�գ[�l�)���e��>ۄ�:�/�Ҕ}[D���J����oA�Y�0q$Ĭ�_�su���@>�*�����tÀ��@R����gF<E�sT��m^�4��C��7��w���[	�!/l�cL�Mv�̯��x��E�wR���h�c�nJLf֖�n�ڽ��aM��\�N-?m)6�¸���qHi����s�+d�ӑ�_t��Y�_���3h�ۊd��L�M��W����V3�Ȁ��r�Ŀ����&&���*��X3��g���ut.���c�-�m�SN�ߐ�$yQ���V(P:$C0���4��<���]�n �e�ƺ�P�S1����������(�X�	l@�Lc�@�x���)o�nٓ:l@-ՕAƞx��ʣ2ڟ݄N�6���b#C��@�"l�ʋɉ�d��C�z�o��������������n�䣕M�c랣�u�rPl��U��c^��e���l)�h�g�vW�z�>E�������Ox�]cmgX���1�TK�Fh�_��~�Ԃ��S��$�n�:Q�=R�O�e�����Jm�t�����J����P��}�S�=�ل%�9/Z�+xR������ےh"�K&O^C��`� ��q��FdS^$�x)X�!�4E��ᡶ!�P�`��d
}֞���u���5��n��R7�=�F�;4��՟��Yt)z*0/�S�%����>�7�}�%�[a�[��!'�s�Ʌ��N�����O3hi��Pk���0�����\e22K�W�]#����z��3W$��9�\/iCrx"Lv�_���f��gy��۶�s�t=�~��vs G�	Q�	��`*�G��\U]_K�	��|��@3���	�1�e:���ʈ�q=ב��	1o�̿�4������=�jK8jE�X|t�;��lC�+ݍ��đ�d8�
W��F��t"N���?jhK,�����eLm$kC�9Ee�B:e�w�-#���;c`�xc�ʋ"��|���S���DY��mLVQ$_����Ol-�V*"�`uoq7��^�f�M��g��x'X�ͺ��X���M�a?Z�zd��3�0\^�!O���i���G��T�L����I$�3D�p���bΐ�T�O^��Ş������\��̜���3��DS~Yn��5M�q`ا��h�OGuN�w��#q�,��V�s�E��]>P��ZZ��D�2SK�*�n|7�m��ƪ����ZǞ��褛�X[[����|�Ot����M��="B���n��}B��(�U����,��}Ǉw�����������k�l��~���^��pGIE�=��5�M_��*�v�h�\�Q��{���h���"56��e���6i$��sE�;�*�����v����;"%���T�v���Y/��o�����yr�x�/L����QQ�[�鴂�*��"ށ|@��	��*WJ���r�4��X�|u�t&�m�M%��Hj^@|z�,�F�W� &�u�	8s�OB��t�ʄ�rސ��B4?76���Y������9U����F��ŗ�)����4�2��:��\I�?��^�]ō�>!I��Gd��R%q��	$ť�%�ea�\���mF7�Ii���wM�����mAm�8�%��wx�_y�������� �?ptp�!/�/�1��Q,����x�Ə\^{Ty��6�M1����WUs��N ��x�ؑ0��=�f	[re�^�-;�.
x@�E�>ʊ�+�|� ����[<��^�e�;��0�bl�L���]��6��ֹso�s���kֶ�\����n�;��W�Y�A�����\�d��,�)�\�~�EH�*Xq7�@��]=�H��@&oH9L6���f���q4="�������4C�\���_���gh��R��gĕ�ٰ�z��13,���Jj���D��bbXͰ�tx���S��|���we��o���g�B&�£�ʊK�{@�����m�9rb)�A�����l�J���tTu�~������z�������`�s[	B6�|��oY�q̏�.��R�kVP�J(V�a�f[˳��"9;� ���d�{���۝�:�ZL@2w�[0��~As�m�0��,����"�,r񠈬QS��v8�R��kه���[�����(L\"����O��O����,I��9���N�1����E]�DW���VC�Z#-壋M�.�_��N�������yGܮ�&Y��qi��u��m��sA���]ͦ��N����@F�����&H�]<O���﷦�W��c�R���MA�֜2b-�N������D~���˲a00U�=+�_Z�5N3[��+a�gs�n����A�ezq��U���Ki�/(�k�3�@y+��q�k��]�����+�8B�?��� үV���g���7Bk���7�H���4�5#�1׈$T`�(�v��%�, ���l)J6��W�����p��
��L��������m�plۚل�~n^k"!�� �%�!���l.��;���O!�6C�aS��jW֎]k����哛���H������$��H�1]TC=�
�"�/B[���3�e@�; |8F�v
u�ްl��?�<%�C^$��n�eaX�m�U���HrY��#���u�fAY*�%i9"/�%'��V�"��D�{�+�E���&4N0OTC Z�2��	S��6��A�s�p��.�X�G�l �axn�]W07�RF��	�����S*����0��Ʉ%x�� ik����*�I�E�o�z9��R�40�`�s�n�W`�u�)�-Trb����S��l'	���*YA�u�>5���gp�gL�k��kW =,�q �uṘ�@�wd@��LCE�r9�8�}@�
f�R:�,�����o�*ʸ�v4J&>�.��D�R�5���h?GF`����~������ ���8k�D14����PƦ->LJ������m�D�^�E�ǡ��I��)�����6�Y�Y� ��ڢ�s@���*M�3�3iT�[�#OPɆa>�m�K��A}U�¬5�rDNr�>a�N�ӎ��4�D�to��dV�bQ�z�O��C�`B��H!�#>�]e��x�R�<��Ծ��v��k'U�l���*��mI"�i��P����5q�}w� �P5�T��O>]���yu\K'��s�n�=c+!�*�[%�1e��|<�>�+�:��B*�*�O��A�R"�u�s��F$����ߙy���N��S���٥�V*߻�mi�'e��L����`Ŧ���I+�\3�v�/_�1��Ak��d�I�t��Mm?>�H�\�+�f��H�{�{��ЀT�
�޵!56�=�o()�/O!���f��9,�)s#@�fA(�\�)۷ߏ�� 
w����J��iP��]:
i�����ƀ�_]��8qo�"�G�C��_\VF�,MY��h5�i�z窆S;0��@����W{n��Ϩ��ii�D)ꮛ�}�%�>�DX����ׄ�]��I�O�F�ù|��@[��b�d��D�ؐ���D�5@B#�ѩ~a?<�G��O��w�g�h��"J聂<u���59>�Yu��؝��o� b���g����Ru�R��V�,}b��fhs��g�� �N�:���O2��̇Y���� `�z �[�l��3��Ѧ,{�r�b@$B��������Fɥ��o��ҵ�.6`,>x��W�5)
�� "n!v�I�����7��{��6�^�A�4gu>X�b���kv��;�O&��ul_�B]긌Dߢ��8W����������pN��v��MG����Aǋs+�X��me�P۞�Ƈ�:�R�{��a��>O�h��x���������{1�<����l(۹�R�i�w�~c����Ȼ�d'���)<Q�#�^�W\��:� �~���
�=q֫��*�xk�mM��@y�����~C� J����|ɧ���j�מB%�w�Jh����&�&���_�j"/{P˾�m��H��b��"��~&��ٜ�[�IM�!�_�t�VB�2�+r3�awn�<�瞱ש��)&��e-&����Y	�	6%<o���b�|�]�� 8�
Gr�X��fHh�u�(R0/)(}��
�U)�M�6�t�~�H�X�D}���¹�+�x��C��V�-(=�`��8
f^ ��*�r
4��8����KwN����!	��y}LOHUCY���;?0���a��)�<��5qw:�h���Џ?xC�3H�pHHn.ZP��* ���?ȱz�;7_���g�2?�Y����/<dW-�L�>���.��ܞh�b�q�ե��2j��w1C�'�1"�k+���22��������?�ޯ�����z_y������ �\p�.Y��v����i9Ft�L8'B���f���6�$5Y�<����3`�(_�<��a4*�'YHK��B�����I�p�ҏ5p�HA�f'ꊾ^�`r��	=6�FZ��g|\I�l�V�[E������U�����ۘ��f˄u20c�t�}���X�D��5 $�It��΋��6
W���uS��������Pّ'|>z�^tBpŸ�-�`�z����T�l]Yz��ǿE���{.�9�`#:�Hj�MM1�+�Dr<�q~i��YyĬ���'JD9n�;�c���a����}!�oHЏ�j�|�^p
�R3_�m�Qp�MCk�&՘��"����P�o_���b��J�B�/��1Z����ĉ���1}B,�6��L��3��E�Ƅ5vDu�E�wɆ�#��بי��#$�B�M��)�%���U���n�͸�"Ӆ`Ҟ�Gn{����3�c��	{�����h�;�%�W�"��H+�F��U��.�;���&u�6���wPfK��H��k�!��)��ؑ�-�]�0�,Q<�2�^5� ��������On���2�1�;�+�� �g{xR%�Jl�uh�*��r&+?�����l"劀�7�S)3

zbiIk�S�Gq�~1F�L��xB����N� ��Q;��00 �x��s4s�sZ����I�)9�95�}Yu6�/FSN-�jִX�nغ�T9��eo�����ȏJ���#�����4:�E7�$��5��N����.%�dy[+{�8NF�-<��<�5�[��p����0�?���=����5R��5�~������O���~`�e�����ʵ�]5}�
'��[�����*V�@��U���}�L���J�95 }]�����J��-1��D�B�iI��ﰅi$���>O��7����I��k9�����<������,P��)�U� ��y{H�%���N�O2@�l�EI�{��A�`vc=�����igG�ef�&�T�Lq���T��wWRdT�8�26�����27ܭ�7��O���~�Epf��ן,�ߚg�Oo��u�@S�ϓ�s�!�����#E9�Ҟ*���G���Ŵ|�!]��=����Cn]Y#�&,Xbq��)?�G������v�?�M�(8������F{����������)��K��R�*=_�R0��^#c�,�ϔ:��k��Ɛ=�Hl��cñ���4_�Z��s)�s���(�L���WSG����E���xaZ�ya�T��+!y.U�ױ�w���Gվ�iˀ�Zf�E�-���2���x�9���']�a�]G�߉�O�^ ߉5A���<'��4�d}���p��%�_P.�\�E]� �X�����O���%L�D�� 4���6�L��䈧ϝ}�-[�)�e�J�REAP�n-���D��u0����O�㹻�y;���盟s[�'�Xf7��b�uPK�M� �
6|��^̋�v��~�A�}d�ė�.����`�F0�^4�!΀��+��u�Չ�w5^��(�ϭݳZ�h�"R�WcR_�R��Xk[i�Y�~�.���|���g����t[�4�߃�@\Pmp=^a69�2�u�W>�rnO��">LP����]W���2�.l�L�"Np+�o��曻�����BZ榛�L�c��I
0���7(���2�,��S�W�e��K3����$V�Ք�K�A�p�{�caq,RDHoS!9��Q�>-����]�(���)��dM�m|I�XX��j��
f���>4*����r��P�+�I����´	�A ZT)�jz|Ub�Dx�52�M���5��*�E����u>Bu���m=���^���5�켟����T �K���$ą)����h6��_s�ٙ�(aZ�ľe,���%�n:l�u1�+ԅTS|]"�rel03�ZT=ﲘm��0�i�՘�.#R�<9�'�+e�j;'�D}��=��iXs�⫞�I��4v�6�q�D�Ϲ�uDM��.z�Ŕژrw�k[vq�=|��M����T�B��d(^n�M��2}m8��=�"�=��0��/���}}r��D��R�!ު!�K�.f���7NBG�6N��*�5��+�����c���r�Z6�t<��C:H��_�˿���&�^��H�ڿ��0���`�4�<DӚ�v��V��\�8*v�������8��Һ=�	&��>,��k�(=�>>��n������՝< ��0�6�+�7,+��Rh��
��z�.�ֈ�ȴ�bc��K����;��Q�D�١��:6�Ayn�9~��J<ƹ�#y1��e�W��HԒ1��U���}�*w����B]������W��>s�;7�Vf#��vp�	W=KW������˝+�,�H;�5������ͮX�`����(��0����d�����
��߮��ENTԦ�1�$��YK����0�Z��dϵ���|�~D�'��p���;�������1z͜�H�#C:?(��Q�q��ec��|O�c�u=-�|I�?jҍi�
4�9�X/m�t��g!?ze��Q<ؔ����%��Ѝ/��ً�Н�M��D��>��{�Q����=ɺ�'-��9�Kzc�'�HF%��gLm���n��E���A;�ء!�ŜA"k���J�-p*<g�dGav� �Î"\��C�
�/A���d�͡?7}%
�9mt�+.��0�K��&�R�X�B��9��'�b�ȣ��3��ٻ}�Y�pHK5�0�O��q '�]�����Y��[43��P���:�ˎ9���㌍��_�)7�O9VBS�5	���h�9g�������4L�qq��a���M����*u�Q�fb��{<�����`�q_�����Q �Jيe�Av���2p=���]#�U[�.�p�kx����)C�V
>N�[ᕪ?۽9$<�>�҅(�D�z��Ra#�?e�{�Za 0���]�ۀ�;�=^�j�!?��������-����GzC!/ѽ.�N��cU_��Y_v��D�[��h�pQS|cv��.��8����Q)��ˍ�v|�"]Ղ���!��$qn6G���������-�S�˒hD���ݸ�]V�]eg���w�M2R��w��&����\�D��¼�ׇ�fYr�<3�& U[0ZΜ�rĳ?�g3gG�?1�dW~
����^c�K8ґS<D�!t�d~?�X)|=�L�y���P�)Z�UF)B��~F��y��Ͳq�)uz]:���Ն�OU���c��*u�1��j"k��!'���u�|���>�GjĂ �p`c A�%�	��&N@т�$�!��e!�ֆ1$Oj�|�;�>����l��`7�M'�3b˛5{��^-��-��I|�1�RJQ�e`\��X[Oƥ�'�Ii7�/�����NkN2��
�Z:��iJ�8N�w/�%6'�8�
�#��t���@!��m�*�d�S�U'<�S=a���6!�ό��zy�!:�jfTV�]z����br��<<�SR�XP�"��
��2�(�t���ҩﮣ��=M�	1�`� )QF������R�S�l���F�j?�N5I�⭛�ym�����H�]�u�%�������ip%��uR�D��z�OB0��O�p/'.)����\��Do[�S��|�C�9
{J�/~h1�O�ZK�u��'������;Y{!�QzfXn\��ӈ�:�FLk}��t�>���ZTP���s&�u�u�אv����	[�i�%Ra�f��)bA'1�[񆆠\k:4�G�f� q�<ci�}�7NS�����rvF�eָ&u5!^S)@h�|�'�P����\��w�A���>aĝ\~T�8�O�Se�1�g��;���gJ���8�6����&)�:?M��by����h�;=!4G�aH��J/sB��p�v��@�[�T����9�pYZ!�� �H��Xb�&
E�d��I]���L�j���9Y6c����A��eJ�a-��YyC"�j�C� �D�-��Hg��u◜~ES�Y�C�?`.���K�U�C+�Ǒ��@�a�s�R�14#��yF{���a��'��E�hmٺz��P礡z'�Q`f�i�g�LI��o�iy;�W?[`lU�ܯ�A?�(|*cAԼ����*�ތTt���i��G��4�/Qh\`����x�BS���D<AK�ޫ>�˾]`u��24��Ed;�`�Ӄ
]yF�f��y�=%�2l�"�z��]�T���L�s�qW�k��
�`�[���nX
1ga�6��X�EێR����~�){m������wq��Ё}���,k%7���^��<�G ���5K�%��ѥ���̑!�rY�����zH޶�d�_��7���Vhv��;~�	���3$ �/V;b9���j�dN햳1�.6[[�eO(N�J�+���B�-	+�D*1|�*QE��b����(�Gt���FE;q����n�'�%�_��zk�p�{���fM����Q����mp�c��|�[���gK��|�C���e<b��n���:#%�N�6oH$=�N��y4�ű�`!�/d�<��{Nw}�5
ɲ�mB��W�����ru��6�z�Fy�ͩ-փ�7���f�I(,�bպ��`�-�~J�f��8�B�֏1�"�<dwz\>(_�T��\����Moyw���s�h3��x?5�rN�a� ��3+��	����T��/�:D��X4����	���"��qX4��æ�o�l����e��'@��f�5��^�����B*���S�{�m�]��ei(�Ǥ��?�i�?]@��a)Q �s��΅*9��^
 J����IuCmc�9��q�դ&�x���b7���q����l�>�����?�虍�Ntmڰ�F�!��A�{�r�2e��x�=7�,n� $�X��]kb�@��W�h��W��ٕƵ��ǡ�H'u�߫HZ���+t e�uAGQ�H}�t���XH���"!aP��MU�Φ�CǴ�
�`��}�����g�쪛Ր�&j��&�CE�rR�`n��xl|�u�)<a�BH�6j3����n��s�X������]��u[A.[`�t��EKd7Gu�g�L�K��]΃c��Ͳ5�}���ޑ��t��&�ѳB�ݙ�8��z�*����i�Ƞ���]��٤���92�K<}�ӗ���S[���O�
k�C��ee�E ��T����IF���5�`�(:(	ye���#��f���&�x��vC�~^��i��Y�;�h3ȪmAq1���Z���IR�kQ��L�P��2=(�)+
[�����B8����\K���H}�ĭ'�M^�P���^y�J�g�_0��s�.��8sH�%&2�UƎfg?"Z`��s�����	���Q^��6c�#3��y�	҅V��&�h8F���H.�|��J�rH`N���ì������^�����0:�%K	w�V9��9K:�g�r�]_= ���Y�Ivg:�7�����G��q�������㒁z��cd��!2�y�`M���V���w�*;k��X�IS�_��w�Ų.���1vff�	M�k-xPh�t�OF����se.���W���T�.�
~]�g�d0Xi'��=g�Q:!�U�킦��sVیo����O�iIw��E���u+k?��h0H0���fd�^f�L(s�F�FE�dQ�`�X�k�V�-"6�O�ÅT�"��l����&-~�_:�`,,�ix���z^C��6�ϋ&�9Mm�^hE)�@�q'�ח�3c7N��)�n���3!�+���e��&WO�6O�	�G�z�/��·<^$
�A�rg�	���fm�'�exG�$N@틻ى�������}3V������1��M0>.�$�%�W���'h������R,�pR��D��t�)C�{~���u4""f�!���8�ި4�����*�eL�^�I�{���*��WoN��#t�f�}���a�;|ߊ�*�]';�TJ��Va��9@b� �~��A�_0���5�^��l]��	��=�d3о�!���Cɖ�����"&k�5��%P��p`�(w> V���=���R��覝H��@���ܣդF?�����bu~������mGE[�o>�ª������{n���3�'ʖ]
�6u�a��CM�9��u�Q�#�ӌ'�������+/y���[�[АQ�~'Yb��ა"�9���R7u:iqЂ�����^@oPu�R2!�Z`ͬu3�S\�$h��2�|PȈ�O���>�䔾��(9*}��Yex�\��w�1�7+%>��vM����&��XH��1�+�ӷYF��,�x���z+��@(V��4K�AbX��Zw.Q��0�kN� ��O-�O�JP�+o�+2p�2"DG��8�{���N/��>wͳ$bzV�})�ױ[�"�$c}� s�=���@g���6�� _Y����Gq�VH'�{�M5�"�%R��;.�e;%����ea[��G��Wܯ�3�?&����{��v�y��z��Xr���eYń�F_}ܠ�
cڼ�im��[�m{s�Ay:9��e+�;�m�sa�^�}2-]��GU�c
�l}��sh��b=��@�Rֆ�*��X.Qu��<,�[ps�F�U�A���P��Vq�@��̷�R#�3��@�0o���8
�hn��?���-@��܆��u����!�έMs������?��;�z�(�FHʹ�߷ "�iÆɝy�4 �H�T���x�?�����[pΏf�Ǐs?ť���s�OP��y�i��틊8��&o7o
�\�����+H	��"�gZ u�� ~��bK���~��C� ��-��D����nM�"�~����_732�#~����$jɌ2%$��q���>��Q+������2�',:E+v]�._�f��j�w�K�z��^w��n�̼� �u�c�A��Wy��ɸ��e�IWON�l�e�T�K����IX���MS���b���؜�k<^��"l��Li�N���cY�ζ�Z@�!�Ў�(tZ8�x�`"p�x��#d��.��OҞ�s�$�5�eo�(�(3�>v�_[���_������-kT��%IA0(�I=b���E��A���ƍ�R�Ր�)A�Z�͆nj�zFX-J�%Y��V��J��z��I�8�@�YvF��8��4TU-_�H x7�2q�pj�!�V��zI*�����:>��m�0V��vzu����H�3⣝�8��@�xfb�H��Y��%=�om�[8݊�Q���Jd�����\z������<`��Q<��VE�d�3z�I�;�����1��c�fxW*�p(
�/,�Я���"��]��h�Ȑ4�G@s�o�Ƶ��E���ӑ����i?�O����[7�bM �:�j���(D�Y�/�����}��u���i��6���|d��j��+�
/�6
���	�#�A����?���B�uT�M%"> ]E�ba�������)���y8��S�g�I�n�>9�s")I��F	OLo�{J�.9X�ܿ��>�L�Ʈ�K����a����8+��W��8�UDf0��&�#�����4Ы&�H��1�.l����>�+���5u
��������0RsG����YJy]��bl ��	��k�_���M�D�R�X|<Mv�'�+)�:}��� �"$�]5�����XӍ8�ޢ�f0M}�zh殡�+���yƦT+Wr���M^}���s�/z��x-���+�g��$�_����C�ِ�{=z�W�6G� �w����@۩�R;��<vtWt?�:7ب�����)���z�c "]� )n��hM@=�~h8sY�>�q���7T[�y8��j�S��T�m	���9�;�S�E8���7��,���$�0x�*��ѷ�o2��������I�'�H��{�Nc�~�G��~�@�<~SPXU����7CI�H_����[2�҅+2���C��`���g�ۄQ\����)tV	o�ȴ��rS��&����)�Ѧ�Fn/����{�,�K�\�Ҟ��YI`���q���]H���旒��Ic3s�O<�^������X�H R2C���?���I(��#�Qn�q�M�X�ԆIp��\O��&a�f%^U����1��h䦺�fo��a���\_TV���"���6geF���A�2��Pa��s@���k����%f(���-���gu[8Y:ri��;x� ����Y@C�l����]���_����Ck�� �Fi��?����6�?c?�vTl}̏�H������fv9RR��Y�l�g���ݑ7����+sG���sh��Lס���GR�}����t�i=?��d#Z����բ�x�%kĄ���v��T!����%�G��[J-�>Gl:�b�s�h�\�mg&�k�~�O	,^�Dq�d���u�Ĳ��Y0o�����I���<����W�*����6^���ĒN��FS���@$�NC�X�w��t�l`7�-���'$���#b�j�@R�'v7g�{��S`p�a.��:ӫ�N��|���G)���"$��3x�p�PA��w����HE��U�������G��H\���nG��ồ���w��ޞ�F�W��kOl� �$a1��9�
�j,`��L��Ǚ��m��N���NLbJXH"��@̹�b���"����QnW;�<��H�6L`B[�:��C��%��Ń�W�z�>��͚K$�"Xo�߬�Y ַ5p�7���%����>5 �z���(G����\�5���&��18�>��n�`�G�t|�r�`Α(�=��O��h$�a�aT��JL���t�B(I>� ۱����5ˢ<[rR�Ϣy���o���{;�d�R�l5���\������6��f�!�\�#�r���QM8�����F��t�t��ª���TB��0e�e�`g��16B�̵��N-����Y��qaUT|�
%e_���YG���; �P�~p���>����#�)_�߶�]aU�����	[���lG#���T�٪����ܿ�.�wI�bn,�>)&�xG��Yj�W�PK�-��ܠ�Ƿ,��Z:�6�D�q(O�	z�|����JYΖ�~T
�R�%�_�r��� 6��-�����>�17��Mǃꑤ8����l4m4��gȑ���0�uFD���m�k-����33�.����Vq2P���׃��y����Ͱݝ������P�a̕�n�4�SXD�}<��w��>�\^�Ѧ��S]�5�}1�T�S�iy�W.��e;ޠC)S�~�<�A!�}7YBͪj�'W�N�`|�?7���!���Q$r�����	Ђ\��d��j��oJ�i逡����u���\��1D��h�]�+Bp�F����&����5� �e���}�0sSUx	�
�?���?:�i*g>��2Q�}����+��Ѹ}�B��6��P(�'_�ҭ$�q�?���X��E��7��7>9��l(m�S��]	�@F7&6�,�D�t)��v���'[�	�h�B�-��{��@��#i����ҡN��/�z
�խ[ӵ�ٳ�P�԰�0�,��ц�e��I�Of��� 9��)��7�~�&s���3k
�W#�m�6p)�����C���x!V���A����cRZ���w!%� �>���$NP�H4�aɕp�D!_|����T������4��Z�ʽf�دZm���Uq�+�2�P;R�y����2�q�X&����y�v@\�Ç��8}&ƌ���_
Z'�B�k\ZB/&ޥ�:�*R�I�˨������#��$P�e�u�aܧ�_;1��>C�\����e�Y�G�ʍ��e��C<�O<�ݜ�Wf(�,�o� �Ŋ��.]Q��=z��R�g�khԧ���a%��ԀyV_��\�hW���]��[�.�Kp"��s�z)@�ώ�(�0�!�g�@�Uw�c������J�͌7RU���i�'�1��ܲ�Fgѿ���(^hߨ��z�L�b�47�;��(��8@{��G��Z��CK	�q�7���M<�G�UI��O�6&ј=�CRO�n��3�'�����W���*�L�q�}�\;�~�� ���ڿ�;�7\�a��D_�X�ng1^:�J��1�Kk�S�-�%{+Rul. �Ċ��ؠy-{�\�9����T�[N�7���B� �_�˓����^_C���6#�J��K�W�Fb�;|�n_q�񦅤�=<t���{���8�-a��B�- ����"���� �=�6�*���-�7R7�ۛo��I���!�W[LP����5��}�F�k�˒1�V��$�����;�l.���3�KFV(*���V"�W%mCn�AH?�R�3�}�:��s��VT@D�~���c��]_������3���Y��ڬZE�Ё�ږ:J�Ns`2��XWԘ^Z6e�3����-�4M�',%�9���-�&k�Y��,4�y��ӣ֭|��17��Ac� Z���b��Ϳ�4��J/���O/L�mfJlPqv�ޥ�N�ɷ+uU�B�޲ �>A޷���fHߘ�XK�,��1���G�ݟBX}��}�/��z���i������<𡼰���T;!{ncl˨�9QO�����x�<��L&$mb��1$2���U^�9cZ/g�o�ꎉp��V��7��؏��;>�[PpK�e1}�n(�1QT�%�|�J9,�S����J��pov�i��1��'uv>��ab��G%r����C�ob^Ȟ��V�n=�5Ԏ#蟾�`qW�0*�/���P ��c�Du�k�BFd��ě\dk���>�b9�K�+�z4o
`U�-��&tyUr-s��W}�܊+�N�
�K�9��w
 ^�A{y�(���Nb����b���a�/Uðk)�*�����^��u?zI>E��P���� ����u���q���:"��º2;�������(%B"`��~��t��OI�����enF�g��ёl���d�Z��3ѱpymn���=�ܙa� 
ܵT�q鯋�T�L��)shli��.)�7EC�1ж����wK&I�>3NA`�{�� Ԥv8$�׿X��\�7��띦4��]%v�pTtT(���a��J.�TȚ@���\%2C�a����� �k�|w.����pgդ�P��=�"^�p����QXW_���.Xg�ɔ\�uL�(C��բdլ,2t�������SoO�+�� 0��ٽ�S�h�⩇h��������[1m4j{�㘧'xVJv(k�M [�ډ;^���E��(���U{<9	X������mL�B�h��p����}��uI�A@�V~I¦�d�����X#}`<4�"ʢ�-:v]�hd�P���OF֙2/c�e�ݠC~f�'[��'f�ԃ�3�/��+�#�?�����-���<��*h��n�x�C�At�m7�2*��_kJ��ܤ)3AʟeĚo�>�b�\bPK@���g��L�'��$|�\j��[���I=��n�P��]U'0��z�K܏�w�����,�^���=^e���b��
p�;�!]���ڪiFsБ4��x;:f�W$l�IZM�Q��������wbU��b�}� ���[�c�c�<cn��f�m�
,L2q��]�p�`F��~��f�C?�H��/�:Dyc^6K�$lҲ^F�qe�}�jռ��L��4�{ɨ��#�@���q����у��C���l`3���Η�?�|�n�g��N����X���d#��>����s�������>��電m�&�.���^^��H���-��>E���_ʘu����	�ڵ5��|��@l[�:���m�4���s��Y�<�OKR��ؗy�{gV�;�z�q�*�/��kR^m��NO+�l1�Ǚ��S�l�'�eېВ1`�KK��d�T΃8��א�˻�L�P��/�AS�3���"$#�r�+t�&�ʰ&i��f�"%7Z�� hn�]�V����l�P�,/�N�'z3R	���\ÌqFq�>H�*�xz�� P�R�i՘k���C��[\5���\I�H�f��Rm<֦�d/U�̣�Zu��
���d����!�桝jz���9/��8<(�%_(�Y�GO�_{��-yr��E@W] ̘_C�m�=�o��X:2��%I��tD�3�����,;jQN,N52{��*�e��QM#[rG�T�����9����Cמ����O�um.9XL��~��lzv�BJ��&Dx�̠�%G�aY�8z�ݴ�˴LՊЭ�[���K��Saa���Xp��T}����/������0A?o<�E;�+'�)�o筬�{W�6�5:�bA(�-|B�6 �Ė\E��z����	�7�9���	|z�*L�ځ��0@3#�?d�����.v҈T����O��~�_��㹙��)!���<��"�$�Xwy�h� �Cm'�8�3�׏��Ϗ�R���%k�6�U������� X�*_Z����*/�QV����M(+m)i�C�=-�1{������D��M�Y)O�&Р�����Ԣ���=c�!�!jⴽ%������5=-���TPes{xr:ɀ���&0���l�yѷu��@�Z�(�{��q'L�G�ߔ�j�6�3ch ��@��pN�j�A���G'��,/g_�a��\���`&$7�饺h���>��<�f��X�7��& �qMࡧ䳬U]*F�v'����A���[��z�?"R;Sg�j=FL�[n��}�9bY`��0<��;�M[1�p�h4�����HgO��))���4cI�b���5x6'$��e8�5�,*4�ޜ�;� {�m���婣F*U��_5k>B�	.K�:�������1��j.o�Vn�-��,ݿ�S�4���k��_�Q�
�5C�r�9?��C��T3��o��t�����JpF�pp�6�h) �J���h�r	�>�{�+3��
:3�K���^�?;Ic�6M�iÂ�P��& ؄�KF����b=�N��M�\��s�L@��=�ح��:Q��^��	���Y��jz��e�@�\�Z�+��"�u�ު0+�o�wG�ńMn�d��J�C�`&�a��s�khG[wО38��rpK�nG'�$t�{�U��٭�ڍ� �ֿ��Za��n&�]�-ul�F"skM�ےR� Q!z���fRV�`��Cʿ}4���@0��9|��l��s|;���ږ;;WBYB�&hX���\��_�����X��ln�/
���^F:�&f]%휄�H4����ɞp��A��Z��W��n�c��]n�l���\i���s�!��z��.��
_����(R����3���=S$�o)�l�|��r���Vf�F����v*r3>�YZhX9����**���xn4/#\U�I�Lԡ���y�w�3�DO�nߓ��5��q7� �(�,�m$f�Մe_W�,_J!�wE`3�@3�8��ScdM��l�r��閼<%(7�;�A��n��ܐwg�)�.��iT.{!*f�4��W��>�����x��o�Ǻ;�?M�-0�V4���AK��;�#�Gd!��j�.�H����C�nA8V�=%|y���h��k��#�L�H��>���&O��I����~̃DyR�P��`�Ў�ǌ� ~~�Ӡ�cǱC#�B	��G����	@��NK�ݾu��L;���J��X_�k�1seTYN�#M�ÒC�/S��/Vۃ!�Qǻuq���zv��hW#D��^�����~^��Ә:�63M6DL��!&T��ɓ����[�O��t$ 0Kt�#wt{u�(�*��T��r����v]��c>�hX��2�+�֌`�7���K�HlS��U�Uw�fs�*�c���MG,���8�'��8q !�#�j6�8H��U}T���K�?�z����1��`�d��Fq!�i����\� J@a'{$��D͂�Z6E��y��B?]��S�E���3k��App���D꩜�
fzZp[i*,��h�ԧ�"����.�:�&A�)��󈶶����k�$����
�!g��.m�EKϒ����f�q����qTYi"Q�ĩ��V����%`�n�#�8�dY��T�$�U�'sЫTf���?�kWg�+ҿ�NԺ����tM-ws��}ɖy�~`�9of��W��]˛�h;>sN��ުW�n��N�gzJ�l�)�SW]� y�L��1#�.��F#ޘ�d��ބ�g
`��=c��8jo߂�Q�b�� �r~4��L����p�5a�i�U]\��~w����w�]��D�s�pd�?v�ݥŝ�ʙ�sm�? ����;��3�$�ϮN���}܂�d��w�|�P��{���t�|mV����`)>���A� �s�Tֲ�>�q��	�+�1L`������bM�Z	�z���UL��ڝ�E��c��F��QEJ8�����U�F�B�} ��p�@y�i���)ɰL]�%�tpEܣU�Ҝ����η1"�#�i�
��Q���#�����'���K��W�z��i�����2^�?����,,��v?�Mu�8r�]��m���,B��d����C ��M#R��R�PCZ.�-}���{(��K��mH$bN�v �f&6A�����n�*\�5m�L����uQ!f��6��#��>+����(����52�.�<��8V�py;Qg��+��9��o?�f���Cd=T���ǲ �p�AL	�����6�^`.U��+?��0K�x�s`�{TbeF�R�+)���{��_{X�:6��~n)
=C�L����ex��We��D�W����Q�Ҡ4�ݐ&�|D��Q�O��h^1��7��^������}��P�3d�����Ŗ���~�a'�b�'���.=K!dJa�y��Ǔ(�mhV|X�K����Ј����_�]��|r�6�m���ۋ}t��F��3b�\����0-��xS�n��<�M\f='��� �KǠ��~ԏ.���%i�W5&�Ӗ�C�<X�8�6r(�ĉ�J��*f������,��p8�\_�$j{`@�Ls��k8_�)\�~!03�6�*_bT%n�f��r�9�	���� �4��ܡƥ�N�� �#��"a�'V��P�<�m�D��yp�[)y&N'^�*�Mb


��3����W&��埤<���D�<�	�l!	����y؜����u��9M� ��S�E[������G"^v��ߊ��Q�:H|uBٰ�	*_�nO�`#�T�P�E��No�LeVZI�ͻ�R�_BɥH����%Cj�E��΅��n�s�4s ޢEX�A9�n��⬲��4��Wp���O�һ#�M'�� �>p��CV؉�����՗T�5p���
��C���������6-s%G���E�`"z���.��/vˌ�d8w��G":y�1A2жS!�N�ٺ��,�:�=�*������U�Q?)��k�è_��9c`y�}��_��u�o����`��/�hh�i���>>vg�u.�W��\�cO뗟��+IM������*����gq�AZ�^5�K*V�&4_Ǔ��R�r�r �b�(��mX�i�do=�`��;;�ʌ�w��id�qbi�]�>֒{�v�����x���l������6z�R.��`'��Ht1y6?"$�x��� �[X؞kW�~�Sg3Y�`D���_��0�T~˯=����I�Izj4���Q�9�n�Vl������@�sM��q�D^�J*��ۃI��h�vC�X�@yL��0G�*Kؕ��ju~�J�҅)����_��k./s﹵��ƍ�-���~��}�����և$����q�*ޘ�K��^V.$��O\�׀ዾ����4\;�J�/p/&[U��y�O�C|����$��1�oD��U��
��h���]!��۶J�x��*?��`�j8�y� )\P>��٪MC�@&_��L4�@�g� 3O|�(���E!�������c#璒�j�,�)��X|~$�#dZ�4�]XC�
'R:�y�k����,���<TL7�����
��m�qhi��Ui]8F*�_����$��
4����m���-7��Y.'���G5�����*���w6kd��'���'ο��k�G �uqX�o�C�8�Pj���:�V8�piz�9�ě&{�^�&)�X�f����)#��^� )���k>+5��ty�9�<�z��QK��֐܉��X��d�ݩ��S_|͉/�np��Y=��;��_�}�A]@����"񷵴@�E�_�ͺ��|/#ݿ��B�麡��iSt9��S�L}�w��YZ#eE)����C�8�n��y6�%y0.#͉w�l�H4.a�Z!��5�\D�;NuFN�=s�0k��X�Y�`���90�� ?��)��hrs5F=��0�?!Ơ��'��&�����1
�A����y��� %�.�:��χ�� �j푍��llܲ��eCɛ`��Nr��ZW!U�61L�����$ú\��"�V�n�Yy�a�S��TQHreZ�!����r�*�q7�R��ˤ�r�����Gt�9�s��Ι8T���njG����������jHb�Ԁ�1��35i��P�T�����瘝��ry4U7� ؤ�i]��P	���_��&��Y��l<r����TOLȼRJ9�����|��o\�HTG�DelS]��N��UZw�/�]f8i�6s�{3��KJr�L�x$B�!��궴7`�p��%#2��w	*���&H����o�>��M^�r�Vٵ��	����z�o&���x�c|�q1�׭C�a���.(?�\3�Yв�����Z��T���c��+f��bC���
���9����/��bR�y-��Q��=X�}s��rt�?�uHи�L�Cd9�vʊ�:��Kz���
��`3��DL�ӻa�k�"Xo�9"Fyx$8��.G�C��G����;�j:"C��ȗ0_�O>7))lO(P� ե�ڒ�.�ц���Itp����`��9�iD�"h�̬y��Q>|���^��Q��0��e�f���
JB󽞪2�6l׫A���+�OX=\�1V�4��`�ݚ�g���8��:�j9v��N�ʢ}�OI/	e*Ʌ����ڽK1��a��誮6>����Z��nmv��v���Û�؃�\Ի�e���ە��]��b�<ؗS�C�10 �˿Q��D[���ءe�X�0D5B��d�=��򽼢�C������V�c�KXG?�K����xoتu����T�8^Qj�.n/(�^.L1�~q�Y7I�Si^:I]|����;�Æ.ro��81���yV����3�R Z�r'SKA!n�5�|'���=Г6kp�ƅN�q��K`l��g�d�m�?���8ǁ�|b�|�}l1^m��"�*�e%��w"���/�>�N񊮑¾���]p�^�wW#��a@,��_
<��0���<���Md@Ph���(U��1}M[�%/·m(�o�1�M�X螹}Xu|[]�&�\�{S���F��Nf�6}ǀ5�rX�&yһv�ӓ�$T��-�]��~�N��!V��񐵅����g�΀H[]'M>��Fes�T��[���|�NC�ef~Z(���:��K�Ti�#�Q�049�r_�M�&��~�H��NpG��4h�i�:2���^oZ�����qߖ�D��4;CL(�*�U�4Phx%��y��j�!��H���.9mIk�Ǹ��f���XZ	j2ƣw�C5�����F�c�/|Yp��}��Be��0>�+f��+�M��
	_�ѭ�9�@d����&h��$�B�q~O��S�V���8�r�X�Ѣ�_e+ƊM��;��}X��b�� ���c��b ��ď炑����}�gⵅ2���I�6���W`��_�E�(�rU�'9?��q`y�Jg+	�>&G9,�#{j5 �`{���ۻx�f|��QqҞ	/!w��mzӵl����|�����%pe��"͒>��G�Y�{j�z۽�K$~�����xO!Ɉ�g�g>�S�6^X�|�*�c�^�5%82P|j�7k��Y-��I�����s�|�7��v
�Pg���
fjT���c#�S2�L~���� ����恣�a�aurnB�#ŏ,M|eKؤ�� U]x�:-�?K1mG�،�i�Ch7�y�4%Ku�~GZ���@�M��	*SCO��_|>�p�����|��j�ů
���l��jpz�g��Nx��Pېp�)t&5��l��p9�����5<\'m<>/��(rF�3���|r��z��h�6����>��Db��R�ps�HD�Y��ʡ"��p�rad}�M����a���#Xv��3��б����P��B�"2QΖs㲴i�?���k����=��ELBYaw�`�5�@��?�yT�{��ODQ���\�} �^��/��wk�:]W�(ߥ�������[#��g�0��O
#Y7������b��j�ήZ(zȁ5�����#�_��j����6���!���R3p���8n���S�k�,st��R����얪(�b#�Q�sq�f=ʹ�JR�lkw���d}?ʓ��-�<���[A
�ʊXu�����	��[���6�=7]�ZaM��7�`k�3���ٿ�C�͘4����Ǖ���S�^�����^���hP�����i�݈����:1šPsP�,W^�r��lb��- ���K�=�+�fK�FN����?��L�}ۖ�'�����̔=�@��z�l����B>���� ��,��`d!�.蠿G�sL��&K�(~H�����ڛa�ڽ���0�%m"��h��u�x��V��k��P(���?T�0l�Y2�΁&ikS/�'�n����� :R�Ux{��+�α�e��[�G�pӒ璈	!���(h�:��/�l������Z�F�%rSi�*�Ҫ>��|�*Wں쳽`3N��5�� �s�*4�j���Kg��r�y(�t�'��b��}AL��,���;Ԓ������bФ��e�gj�� V�&` ��+�y��}Ƙt������5W�0e�y){vO���â��M��a�����4{E�-��<�8��2�:#������|�t�N�Ė����&.�Ů�LY(�S�=K�J����,(�ـ������tb�f��.������������"ܕ���� ��OG=X8i;�/�X�s�;V���x&�+I��R�$�8A�|x(я�E�\8����u��Bin����_��N2v%C`WT<o��!�*�4�+}�Ǯ��в���y�~�]�����η'�S��=q$o�B�������P��%6ԙ� !�j��<���(�!����b�gܨd���]!,f'�Aw�cIZ $�Bi��ވ>0����ڥ/�PE��*����#���o�s�ӟ���ve�^L�xLv�A��V�C�u5ẅ́�f���U_������@�)ռ��;�CxC?Lh-p*�'0{�l{�y�sg}��%cc�5�Z�r����,&x��n �u�ͧ�wC�m�&"�z6�rr�t�:6���B��#�Ղ�A�z�-��>��cA�2I���kδ��+�2],����Έ�+K��
����C�MKA���,���90#;f���SΎ�������ǧ��.���r9N�?~�u���G̥%�" 5r���P�Υ�3��Ǝ��iӸ�Fy2=q>�(L�^C<�1��k�������#�{�����c�K�����d+�_�X_�ڽ	�{�_��	~��Pl��Rb���s���<�uv���N��q�m���_��	�5�FY��YC<m�!��9�[c�kLKƯ�X��WH�xN��6V�����?5��b,j�����c��Jt����|�pLy�\�f�bP��p�h{�"O"ߚ��%�����r�;�
O�������e�[��K�d�m*��>Y$���[��@a���Y&��L���f��'d��,�&d��_q*��;H�`��4��Rm�5n�h� ��-�lp4Kc�0s`,qF�Nnmİ��C���|��3jN)��x�31v:�"����y]�X2�։���F�Sy�E� vXBr���}l�q��zf2��Ѱ��>�H��>��.Xb��V��]�j��J�ˊ/3�:����5�	4�a>c�>y�����3�\��(�k���Zi�0]c��)�"��TG�����>�nS9�i$7.|D����>����N���4}������سA��.^073�e-��A�2=ǹ���a�.�J5ֺ4�Ht��7hD���䎨��<+�W�Sw�+ǉ8B9a�P������px46h�����t�D�z���t�� Q��Қ(R�6ZSMۑ��q���/�MPW<��궎	�P<��HHHP�S�:���NN���x^aX�e�U=���xXe^��Q֓��9���YeR�D撾U�\1/�ou;�Z�$��]ܤH��pV$����$�Q`����
﬏�2�Y�s�ŋHt)�jt!���\I�g� 2�6�"!J7�F��>!�t ���z��ܜ�3��1<�����mD:��*(cWk.z�o��Χ��A�a��|B���3�=pR���T7p�K%�q�
R��yT�R�jy����S��V��o�QU �J�v����w���/}S:$��2Y ���1oV�����9�N�V�����R�4��`�����Jk:~���t�-ǘØ������O���Q�)y�,��_Df=�0��Œqϒ�cb��E�S�-!��`lˑ�חb��~sm}Z�0m����qw)����{��20�2�2C8i�I�Z���@Ճ����%��BMvZ}�9��I�4O�Ǽ����O�/�p�a'����U+4+ݵ����'�Iغ��[��yr���ݶZwus���
����X5ʍ/կ�WG���ٝ|m\��z��?^��h��K�I�)-͛*E�B�������'�ձ�2��� ~,�?F|ta ��uD��(__EI'�Ә/��v�H�P��Kc�,�5���KDs�8�N&gd�ڤT�G_�	���~iݦ�Ҿ�nd�:��qr(�]�C;��)	*����u������q
���o��G�����Q��O�O���l�{n_|��&�{���k���
2�� Ͱ�:/pe˔�<Pw(�){�Y���L/��{�ݎ˚������̸([�sߥ���[�لQ/p�n"Ek�.�Wl������jP`���������*�;g�r��8L�o��vB��r�guPU�:sC+�ہ������hҘ���"�������U���Ez�uU}�gĲp")��IԪ�RE�B���z���j�O7�� �
^��W����?�_Zh��+ y9scٵ�kN�;��FX�Z87�0��6η���������$�+z aʤ.��u�NwD�&@
����\�9��9�/��j;�[&IMtd�H�m"��m�n*-�?�~���ם��|/����Xix���f�vrųY�:�z����v%�k���6����,�|��KV5���]_@��0�:�8�_%�ְ���&�#��H��d�n�����o�o��-�#{y�'l�"ڷ]J/o|�m�K|����ܴ*O ��T�N���"樽���:禲N�à;��k_*������d�S�l������;~4�kU��0�`+�Ý�� ������_�% :�l�^�JٖU��z������MY��p  TE[� \Q�ꅀ�Z~nb���To��7��UBG��N��x�Ys���Љa�M���Q�d�6��f�
�/4A�VE&FT0�D(?��X�檾������k��S7P�����R����B������|�}5�x�ž��q�Q�Nb&��v!��"x*��l�틧�qFkC���G� � ��\<S��^�n%@G����v��\sy��N�{��d��k }4K����ٙC��i�L$�Ć��\����Bu��K0.����Cօ��:��BH�JO����SV�i�<�V�0*�D$���!q�M���]����E�oν8�g�r!6<��e�}�G�s������Fmt����r.�V��Ceb3W��<Pq�E����T�&�[<����j��ub_b_�*��w=hquqEW���*�rpV9'�SNT=Sf�ъBI��k;�6���>����^2*���g��(��:[zP��rG�mO?9�Isv۠��*�P����I���9��x��X�Ȧu�v�X^ӱq�TM6^�qT�_�%�b$��o���[͈`? �Tkd,��n�L�O\m3y�CM��!g?��߹���<�ު&l~��"��UJ���M�P�.l��\8h�Y������Sߣ��R�;x" :�Oq�����l�
�?3C�ֻl���������za�,:}�HTx��/Ja���!��
ШkD?{A��cLTѠy�R�'
�j����K'N����<��۶�A
���|�����g��� ��G�8��)ԛ��8(��	��:����B���~��=�cb�6���³�eG$�s�T����% R������i_�O�;3c3�+O*q�w��a/%���������*`�hq���z��R`�q�ʭ��IMa���艭=J�A؆�j�s,E"ec�x����
F���Xݴ<���t��c�W���F}fsk4�4�F��C7�b6�K>7>�ʮw����{0W�xLVHu��pכX]s�r������n���+5K�wI���8������T�V6��ヱ��\���?0;��o��;��˄�4hF��n�=/����W �VL<������0��*�^Z]]C�i��H�C��L��{k��b��j�.������0�����;o��e�^�T��%�?�L���E���3���O�}ȑ��޸��.3QZ����}[dj�
[�^K��ݟ�f����7LK���*8��̣���q�i�Ң-�O7w֫�}>���
B���\�_!^H4^Bm$���޴)s܉=�}n�^s�Z��V!� 8;ŏ�ԡK�^��ތ �F�c�ZN�P�!C`����o)@�/)���]���pIC�B�}_������h0�����^$�i�%�`�o��
��\xr.�p Q�w!>�*rCܰ��-�U��b9�{EC�����2���u�tZul��Wl9��M/���z�Y�ƪ���=뎕��[��.�ƥRՔ~3�@��ɕ�r��ף�w}Z���3m?��jM��|�]�i5����Pc�74j8
���k�F%]��3�S�%1���b��I��p��(1$�߉���V*s��)��;RI7d^��A�	�� L��B}"1~�c}�i	��Fߞ'�K�b�=U,f�?1+��"�A�u!k�Ѐ�����}?|����˫Ӻ�˓��5�8 g%P�`?��������(rls�&&����1���}�BPX��Hz�~�ր�%G:Ye$�F��<�j���: (�$@1|��6[&'n���z�,L�<? �M�A�4�� ���(0�F�����IN���7�Ƃ����M*i(R|��k�����ע�gH�e�5�r�;~�����h[�)K�-��!��?����^8_�������u6m��p��yHW�+�U ��$�����ӂ9X� |�j�@��
o��E�
�>\bڶЋ����۸�-Tᢪ�y��φ�i��~��0[$�ȧT���ed�9��e�2�~{(*}@3 T��b����n�`��V��J��R�:���q�]����0����T�O0H*G��X����D�q�Gt��C�:���늖V����.$c�,�� �*�-��>�E	��y�tM�̦Gm��F�\� ��u�������V��%l�#�Չ���[s#��m�n�$F�,��7�6��Jxoy΁���&,���ۏ.d/�d����f"�
oMϵU��|h��#�=�ܔ�s��vjp���T� �ih>�Q��M�a.(\�$�����m��m���Q�v5�mX1Da�J��F�3�rԝk�+���8*�~s�����	5�{��G6�W��7��a��'�V��!�~�u���v��f��>�G����� ��*�z���t ���VX��� a��9��au��k�m��,mѫ��hv):@.<4�v���߀��y��{ގ����*B^LAs���G,T}��������܊`��U����'��46>��J]�����8��\�i�%P85V�o��Ǵ��pvr�c�cT�Y�����Ie�	�KI'kW��7T�8�K;����|�<�k��Q`H��O��j!��~t��'�v�(�R]�mH#�ļ�y���'�X��	 ҍ]�y��G4��'P�!��	����L�xcO�ON�ACO��	�@�9�����	X�
ժ�d/�B�UF��$3��mY
�Zhy�yO5�Ձu����ym��/�)#�ӵøH��WSٻO���e�F��W��E�+��i�)3��R��U2E��	�ᡉ�����)'�������w����5�-{�2ʂ�U��ֲ�-�F��b�E�Q�s��X�CS�4jF�gz��JF�S�q(�<��{�&�}_���W� �M�Y&��Sآ�
K^(X;[.�~|'M>U�y����C��ǐ��O�E)�\\#HlV�?��
F-�	�8FG�G��y��l瀣�|�>W�I�7EX�_ƕ��l,����AC1��b�����3>T���юFiS�yc� ���UȧY]��/$�*�w��_�h�����n�fE$��r�����3�I�A��~؇C��/���v'g� 	'+3w�,����wI�2@�l�D΍>?��m�%ódV��7 ~3G���p߃c�Q!����u'z{!"�Y�������c!s�[�@B�l��!H3c��O���^���Aռ�Z&�Ƌ��{dn��b�0�<��<�9	�gzܛ�`�����=�`��g�����{d8��i�i�L��e��8i����k݆�4��uK�L/A�7]ϥ��i����A������E����5��M�0����*�!����Zh�x�H�i%��F���r��]Las����(�7�GhP%��d�q�{�W�R��t�%`���l�c��2�<��$.�d�AR���,>'ָ!8�(cn^��eF��>F��Qߡʨ+����EU�Z������}�J{��e����ce%�,��S�b��MoJ:êrw����_��>o9��Q>�B��u[a)�)k�Pa�=�ǵ���e%ޯ���Lw˳ר�1$۩�B���M��݀�gK���(ښ�2~|^6��EL()2���ſ�[R�U�	+3:�[僕����8k�LH����ʚ��������eL�8����4^ʘ(&-��텨ȹŘ�y#��9=&���n����#�>�NQvm��^L�S��)�F����t}�A�7-~�3,yt����"�K���j��z�ڗ.ӟ@33Q?�� �|3g�{��m���8R�G��~���y/�����?q%p{��l����a~�<�P����\T�K��}��!�����T9����/6���]�EmX̖`B#5��~�Y�ր���K���_����ot��<ό����Z^�ܚR�x���EB$ѧ�'�X]��SWU�٣��Cb(6�d�+�?���A�ԡh�Q�s�7/t�@�W�>Cw�����l8�e	�\(��0D|�U'O�z���c�ɨ����(�jY�)z�����Ai�T&�x�����9X� ��eD�k�dϰcG��H�8�L�y�˳�c8�Mn8��b�e�ke]agї!���J^M'��].saۊJ�]s�G�t�+6^o�<�������x��&���٣��|����x�����U�%�t�@�%5�|o&�69]BKZ g�T�Q*k���ȓ���pT}_��z&+��s|�0րH �������R�س�������P�.u�6\덖�?��'w`��6�C;51+�*�|cvd�1bA�Bs��P�h�yⶾ���C\K�g��Z\g�T]���\m<�N���++jg�Y5t��E6����Q�G�/����x	���{qI����b�����,��c0ƯAjH���rT#�_�SN|�p���"$�{�'���<x�Q�2�]x:��gun&��*4��Y�X^�e25V���Qϯ.,<f�LM��S"���mE���@�a~�q3LY2s��\�<�*Y<�d6l|ϱ���toK��¾d��ҩ�@��b��d�ӎ@�~|+ٌ�z�����+Nc�-�P���d^tM�E3���#\nNj��F!�Y�gc�k���5%��m��_]|��A q���k�֥�c�8Z���KP�!�D&&��@L�x�*XO���ޭ!>��M�j����jU���E�T�P�ڰ<ʐ$y*{<�nQ�>(Ru�m��!ў71��5D3$�Wt��$���d��v͑ˍ�}uX@���J� }kv�y�$:��UdvU��PyR
��d0M��6L6�f���'z�Um˯��Ȣe��.O}��u��������k�B�4��n/���{�ƵߒP!a�O�<"N�q��p�
�b�����
��k�خ9XV�F��k�(@� �]v�BI	r���u�ґ�s�{`iQ���1��^І��p�)�HQ��٬ʕ�};By��Uܞ�������y)��W���L]=����#��h��wj�t/��'��I7�܊�G�ظŇ�Hk�#�9ڇy�(�<YX2�b��ɭ�G鳩�*��h$��Uy�d�I>�b�`��<gC�߉����w�>YVm˱���Q,{x�Y4��!��kڊ���Y��U%޺:��"��v@WE#oP���a���gc?��.Ȟ!t�-"
P���5�?��K���3~>=ҵ�;�;�����C�� _�]�z�FG��G��!.���U��T�D���ba�����������s3���e�P�����D��j'�=�!Zy����3x΄A��ꋈ
���xQ{����HAq�b�b~ќ�g�V�\�Bl�剱C30���C��	�pA{��c8��u����њ�pF�h~��]��LĝH���f��6k�N�ԕ��E��J��E�=�ТyQնm{1%3UT^�
j��s�����ج�o1A���ճ#q���*Bp>�(�*�P�w-|�.ѐԥ�q,��1���@ޭ���!,:2�S�V��0^7�}Ԕ. ���-�iK�|-�t!���s�V1~��*�r����E����Q�}B���`
l�-A�U��aO�}����Am�!�����!sa�C�ke�eD��TQZ$�����Ge��G��1������,�׃�'����T�q���(�f�;��mҵ+�wD�B��n��E8n�g�n�(�a�JI��v�$	�CQ�sNi��V�Odl^�^5���u�t(��bbڗ��T�,$�(�q��f�v�h��'"&�t���Q�<k���i��.�R>�,�r��E�0�bAa!�QJ���b�7t�@�um"Fg��OC�$ڿ�U'�A�!0�����;��GxJ:���t�A�Yu��~��k���7?�Oo�.��PS�|�K,v��_�p�@��Fx_*�����<Ֆ<�]��b��
\����Iv�58@�zrU/��od���&��q�H�C�'ϸwy)?c�h�+����.��]��ْݚa|F A	1����ӡ��B��Efk�`�w++�x*W����ia�:�T�E�(h��Ϲv�!(�Z9S�\�
�@�Cx��<��؟7RJ����5O���ؘcz ��֙5f��Y����W���_Nڮ��'����0)�i��l硟f��cH�I�*Dl����c*3N)�5�z������
�r){�ON��;$<A����a���*u����
�H�R������_ �UBgp�Q��Bȯ����e@T80vW�E��#c5(��#1�f�et�`���b�F����S�������Nֺ>W3UYݍ<]ߴ���K��.�ʃ��i�,d�<素Xx���x�Ut�A�Uz$�`��Ѫ%7��{j\����8����b��g-Tf�g������H�s%���s��K��'��j�U���[�{3MK�
z��*�I�����2�[��n��8O�Q�t��6�x���H]8R|D%�RyV2s�'v�Š���vO��.!fU&T�MAJ!U��k�c�P0Sp�$�����:A؁���|�@�9=�b��T�e�r�H��%�����fsQ����:���k�<YC^]ͥU���MhS%�q�H�<����Ǆ�!S���	~��V�$xZe��J�Oq��Xq�����VƳNu��YZg�R�����}>ÂY�GO�?�FNk��h��ѷ;�O�ņ��m��	JȎo2ɣқȉuZ<FC�80G�̂��>9�-� `�"_f��f���8��ܱ�Y�-61�t�J������p�i�Bcz �޳��������պ���ME#��m�5�� ��,��SW��hZ��g��ʲ���p�H�R�/�~T�]��ך����dK����~�.U�����J�>�E����3d�z�"y����IƜ�XJN�*6�B�������*�w#�q'��Ȟ�P�c^X�	#B�a�p��D�l+�D�z����k�7�/�^��e�C�靰�/�>�w~:'�t`��*��V�Q�1��9��D䅜G�kZ0�?�2Rp��3��sy$�3EY��A<�",/sN��ō@���B�N�fDR#1�L��#���f��/���YaͲ�tl=Y�x�21�+����#I��Zw��_?Έ-q+k3ܗ�{<�Y�*�z��1���I���B
������J(�@�cT@�!���Ɖ����X�.��%s\e-���gy�׷�R����yawG�"�����`E���3�`���SN<�Dٙ� �H�ԨAN0������R�@aYQ彖S��m`Au�#\�9��������h��l�7�q5Q���争7y$�V��I�Z��;����Au�[�U|C4*��[B�tF9��_�3��z2�^��J�����!x]�(�����pwj����'H{{X��C3�cX�|CEDO�S�
��5�|����s��W7�t�����e�3ǝ��p�C�O-<lV^@��GN,�p��Յ�2�XH�����
�>��`t*麵������U&�>�Ot�f�ތ̢�~�<ܯ���[�'�+~���(�e5���:�Ħ��2^A��e�����<$�5)'¹K,��̧�#KTO�-(&��s>!Z�\���˴e>�d?�1�۪�������6&�J�3Wz�a3�ս�f��"�3��"[_n��"�q���А����#��m��m����K������3�n-�;��n���0��eZI�21!v��'�kB��𨩐��Bm���1`fG?&'������+D$�� ����{���J.)ɗ�\�r�M�h RM�J0�]8�R�bh�^!��4 LT�t���`��*ؚ��|���_܀��c�T�tCt�"����r����N�ۧ��^ ��)��'R�"��c�.�<#�[�J�{n�>^��V��P���BY2)��}�q�k3�$��#��P�@���O��m���2��y�%�ݸ�B*{��B�1P	�??�e]�^JZG�ߡ<B��Cw�*o��Y�nW9�aR#���y]�� `�6B[��BN��6"M*S.L�~w�P�l�]^$�p�#�f�!�oʃ0���d�q��ʭ���F4��96�v�>�F�
�]Vo�����e�c�D(4x��O�y��"�%���6?�_ド�@��3r{z@0���)N�8o��8lp#����&��1�v�� X8#r}���f��n9K�as(%=�f|�V��ݡE���eCξu�S,���5&yR6�����a�
�U7�B�����!J�1�3�{ta�kN]��_M�;�G�u�����UVPhҹ��REΆxu�;Q����MPn�l"4l�4��)骞|���$��P���l`P]\ӚcFLgKY���S�2�ER�O��l�[��D����~/�$�gT]��8�/�`A�A�>A�w�(���n���`����J�(:�����Zl�82������g�\Ej�x�9O>���U��n�I���݁������kCeO�n	K
��V!��ga@����G�-/�^��9�)���M�W�d��'r�]�����	�T����?�{$1Mm7q+b�R��G��N�qR�R|�?��a3
���{�u�����LҒ�;8�ǅ0�L�����t��(5�)|p����YC@A�� ���aqi��5-B���F U��)�:���|�yM�P	�J>�iΩ�Rˮ�R�m�,������\B�ￄj�.�r^u�����By.�\�cҷ�hD���+~ �9x�3F]��]��z�i�˹4˘e�0�IbAV�N�|�wJԹU'p1s�S�����rj0��쟒�Q��}��
�J��a#,L���'+��7�v
��a;V�Pt�|��?еֵ�XXd^ʩ���9<�|�t�&i���fC��w����kkU��e�G&��q�iq L���_��jB����=&�E��;�
�˱�g��#qSfNb��\�ꝱ���i�}9����v���W��%m[��oD� ���a;x�w�X�������.�9�F�l����;�!O�Ҙ�HD���?V�E��#ln%vxƻ��cA3��չ��m8��Q��p���n�il2�����<�Bd�����U��K��fjZ��Ӳ������Č�y�s�����J+����l![P*
������[ �nw�%&���g�{Z�4U��2�j��ɤ�.�ũ�rBkS�L�a�7�i1��9� 3J���`QQ�x�i�Ҭ��K�@	.�bt�I�����/��>��C�Oc>d7~.g~��V�*�y�����
�Zw��^��P�	 �;@u�,��}�"�W��^<�2�Da�Є�)�@v����s����Xc������3��3v�-�<B��L������!V.�y�f���E��ٗ��[܈x�[�n/�v��#��䗈�q܅��ҁ�l�NN�h Kid#:�C��yo�F��i^��d"�0�J�]=׮���� !
j�W�D�!n��C�]ۗۜo#ۮ�pb��O6Z(�Q}���: �Ҽ����E��WA`���2�=MpBF�
ě7�r`�	`��E���	�9Z��?)G�E��đPXFߎ���5B5So����|��C�;��<��)�܅(]���8  *LZt�f���L�PIWl�瞬PY�ũ �r�J6�L�0t�FK�*�i�3Vܐ����\"u������an�9$�20�I�Uq��;]e�S�	ܚ�E�˵���V���%�2�@�L!�PC����-P1��4:���؊Z����}�r�S�Շ_&�<����h�lL�j]��-���~�EhV�̳,"ʋ-)WU�D���:ҟ�,�đF�ҟ#��=zY��h�!ĩO��tÿH�h$�BxE�����/��ߚj���-DF���	*���O(�f�h*M�j����Zۜ�S�S.���
�VS�E�s�qS�듩��m����i��\=�������з��s�s;�Xg2o��3L"���̙>��Sε���	Gs�@��0��a��cG<��;|<�A��G�<7H��1Q�p���_�e
��֘��/³:�S6����Q������q��_�6؛������7^������"!�+j&���?w$��u�* O���31�%���!"�������S�C%��K��q�z����Q�wy_	~��yJ�yM֎s1
??���#>�Doh������ Tg��#�r,�X	�vN�ivS�柔�{Q�0�k�gw�3�F�8XoY��F}'�;7�+���ǫ��v�*i+�z�?���!��6��n�h�c�hD�3��Z�@��5�J��i6���wv{F0۩5H��6d]P�������iu�H����<}�-�[ڜ�w� �k��简Hs���u��Y��9]�
L"�>'��dV��d���gF�n�]�X ��m�����Ƀ� ��Fl�Dq�r�
t�D,9 �*�d�>�O��&�y������o�ǜd�8U͜��+�Z)z�0߽��'���e��Vd�����O�\��q�I�7��|�'#�/n��i�X)�"lly\��7dVn�����g��j��f ����D#H٭�kKʁ�fU�m����Q���}qJ�������~�KjB*��mg�u��2�-���q!�I����(�� �`T�=,|�h!(��)dcj/^���0b����

�1�����A�����G���©ɱ}![69d�`����}�]Ĺq�S��=�̯R฼'�ϲ�M,��k �a�@���+>�c���p�MP)mc*�9N�q��Z����F���y>��J45�5_ґJ���?�s��~�B<Em��F��6����K��@����~��K���y3&��������v1yk�0v�Gs��ߑA��O	�Trr�b�Ԫ*�IB:d����r�'_���y�sGQ/k{%8k=oR?����u��i`H�4���Ԁ�_�c�6H�mX�[a��`!qa�iBq�C���k�tǬ��3L���G�+�ߒ�z `�T�I�į�0O�0{~Wק[�� �����'}%�~��Q�������Ʋ��Fj�q�Q�Gp�����Ox��Q����r�p�5�(*[(ct �f�̙�Y�}�w[ D��r�]���-�M�@�	�-���e���Tԁ��b
����b�w�t�!-��o�%�c�˰b���A�l��������!V8u9a�zd���8�{*h��>�l.2P^lT�"�*Փ��(��hy<����f��d�A}�5kQ���..� ]�7S��I���e4���/{�Ld�ʲJ_��f�068Ԝ��
t��1����`�E"S�ٶ$�ؕ�]$�!��)�ɟ�ڟѻA��I��Q�����U���3��"�J����$KTT�E���M�+��[F(C�؋��-m�"�3(��D܆��C���c�}z�3��\H�rj�w��7� Yܱ0���� �"ӟ��W�H��e{ubCvj�����%��i��/�Ƙ(�d��q=8Z�l( �F"�{%a��`�y��!��������r7�?Ħ��P���j�&��~/Ѧ�=���O&1�h�����~x�
Z3��j݈�-�E�/Q��2������qc�I[���=W/DX���T��]4 �^����v4+� ���x����kj��K1s�"�6	��,�����ipl��l��߄;|a�L���%�>��O�MIPA��~��n
Kc?��j�ŝ�n���I��������Y�{��wqPQ�_��,��x'$���F���\D�Ԍ�u5pݻ���]d>�6`a�RJ�E2'+���G:H�|e����'��7h߀a�ZaT�f�pϏ^�O�������1EW�zFD<Z�2����S��L����c%�A�+�o�̂6��6�	�)T�"�IsF��	yuێ��{kȋ�$��z�e��ɳh��)拻��I9��,�\u¶נr{��ϵ��*SkV.*�[�k��%v�SZ���<.C;4�����^iA��]�����RP�6;Ⱶ������@���-�<�v��{����	�q�F<�f�i��,�}�4?�.�	д��bEFh=>S��5X�y�(��&� nty�(|=�Qy�:,������iC0jL[!:��8�&�kĪ�v�9o���?"��Isē�������:v	��hO����V�@%�������3�a���0ϣ���R]��Y2�7ǾiP0��&5� 0��	����[6�7Q߮D��(���5�2f��"P+	��!� �|j}���aD��eU|E�/zs��)����e�ә@ƾ/�F����� �DW�Ҏ�@�vН(,l�r�	8	�=�|�H_�M���c8��������i��������cX0xm�N�̃>�+��|%�E����@�� x$�`~�_1�o��T�B���xo�V���-K6��6��`⡋�-rh��4�S�6��@�{d^G3N�V�I"R�x�������A���E���B��k���v�6^AU�>�J���\kTZ��4<y�&��5�Q�G�C'NÍ(�;d;��G�����.2hn�uvJ�/	7ԛ�����]����{H�rq:(�h�nNo���d.9��1N�p�f�g���ÁT38��z���ÉӪ�#��C��uHJ�$�h<�ef	��L����Vv+�)����%���Q��� ����{k	��%��ax����Lwg�inN�9M��U<o���73�O��}���Ʋ�:I�,�yu��D�����x@��։���f��+簈L��p7�bo�w�\AT�]�w�lʨaX�jS�8���Y7�����,3����˲��6��ȶ8�����尣�k����S�$#����tò�.��;�ז>p���]��z뾱�=������oi��}!V+���A�l)���.g���H�;!X���]Iw�*�E��LyR C˶mg���_��ͤ���T&esf��H����|L\�Z��z���Ic�`�`n԰Y����7@�k�a����!ZuX-	���;�g{����J_ ��o����(|N���a�1�� �ڤ��Wp{�^8J����6��gw�^�2���2�zap����,8 k��?���K�M�rj9ή�BU���#�t�!�s�6�&T��3��p���| �﯁��w��Ԇ~��H۠��I/���,�8�N�f�á����������W�4�ㄿ?G�v����/�����߬����6����{.>�Oq5�Hz �������Í&�t�̶�T$ot�Ԩ3'*�������S�M"���Hm���-��@���5"J%�M��e��i�1V;݊8�����@
O��;0*�(�Ѣ�����M��SM���K�|`93<	J$�Y|X ��4�m�NRP�Tr��T8L �y�b!�}=9�^�R\����٣�`/�4��m���]� ��U�?��>˪�l;�2Oj��(�Q5���,��$�	��ᒈ?��8�w�7w�B��u69��tk�z��>���,�rP��-�B$ڷ�����K�=F�g����ϑ(��(��>j��e����K�ְ���'_�&5v~�lZۥ8垥� ��o?PhY[��4�[��O	��[�t<������&l4�LK��'E�����(���yX=�d��"x�� ��!)�+�,�c�����ذ:.���\���1�JY1
�g'c� ��HA�.sg�*�]X�Խšֱ�g1hO��NGE$/�?�P{C�ϋo)�-�k�o���{�Qm�_�,'/�^��b_�	Ij��))X�=\�&�����-$rugȺ;4��!J����ci?Z���u3�� W��
 ���@�I�q
B�ήd5�rL%n䏉�և������f��^� +�G%n'�/�x�n��j��9`;�#`��������`���(
�͒B��cowq@�ݫ��"�
��5��f/"pҍ)~��:�:
����6i�PS�Ƥ��z�H1�E�ł ^	�2��xyz
��5����p��H��@�W��t��"O5:�2��TX�b�.�~�v�
�q\E���������{�_��ë���1=]#�������b�X ��z�dv��J���-��U�S���z�o��Q3� ��+m#�L�JH̭	���4]���a��.�1��mQ���aR��}���E4\l��=�\��� r���|�N}(y�H5��W��	>ॠGl�G��K>3v������]*�(�iE�^�$Ws*1\{L�[�[�c�I�iS�@	[-͟gT���0��:q�T���攓�C	��SS,���]GJ� d��_T�����V-6�^#ʥ%��ό����)��zU��;��/I	n�>�~���Tz޾&���2E�n|��ϳdk�T�w���!��0B	~�G���X�~ǅXۉR4	�١��~ߗ.�5䶈#��+j�܊W�K�fo!Z `���L���-�Z*$�DӫOP^���;.�q5�!��{zHDɧ��e�2Q�dfş�焜��x��m�Ӌ�N�4�~K��N(qUD�nW8`�82����b���y=�̉(����GËq���80bNz��E ��I�1cLm�&R�)+UwU\[ǖ0���!��/%|"������8�@�=���%�C�qVN����O�=�t3^f�o�Ե�yK2"F�jQRy����
X�Fl9�@��;���ܽy�t�f�m�m�q#QL�Jj#�?2���"���T�O �N���}%�,��?>�tO��yx�?�8ﳛ�Q�kL�������x�t~t�L�gb	b^�ܫ��n/=�⚚8�^H�x�iT�=∅������Q�v2�&��
c�)ǘhd��u>�i�r�GA�+�G�&S�^S�j�-C�"x�̝���E�Mhk�V��Y�Ţ,��|���[vgN�ȉ��������F�$�Qo�֬����u�y�YI�@�y�1/�s��q�h\�G���~�,�-�"�䡻�ՙv[�o�3�z��On���o����I� 2�k�fdki��`�� �Ynq��e���<�e�请*�^�-��_s��j�N���N�%wq�C#
�$�C0�����R���L&�I�Pc<�w7)��q�X�e�dHٮ� o:i,�@M��v�"�3]�ޕ�[9&����eN��@V���J���.g,n?`._F�M�g��h`^��9���J�9��R���V!h�Q�k"qu�P%\�U8!{�̸�E{�T�ٺގ� ��a�GGڣt:�����T�ElXV	.lK�j��߻:��[���9cߏ�5�Q�x̎�M�Ԃ������jF�V|��Y��a� !�$���2k�n+��Z7gMHFSs�&�u�:����Q
B�(�LS�1JW&�K��n}�
H4F����;&�gу��`�&l��&�5l	̔��)H}U���	�,9�;�������Q?��$�#���`ň~ԭ�M��ߧnK �Xr�5\��Ak2�0FR5�z2�:eԘ��p���$��σm���k�S���̶��D�U�#�
�JR���A7[]N�-��x^�U�+*�o^��N��^�?�86	xE��h�U�(+�G��h2�`O?.)�����Z�?�+�e엦��A�y��O�ӛbq��-0$�Ѓa��D�i ��D�D��nZ��'��m[ܪ��`^X/gZ�4Ii���%�j|_<H?�W���>9,E=���w��R5._������۽S��i�D�;�!���������M��(�(X#�����S�C���nD��o�i��^�����Q�a���L�J␆؂��3����p����մ�I��#��A���Yu�r� �Q5�Ruɝ݋�m���w���V��H��dZ����Nq
�3BC��CB 3S����G���O~��
����Rq�f8nM)� i��d�a�ؒ~f/vA�)P���!����,�s[5de-�Y��尐��H��IYG-�6���V���`���/�gi5�;� ,�<4a����yf:�T޻��� >��o�2��J.�ݙ����@=sMɟ[��VH�CV����=7.U�YxDG���u�B�Z=Ż�:E�Ӌ�ߝ� i
*��HEd��4�M�ڏ��`�{! �[M
2{�5��DZ�!d���*�p�<�u ��� �z�{l�ƨ���8����v`�ı)VΒ^�/��,���x!k&%��&�Ъ*��~�.��Q?�H�m�o�z�h��,3�԰�=�(� ~�k��q^�J���Q���V�i�Ѫ�;�~�s}M��􌚨v�]��]���u��/����M3����z+�hP� ������ѱ	�&tQJFT�a|��p! ����:��߉���A�R���!��8������giG��d{tu��ʳ++�\x�Z�[m��2vrO�^�N��z\��!4h�ս�b1�0㾺s�g6��o���n�� mØ�݋��B���`�֜TyV�(>~�](���_9�/�O5,f��;�{T�x2�J$7�8��ϊ�u���R1I$�sϰ��T3��i3�豑E��Kc�E�9i��=�{��K|`�"�5S����OK��޹�+TS5Q�!=3��v�����l�Kv~�e�F9m�av�wf���c�2a���ls٭PIz�&�g���J�����g�:��©P(�O0��6*�Ꙋ驏��)����[�e�x�[ÑztDM�'<�C���@A����@M�(�L�ƃ�a�	��qY�%J[<�$�ؘZ�Ώ�L_M}�ij�@�ux3���4j�+��32BK�:���
����Թ1�(�!	���j=&X�!7���~�*};pߑ?V����b
	V8��-��i��K
�W%�����岈�q��w��!e���HSU���J��c�{҈�
�K>��@�	径R�Q�GDz�{z�'B��B?{����`�����I���Rc&ͻʪ<���z��)XEa?{�e<�M_k�
��񕙂]�#�z�w����`Ǔ�K��P��D����(�3� �nmUO����KRg�A�jH����G[�����7]�Ҳ�Au�����9�,.}�A���[ ��F�	��g|vb�֠c����^�a�Z��q �y�p�̿��t��?'�3F]�OM�Τ��`��ċ���R�qԈ1~��T"��_���cP^�u��e�/+�sÌ�+�]9
�D�
����%G#E����8qo8`�Lqh�N!�_xm��n%�N9��� vi2�//Hj�c|	.�G�ȑf�;�W؂���\l׹��oq����R� �?5�bH�C�	���-��ܦ���ͷ��'F�@�v�$�I�yI�-}��0_��+���˛{�tr&�q��������{I�T�ko+y��-��z�O��٤ �Ϙ=�Ϥ��\;�^G�X���vcY1<�6F/,��v���'8�ʞ~�Kig������-���4D륊��K֥�%> \.^��	�W|L��U��S�(>�2��Tgo��nl�Ȃ�)2`,5����x:�>���^[#7$�:�~���x�Q�_j+�%El�-E���[��v��H]P�������:Q�oM\�5�R1#�H���A���<}�:^0�n��Ī�4��AP�$����@��{��-o��� {ӭJЎ��P�oT��s����������n�n�%`�Z��	��y����͌W�����"$�tKќ��)��������>���4!�#���t��!�_7�/a�]�hʔ*�M���4Ӂ2͊��Y'SS��O��x1K:xǀY�����o��d��Y˟�9�N@5 1�	ϼa�PA��6�����>�dX��`n�������'X�.ŜP�4�d�LTB*-7��в�Vx{��5yh��N���������f�*���5�Mu#�8��E�Y(�ytW_j�a��s�/ꏼ�;P�ܜ�~f�HѺ�M���˞/9�E��˓��_�s�6�/�q�bp�Ƞ�U	L�	���x��I����t2ES��4r����6�=��m�	�'�	r��A�)�b�`�e������P�v�>����߉Ի������i���I��.�C�&�DG���i�}���{�����+O{p��:Mu���/�d���g�+��[�p���_����)���`nj&p� ���pc���u�%.�K���O�Iݟ/��;�p7�G��>�p����\��JԹ���k�͙B�����~i���_�E�)�w�y��������<�+g���z�?1b(�@m���|��N�.jї��0��eO�O�ҟڈ/]j;lK5�MJ��͆�qT�: ��q�fyI���8��MK'��,�Y�n�jn��F�lʨ(�- �D�s�ಲi�Ey7���0'[�<*�i�������6{M�Bζ/�e+6�%ޙ^-���f�.M���~Wsƭ�p�9e���wN�|ۡK|�[�D�T����������G�5���Óɽ�t8�q��x��i��A�l~6�&s���q���\��d���w�&���E�0߀BkA֢�t��BA7\E%2D	g���F�ٷ��֌�ZymX��(�e��w�,M�+`�6�J$X�T���l�譋U����a%M|F�o�ɼ�&������_\���ضP"���B����Om�M�j���Y��R�ꏪ����$-C�bu��3���pc� POl'��Z�Hq��`{�7�J#s3���l��sk�GB a�vB�Aq\�z�L{X�aP���usqX� 䙌��;Q�D���:;��z����ɟ�K�J�K�8b�Q����|��	T�%[*�+��mHݟ4���5�Y�W��5��c�95%g�Y#�ʞ���O� M��-K�~�N��3�
����ʷ"gT+b�eya{
Ѿ��˺�e�Q'�=�n����`d|B���"���L���'mÎ�c����$��7)$5�5'�F�v��\gw��y߶�
�J�߃g�&O���יh��:c(eP���j�vIm�d��}����@^8��߶=�bC�Bul���i$�"��<�}nT>������t1"���\�4*�ϕ��%��P�q
������gkt�Ɂ�u��'EK}�i�.Qy[��}�Õ��p���A����)������Ϫ|��O 1,�>V	���(V��(�@��ʝ��fl �wv�r�ʯn"§vKFS�1��;-����2�(�x���h�����[�q���o�˭dޞ��q$��Q)����K�w��T�2t��0������YEPڹ{� �Fy{�&�gސҺ�Ս��E$x����A�f�u�p����'8�l�7�~�bS �ڔ��㦔�P��Y[��̺L[},ʊ�$'�x�|_R��xWpg�7
����|&�F���Xw��~c�e	�~1,�O�"gty�f�?&��z��j�p3�Dj�8��2zż\��9	���[����9�T�j��5���FA�J�Q5��h���1�/~UQ	5�e7�	)G�b��$��(���6Sr�ث�|�Z�ŉ=�ķ��Ƚq�[��<z�ѯ��X+}�U���j Qp���4�{C�8;�g��e-n�R�i�+�+��^��E�g�Ee��1��uB��;��9���^Ѷ���yPle27����'�����<'CoCX=�k�v���Å�w��ڌ�&ƹ0�j��Xɢ�����l5��=Ǌ�r?�����l��I����?�SsK�P�Fz�����[D[���Aĉ�Y���V������}xǨ��hI�.��`Ĕ�Ǳ�r^N�� r�M�<������6�g��(?�&�rg�	��פֿ����M$��fIAS!v�$�t3e��!l�N9���l.eQ�D�s�QӋ9��A�6Oc�2sU$�+~�V8�\��?���<=rW�Q-�skm�]b�3҂�e4�E�0�k�r�]��'��p���@�N���i��2T.��&G�:��K���7c��2�w�2 [��wm��9������8|���z�2JFs||�f�ZĈc)�F��ؗ0(D�fl��r���j�zi�} ���E���U����Q�~�ḭ���K�-��j*��ON�0����a�Nx�2�����ƽ�T�gj}1a\�\Y���e���@ ��j	�;6y?Tt�ܑ/ڰ�ma�|���q���W�.�b���L.��2N��@�`���o(vh��w�����7�2�5�� /��ƅ�Z�y/��<��(����`�	A�w��*���iB�C���E3�e�@�]�M�u�<���m��nATLL��A�'Zot����&,����	�؅T̽u�&�h��9j9Ɠ�5ƵX�����%QN�/�܄$}���A/k��}{���CȇR�(���+��k��)�R})\�MU�峳�~��e����w�����䏞��"�x��Qn����b��.��?v�1��k,�C�.D�=��w�w�ze�,�� 8���p�p�%�����d ��#�����A ^FC��=��ћ5����uS�y��z�J��ɥ�M&�_JW"D�R�� ��t{j��CM(�p�J����2yt�ɸm�Kc���u�!�w$>H2��#٭*6i'^֗���~�du-Xc��j�V��������|w6N��(�cwe���YR{�ӳT�ey�hX
/��1>2�n�A�с
���
������+�J�~>k�ц	(�x���{[C�bw�1��������ܱ�qCu տ;:���-��x$u�&p���uQ��$I�x'�`֛���x�{J��9��r�0�eEl��d�YWG�x�u�����{q�ɽ�C,�R"�`,3'�Y��hH��a�Z����}�BI"���s��i��z�+l��{�0��X���Fb�������ҳ tO;����9	�F��v%���6+�W�Z�}��T�m;��"h5�G��_���� �d���sW�)�!��Q�G�@�/Uy9��y�O�,3�N=G�D��m�_�0vz���UvSN�&���vW������^�`���6k}:����u���u��M*5ZL��O�B�&-��07XX�*�wlbUP]z��M�|��=Bܭ�aD�:b����6�֗�kg�ǫ�,��NO@��G�m����h%�8}N����dr�?`��,cX=�L�_v���(Q��y�9��L�uE~4���UnJ�ڭ�A?�܋$�oR�Pǲ ��/T�l�������Ÿx�%
3G̈w��j~�����έɰ�#�>��1��~bD����<�(-��4C��˧Fb��N�E�N�a�FYd �^!z��#���Q���ZS��}>P�ȷ��1��5�C5�֨��(e,��v���k+�<N�������"CFǊ'�?�^�#r�_�%����@���E<�l�oj��77;us^X]��H��B�i��GƂ.���%���f������8v74�k���|#�gd��K����Z��(Ϣ�����ט-!�f����ٝ@F����c^�Z="�;�縝�靺��N��4��e8؊o�G<sAn��0����k�8���fB����j��ӳ�X&�j.&��=
[vTbK@�R�EkwJk�qT��fw��� �<�˪a���k�Cj���)7u����Kʥ�\�QD}��D���K6�}����s��Z$��7��H�,zrv�t6����Mv
���,$�^�Vi�N���)���P/�d�����Ȳ�t��M(`ɒ�ǫH��{.�bfv�F_x��E�k6c�=R�7�ZBNe b3�;C�p#��-�1�e:z��$U�&ES�E����3(M���J�/+b8C�7P[%g˛�x �>N��*��У�gHF0{��5�Oc�#��̃o2�F���C-�����0������s* ݒ�=��k���y����	���ڹ���G�F#�!&����l����X�/c�K�����#�Uē�F��"@UG��|��3j��p� �;���� ��'�����+�1<�8w>]��F,�9���4<a&��i�7���zg&�C��!����X�{QR��N��J�|���  (y��˔��.*e�X���x�"ď���H;uo9�����NaYn�	+�@	 �|�<+�:��^z\(�߅W�н
 H�ldO��xP;�%3A*�+�w0����wo�;�Q�f�x�G��Dë��";mU�F���o�i��O���X3oc�9
y��>�j/,����rU���}0>M@2FAM�r�=��i����n��ͩ�&�8����� d��N��턻�Ĩx��	B���`����F�����T�ޟ=�=��g��łT]�<�ϕ5%N�����μ��ԙ~�x�'����k�Ǣ���<~U� ��D2�`gs�W�z�6�k�:�~�8';j��c�4��.�G;ۜ~Q��m�'�%n�u�S��� }h{>�ۦ0H�G�i�,��������uUR3�Q��,L
|CgPIP�4���!�KM��tݚW���|��'������m�R+��]��$�*5�ϫ:��7�omH�<��6�3��Dy
���ad9O��j�&�Omz�j��m`���ثR��E	`cz�O�O*�;xxJ�ԶXC��V�٥�� 8q��Q���й ��Z�
��v�x�!��Q���=�lŤ$���4�:Z�����'ܩ_F9K��j��d�g�0 bZL^�ĆeCd��A�9{tr�=��p6A�͟�-��Cwv���g�(���1A��!�֑t�*a!�<�/m�a��5�t� 
ȿ��;���6��ʹn��9�nO�N����\wmm5p
���?��ѷ-�Úp�(��U�,'��n�[}h:��'����(�`��0�Zɑ�q��R~�g�6Es��e)ɳzHG��{*���$�y*�K��I��7W��}��¡F&Մ&\����dv�iѿW��r:r4�$J@WT����g���֪<r;��Y�}��a�x�N���U�z�e�W�˅�-o��]��bn����?�W�]�p��*9���/ܯ:�c�yb��J㡎dU!AU�w=˼��и�ݑ�=�KuT���Y}^��J���S8OuN.֕�>��I���z(i�;����`���*�i�GБ����璕\�~(|�jE70tU
����A)}�H�Hfr}��@�X�m�JBʩ��@]��߃<���I�j�u{~*�{G�p
pV��gz��P�vK�]�Eӑ�N�&b��-���O�n$?���t}�L�ײs�w��L�y�^u���r�П�b�΀2J�X�&r�tͷ&m� 0��ܑ�N����`���*,H�Ȁ������t6uB�
��F�K�J��(OK���YVߣMplB
���Yk�(���HRn�3x���8s<�(]��rT�>t
�S98FN-��@�E��)�z��/o��dȘL��k �k\��?w� ��%���l�)�{̓�CfR+�M��B�����t�]��b��	�y���4x'���JӖ犻T��;V���h�{Q�R�u^�BL��
��(F�y���<�@�ן8����N����/��yg2e�����S�HI�܀�fٛ��ɍ7iZ
:Hi�~x���/����R�K=	}bQO����F�a��.f�z|��F0yʰ����~w�ZS��9ʢ�gCu����i���U�kȿ&p�r9���v���Z_@�H�E�2��[ϖU�;��n�8���p/ =K�wAn%�f�����C��]hC����5ɑu�׮^Ŭ�."���@<�^urH, ��������/���Ǽ� �&��K����g���V��!�n�y��#ܳ���E��t��d-$TqD�m���w�� �"Ś `�#�����ѯ����N�����륎��ٯ�`w��ޤ�w��l�Rl��5�u;�:pn�Ot3���"�93�h|D���	��\��쓆\[
����j,�w��+-I�φ�G�ȱ3�Cm����{5�U�s�6{-�]�P�t��뛜�7}*,�}���)�I���qO5C��v�Q�x�ԯ���?����l��@7`���ۚ*���[�ď��n��ɇI��MѰnG"�%����v�{�?�x;HN.������+PI�Tr��v��I���{{��}����.�OF���&��@2؀H�Ea|�3�vr���Ǡ��m^{0D�-��X��0JO 3J�,�aC鶏�<�HJ��e�+��P)�-�3�uw���$�<�/B����؉y�j�&GV|�^_1�7gl8:~U���Y�L����o��4Q�[k�����r��.�#3���w�y٦�P���	�"�>J��.����0Ѯ�ˁʭ�aW�Ga��9`��I�S/6��UŐn�T�H��)�ǂ�N��:���T��o�c����i'�y��Hm}~G��=��L��t#��LNI��E]M�D�na����V�{��+�����^�,��o�{P�<��Y:e-��$��Ow��?���D��	.��SJ�
Q�le$��%�A��k��f0V����07TDx�GN6�;��P�6��ؼ��K��O�p��Yf��Yp&��A�0<�Ŷ!q�å��)�`�b��w^'�����3�w�����Z>g�0�Ŷu���ˑ?��B�MO�o��Wd�����S��bCZG�7�WRmW��;��6�͘��r��<J��H�~�P�h��ԀRv��m(է�����I�6ܰ|!��|>�k�_xqG���|ޚ��oA2�tFR�_���*�ĕ�\�=�d8�ĄӞ�o�k�bV�dɢ_���lF�������H��-ҹ!8�<,�A�����v��P����rI�
��%*�R	�`a�g��:?VU��iMzD}x]`AS��</ c��5��b�8�C��iC���������"���!���iB��O*��:}� ���ܩi�� HX ]��CJ��V`�Ӌ	�e~��㐐w�D�!*"FF���1��߉ޣ5���� ���s̛�����y~Ҷ�_-���3�i.,���!_=d�r*I����J��2�$
��ъ�����ta�2q��EW�ۏ�]e�^��~̻�����Q$�3Zb#|�0���k�����K��vO{v.U��f�J%��d�/��?����n�x��/J�\z>o���/h�>���G���<N9e��~>�E:�FPg.d��4��p�]�m1��z�<QR��Jk�h�M��9ɅzPO'Q�(����;��)h�~�ܴ^iK�ɬ���^�������j�Qy����Ӭ��	����ˮ׽�]b�}�D�{��|�/�����7"�B���#<@�.���B���� �����A�9�>��.��,���0&�Խ8�܄u�@�Wv�"���F��M|VVe`$����S��^KY�����?�?��_�gNXPF�гS�!K�m>��5��c"&�\9��+�A�s���x�f����ו��z��e/Ѥ_�4���9L���e�ⓦ22��_3y%ՕJ�"ה..a4MMK3
,B���.@,�Y���R�m�Z��R��":�)������{�w���q�F�pB��W;	%�<c��������<�M�ڽ߮`a �p�[��ɻ3���@��	��Fp���M�kL|�p�j!��dE&;�~qΚ��}�� ���n�������n]�ޣ��zʐ���úH�o�r�@�7�@m��gH!���Δ�����7"U_lV�҂&�h��Vq|�k��Z�f1��C|CZ�쇃@�A��2���NYz#h�_-��^5]A2g�Z�Y����d��o	,Z���)�?��
O����,�1�Zyŉ��c~�G�ʄ����sA��8����A]�c��\o�B��=Q�]�#�UW�@M�$j#���o2�=���O�Vu��~'����\��Y�EЉ[�K5��=V����˳Br� O�K,Y�\!�U6���4U��F�����q��g�Nʿ���h���o��ɹ_4�b��|�ܑQ��+�\$(�\=�II���5ɓ�^����J�v6��R��yѾz�ߡΰB��"0��[J2"�R(��Y��g���=��9Љk 鳊�.������s�ZOu�����̸������7�MUy�4�O����
�S��p��ܼ�3���~*uff~�'aV}"mE},H!w�S����p3���N��f�c�^�Ow��1�QcbV籈�aT�o|����1��6%�iھ�S"\zd����D�E�����q�~̰m
�����:�4�]N��;Mx�����Dׄb�S$�@�S@F����y�x=P��E�E�H�2��!e��8.6缤�eW��)I�� 5\��k}���xw�t�X̦~=.Y�k�5��-�a\��Y��l~<�� �/��	�\�.�W�H|̕���j��꿴�׹v�>e�1�8�y�>��������ϪH�0EV;����矧y$(j,�}�������?���%~�-g*%X�+_�_�{��h�lH�PBƗE��`he�W1BCL���>U�5AA<˩�p���
�	U�v��v�0F�ޓ�,���T�m�9�Q��)�T7�,��גVR�"a�"t�O*{%���No��&.���:&ًgV���/��%�	ψA�Mȭ��H�X�#z����g(���MV�S��.d].,��ޜ_7{}�ֱ䨓��4;/����\�Pȴ�u�;� i�t����X����G�W7�l�������1�g�̠ç��<l#K�9��4Fxa��@"���xj��s��J�DIɉ�6����i�����1�p�-],��U�t`���#���6��"����*/9i3���=�^%�y�x������L�X�"l�oN^$����:YΗ=I�3_�}�̖�Ϯv�u͐�,9��6��}����ͮ]	hB��E��ⴾ�P*7�|+�\K��n��G�m/b��2��65P�G�q�_CF��e�@dR�'�+r�9�N����z�sQs���
�5U�r6q��2�C\��N��#&��Ip4�,q�A�1#��r�˝���F\;���0^?f|l�O����uls�B�h��Guڿ�o�2h�~��uY�<o�G��,�4�b�d�w�u~�2�����[���|���L R�Nq�Z�	�0�,�	.�~� R�I�UݍX~iDZE(^��������y�hF���K5u����ե�56���B�u��|1W��W-�#�@��.���x
��,\_�j� �x��{�v��D�$-mЁ�G�������=��7�`��k�\�D� Y�|d�?��}ՠC͘�����U2vu^�����T��KH��M���E[�3=������I)��۫��|����� @r0��Et�"V��g$e}��z���QU���7�l#��L������j��v�?���C�ۙ&�o	P���ɼ� ��v���}�&a/�	&w�_��^5F%��b J�e����3�ސ<�tx��8w����#vTk����)���:��fė�B���j��0���?Y���`�g��qHY?�^r%#�8
�%��w�N�FH?[�2[xl?w������h��wN��f�K��w2l�aȎ�4����-�b�����v�x���	E؋�%g�� Z��z>��l~�,@	�Ϙ���<�f�1��J�&
��i�2�����h^g�B���$����v�o��}��|ˉ.S��R0�.D��{zq'��|Ʈ+u����cvS9\�#�h�����~;�ȶ���#,�c��� ��)�%��'�`��9v���~D�i��g���4z/�n�H�hS%���y9Mq��j֞4x�{�z�q͚�(�'��]v��M^oBČh�>Ϛ�*!�m"�CNo`.��4�w�б�˝��N���*?
ظ������ֹT9Ӄu�����c(E���稜�D��gP٬R|ntV@r����偷lv�e��n1\�:���c�D�0"oHo��>���^�3k8YQy�C��i����K�p���"\�l0�z���G���\��?�K�w�rJ"Ld2��d�
n5��y�G��]�`UX
��F�Tf�p	~��҃�$��u�p�d򰮮�0���Ur�Sye��E:i:w�-\O'6܎���i-�/��nX��U����DG?bb�,42)�R��� �6�_h�67ԕ��ofZV�B�f�9�;�Q�Ċ$�Ax����t#"�GtE�<'�n���w�Wr�}iEK��jl�-B2������?�Z���Jh��{�$���g��B� >@��rh/E�Xz������I����"�W_[�?ԏ��zk}K�g�t��+6Y���ȁϤ��a&�vS�K���5
��"s��5<�`�Љ�������+jˤj�:l��U�&���?5��c%�|I��h�I�	lOŐ'\7,mj��������:��" �o�x��g<���L�oU0���'���L/�Qx�E�e<��'w��D����La[�oOQ�9�A%���A�z{��S���z:)�%�h.]�l��'�Y��j��5D�@���)*^i��&�z�8��z�����9�.��1��2��_~e"^���_@���v�PCSh�`Eܧh�,�y�43<w��<��!TkV�y���*r� ����^;5�dQP�<�V�t�M�M�%X�]&PP&�Q"@�@ۯ�b���N	��6`�h��(��y�+���	9%K��<�@�O�zC������+���|q}=��g)����qg�t�}�Տ���}�qt�8fyA�e�
aV�FA�AӢG(���o�-��'z}��.AQS�S|�:EBNe1�?�A�=Jm����S�)L������\�-z�=���gu���#��ΛK���Y���R�o��P%)��6���a��xmȶ����]����>0��q�"�(�Jg5D\�U���xE%�".�;�+ڸ}4�}�)t����@�����%oY��b�|�D5������pΛۙ)�yCa�E����Cn�~=���g�_͵�=@������W�:��X�§<2�} �
8����Ui�Բ��_z�[ʀ5����<t�oN����{\�H�T&�ּvV͎�[lQˇd") ��L�ފ%��%U��*kS��8���+�.]���Yiњ����Yû;p��Tw<���������"��İ	μPO�TM��{��w�(��MqR�b~�Eł'�]�����3�L�8|��J} 3U�c/�04C����1H?`���z��r������C�5����G*�c����^� %2�Hn�]"���9�͈:{�������T�������g�ru!̦�P��Ӯ����P���nh+����@0G�<v�`�n�oM��̣��VG�ш�r�#�v�A��Z��Wj�v�}�k�4Z;({��0�i�h�������mU'��_83	}���T�[)�g��L>�����
-�$)���S�LG<P���'��O�)Hʀ��:uH�y��ꎩ�����**�%Gs��X��<a��7G0J�#�� ���oR��%{�?����߂v����lcJǒ<��=]9lg�Q�Ta�?�J������G��R5;�¤	S��{��y@����\o�`�3�*���Sۧ�����q}��]PT�&���6�%?��x�͕��(�S(0��c�L�
������������tgL>B��;C���:�wi�R�8��Cll+�,1cN�&�2�6�˱�H?��|R�qYcuE���E�\��R������]H��#M����j�I0������V�9ы�`rY:<�.�!�PUH� D�z�� ҜOAә4s� ��&��A�/�g���N# �S�?�i���c9xC[�->!-�<��G)zY��!�	������o�MD������'j9'K?�����$��onp}�Hy�5�C�\�u�6���B7_�
h��
>^�p}�JS�pt�G�շ���P2z�U8���Pҝ�@�A��B�~�y/D��B�^�֊��/�������˹�c�F�&��'��13�p����fA�#}�EM�E�~`4A���}�7��N0d>�Y>L[G"6K�S^+�����1������;��LH�fd�|��^��Z�_V����e�Z�o5]�������K�b��~�I�g���sѤ*\gy������r ބ���B�������$Ph)	7��?���x1���h��G���Nr����Y8C�=Yo��B)���Lhp%2��}?F��, ��zOn�d��*�6�8�BMm�o^e��݂��\����be!��芙��lB����144���O���@E�(�z�Q��ă�M,(^�&��K�R����W�&;o���A�,�N[�(�'C�B���0Eb��$o
���
�j~*h"�uG����)��sf N��^�J/�k��|�I �9��6
�X��F~��5 h�W��WRk��8��zDWTw�}kM�<;��*����9���60MZmD��đ�U����b#��[�
�i��01�Æ��q���qh�l����r�#��"�U紸�@Ӥ�JۡU�M;��Gw��J�}p6h��l*�l�y���k5b˨j�ڂ���x���f��{��7�r[��U��d�������a\>ԛ�)0���f�d4���S�;e䟁T�-�����ʪ�F=�B��k�.��7�ȶ�5[׫����I4Ӽuڍ������{�G��g��:����+9����؛_�:����l��4)����=����E����VV+IW���j�<�>,�P�?��F�j8��a��"��n�~���	dJ�o��]��K;��:�MX���wPɈ!D��_��/�S�w/f|n�����]y�{���Q}��v6x���cf���#��v�c��؅�"d�`P[�U�dj��Sk��WS�r{a�.�>�e��O�;ɘ��y�8��	���祣&�GE����� V��h	P��_ѳ���~�XS̼��S�t�n�ԁ�bcL�����eн���;�i>w��POR0�XS�$��HE�p,��<H�+n��}^�w�'6Qx�K���^i�;x�4Nұ0���us�.:���/o�N�%��̣H�#�R� �=ڬs����e�+�~����ӂy����ո�aԴ��2�W�5��7���|��l���Pg����y�(͸jZ��$V5F@���b�]�>V��H'���$B���y?�cTu�]e��a,�S29� �ӛϴ
X��z������hh�X2u�VziZ��i����t�t�/_�QE穲��L/DJ��6>�@.;\��l��~��KQ_ꏘu��@��/���c��G�}��t{�c^8H��Π��=���QDd\C�i�A�)F�Ͽ^�ݏTt��7�ږ^0�O���͛Wg�9�8��)�&u�M�p��k�<Z�F��%jf�к��~"��*� ��"���6��Xi=v>����>�.�ǫ����vl0�����.�����-���(b+<��h `��c����Ec�q�bۙO�I�*q$�i���\�x���I�յO�2��V� r/a�%f��BŞk%v�� ΞRVr+~��G�$����i����l[�Xu���e�!s�)�ND�F�f�[����Sy�sudN���$���3l��C���-g#��v}%�ǵ��f�\�h�������@B$�FL����:��;dߕ�8f�[�Wq�O�|.�鑱9�e)һ��W�?�n����.�^�{d�l��i��8�\�d��b�9�ç�|,���O�Mr÷w�����m�����Mgr��%����K��
''�b�!9���^�\}�B-&�N���aLg�G���1�`�E-9;0����V3)lrXz��I��L(�L�.٪V�Bs�}�|�\�K�~�}�ވi��4kɪ��;�։��)u��¹�q��,�^������ڨC�b��"@4!&���=~>�zg���hW�-Jj_�#=�]��#�CF;�����\к��J ��gjT�@?(O)D��� �ȷ�'�S�t9�O��V'��#,Ʈ��u�0jJ�h�`Ė�L���o����"goe��͏$G�d][�iL�Y�8����߶/�{�$i8��x'ߤ�$�hr��i��׳��>w�ul�N$�t�.G&���;73��T��a�'D5�h����~(y�h�UNI�MR�8�s�%�F'*��V�^��};�i(�(���|4ɯ�Џ���Nʪ�1V�ۜѕ�EU��|Gg�&�f��GT�v^�uQz"l�`C�S��nǘNa5 P@w� �kA1��Æ��u����0Xr\%��{��e�qr;-�R�=whm�^�`>�<���K
�N��ڤ&֍1��|�7f!�f�Y�� pѱ�;�Z�,�b�J�g��f#�9saܼD������~ܮ�!���^[�Q�/frC�Mq�0��Dx�!)�×@;')�۵��mD���d��ۓ��%��^��/�D�!k�v%?(������!�.jB%��һB5a����L��k>��� l�-�Y�ok�;'����FO3!�n\��r���z����_�q�J*:.��̢MP����Juq�b,x�񛓶�l�R}��E���t�viʲ�Cڸ�w�Y�����[�C9�ˮQ��HB��r'��(˱�Nxf4�y����������I����+\)H��D�1� ,,��lM��9"oיsW�B��A�/��/���L���Ѷ�����7O���=:SRs/�gb���L�k�� �\�0<��N}u&�,�c��l$���	�I��>�{��s�i�G�s����##?�&]`�v��s��v�y�n��M�Э��ea�a��d�9 ��U��e��c�mj�D���j.Q�{<ύ5���r67H{i:s i1Std7�����R��j���A��Ab?
�vGm����#ƞgf�~\����K_W��M����
�`8;�X�6���2�Y䟮� �2w����]-�f�k��2�h[�z�}E�$q>\�V`Ȃ��g�~�r�kVn#@J�� }���2��#>�i��c��N���B�|~/����KH0)�1��/'wW~���OmG&#fw�D�QɁj�r�z�*�҄�x�����)��r��B�(���l�e�騖�7�T����ecygg2滤��9����tDe�2��8L��΀��?-�Db@���:#�-���I��J	P�%�l���=�"����]�j�����'`�t��JzM�*��3�j��[���n��+ �D��C�����p�|Q�`��C����������i|�9����>�FSxE��6�,�jѹ��Pi#�:�����a��(43��b�uз����N1�Z��J�ނ����P�dV-V��O@:���j'_�6����|��F�ƝƂ��C�^�ߧ%�gT�T!`��j������W���lG��? u�?F.$��z3@�~Ƕڟ��o��.J��2WV���֖3�Ι�6��]�dw��{���z������c���Uc5-}�ъ���ti �07��x�3�Vk���v>����*�%��F�	oA]٬
$�|�^�7��SU��{,���c�4!�ڴL��`��z�����H8=��n��1H$�����ʔ��-������4�O`i4_7���E��#y��%�wV�_�l�bEn�� ��xh�w#�h3)BX�m�u��Ǎ+J�m�A�jĦ�D4˷5P�Z�2=�%��P��Bz�֘��>�;C�_@`�&T���{�5��{�ED&�E���ȈUB��S�ٽ�f�+tL
�|7o��b6-7���O�*w҈�^:�����X�i�����(�"�Rμ+P+��w��w!am���E	�*ڪ`�C�]Ǻ$}��~I� ���!�o���ӷDk�fԿ���*��F۪"�7��o��E�!�&�z��'}��^�s�,P*�� �!qB�d�n��v꒨dB� 8�'Z����Li�i��D�AԮ�ht[#��'���ނ���NO�F����STP�?�	�-���Bt\5Yz������4$��:OU#���0�L	�"ƺ���gZLU�I����ʫy���w4(��bf/Ti>S�	��N>:�j�ݧ�o��3x�0��c�����IO�l�> �z��U\d�x�zw�d�٨F�
 K�z�F��V48�P%�l�+�ˊ����j�+.Sz)��I������Ř;���T�U˪qR^'�,h�?�����K&�\�q����
��6ջ�a�f�wD4�

9o�A���+"S��4]���ypP��n$÷�?���#�� �,�S�F�x�Ct@#�	�v�XU�{��oLZ�(3WVH�#�<vX's&7OPP��f�er��U��8�睯5��y���w�-f<
۝35�D�4M}��r)�2d?��#Ve7�����ώ>��j��l|/�X͏�Yw�.˞?�UԦ����g�zQ���~9�Ӟ'����\�2�8>5�>��KS��i���YH�m���U��II��-��r��	)Ԉz�[��Q=�LϦc/�ӗs��O�~}�K�r�d��oF�ېZ�:B�B|D ��}��9�^��K�U0NN�0S������{�o!h:��17���l��
�eN�j�s� �9��	n�G�E$˴ZY�4筝��9��J���0��ƘAӃo1��AK�յ3[�Օu�/�~]�%����{�����&e���}"�)�U��O�1�����:B9?���e��;is�����a\�~�`��,Íms���Fn?<o�1[��a���S���R���cR�������RG�������V�s� �mI�tX�� �e��IPr��H�-�����'�����7�F>�1,umu���rUoe\���f5JR=�0�)ҁ�ݤ=���}�YH_C%|+-���6�}wx1��
����_)I��]RPx�8V�U�7��J���_�7�~��/�ͫ�5~� ߰>eeԊ���(�ƻᠶ�9ez�P���	a��Igr:�/s!caJ��=��16�j\��E��1-���h�\��֌�Z�l��w��tI@a�C�E`_�Rʪ�|�Ʒ(>��@��,Tъ�����zG�)"��զ@Ձ�v�y]��ޫ��=��
s0��b���d���k��ݣ�^S��a�th/}��������R�V����k�|�5���ɗlczLmI[����r�J�	�_�in-�7�F���\o�
#�:��k] '�1G���pH����S�奁6 eJ|�u���
����WW*�):��1�ߔ��=������� d��37E����ϓ8Kt��V�V�-W�A֞b��Q��攁(nծ�3֝ټ�^'�����Ps�o���S�8On@�@���CJj������l�&"!Q"���Rpg�F��)͆вsw�����Ҍ����,+p*�t���m���K�Τ���aRn��*��`�TK�������;p������w���+}'&G�I�z�]��	���mX{|>$��^
 8�ʴ����
�,�$ڲ��D��~��m��q�Ui�V3��*z,
l�/�\�ѡ�)�`��9(� ��'6��[�Ej7y��>��%|M�(����^ꃕ�<�IL-�.�̗u��-�fqK
�����T�ّ|��d�1���	|-�������A^����6�ߠ�B�j?��ۆOb�l]��R��]�>���P?�l-� �)����������0�f�/Ve��b�}U���d�;�3f�>
��9ԡ�͌#/�ww$�_�f�%��$s�&�.R�k�:m:�����m����)�sX��1\�s�W�F+>��~YO * >�V �k�YB���	���j��h�&�lF�)�3�FS�~�K��M��\&o�B�ԥ�l�"nE���џDo���>͘Z�Jiٌk�BS��捐.�N[lV��Ҿ��!Gˣ�Š*C�lIh�*\4b �.0��>O0�c�\X�G��WO�c�3S�I!r���}���?�%ر���kr���Qo��8���H�ψ:��F"0�C|#K���2�R��%-�Ca��*�@\�Rc�{������h}�@ �8�O+��#�cn�|U��LO�@��Y�gp�Q��K��om�J� 廯x� T"Y���"��eNռy���9�*>D/L���N�N�/{�M�J��(`K[���7�z��˱_v �ߣ�=G�[���=�B��)�\֕��(6�.�jIz9~	�*��@���0@Q�l�ܾǷ ��W|o'$&����
�_��D>P�B���d����Z�A��JFXԵR�l�� ?,�;Ԉ&Pې֚��3$S�:�d�E�
�S�m0�V��G� �0S�
~ވ�#���z����-�S�u�Jo�ʬ���a���;PT��W�D� �d���O���v�.ρ��!��xd[+�Դz��4�`(����D 6����"�N���ݩ����3@�O~� �⤴�zW�����H�j=��B�����^�a�U�[U���y%��l�:�� @_V��!IF�@�]/M�б�d	��V��� ��������jzm(�
�u�1#��Q��ۀ�\��a�"ׂ�x|�u�r�V]��8�~A����ɑ�z�>m�(:K#P�hx�#U Y$��E2��>n1O����(����U����D�)�e�2���!�O�����䑝���^�O��F�&�/��5g�MQ�\h{�-b� ��-�N x`*�1������c�ԫ;���	���M�/ [2���\�#����Zj���|W�Z3���P�����{-r	UŨ^���TH�h[.ET�E�Q���,�M��-٪2���+�poP[v�JjJn5Ыζ��n`�c5�����$������n4�>����t�zpӀ���(�+�T��-J�j�4|0��9��H��D�A>v����Y=�:[L{����T�DZƁE�7�e��}yJ��õ��]m	��������\"��E��]�1*�ײG��Mo�E�x���L����]�5�=�mߍ���S��%{������ͅs�Gܫ��W(�S��:�W��4ɴ3`����>lU2?Ы�	h
�m���@`'^��������Ir�RB��{}Ӛ�D��U5��&9�f����5ZU�� ŋ2�a���wmL��W�\��_,+h�U�.���(��$ki�#G��\�ЛK���Ԁ�]����>��MFx�o�4�����ln��+���o=��Ʃ�����H�����D#{��f�[[��*	�R�j��Y�ÎFz��i��	y���.z�'�\�By�EF[�cV@��
A����>7���T_'�6\Y0�E�S�n=SEA\��u�[	��_����{�Qh��>�V���������^�h�m+�i��`;�� +$,��_t
��)m�<�`97~�pē��Ak�QȻ�����]`����B�9���9������9��T�]V9يb�b����o�J(��m��Y��0�� �{Wq�����8��/ډM�r�:r���D_ �d���B��0D��u;�g%���S���|`�3���%$f~�GE��_/� ��( D+'��,X�'K�� M<B�<��/~�2�{XD�*3unK���
@�x�?��	�Đ^s!�(W�ګ;��d���#!��ZsX��� ��C�����Q�މg�������b��G!��Ӵ��W�u4M�}�,o-u���LW�r�qIgċ�8��P��z�����K�>��H�.��9�XL97Ȑ���o'θT/S�A��X�a�
Lc�Ca����6<0�W T���ZuEG��AX��e���). ]�%$jRm)~��þy �H:��4l�q�rfՁ?��~��+�{���q |&0��W��,�������4�tTk@�͆���˴�eyM��K<DL_,F9QL"�9��M-��8{�mU��=��������1�q�}�F�uū��[��^��C������:�6�O��Qz�n��lQ� ����s2W���m�%
���\�@��9�D��G��(o�Sy� B>A�}������_���R�R�u���0��xz�H� ��)$�m�67�<�pvw� ���EtS�~��s������PB{]ayQ&zd5� �_I���r��!��w���T֝VHo���
�Y�3=�J
�G�[@����#dn�<$�81��(���	s� ��P8�機G�N�K�T}���wAM����ldL�#$+���t��ˠ���X�]+]�B�4�ܘOO<�����H}+�D���0��xO�r��,��xJ��>��Y�XU�6��/S�#_�3�+�p���*O����G�����5��� t(�LҰp��!��ݻxz;��9i�y��s��N�Et���1̗XUN�m�6v����e)�|`�t��2=^�2��]x�a=C��i3g�py�J��-��w2y�������I�8�ۏ�|�[���vuw4��ܾ��q�r/퉐�dM�!���w�y�Ծ��A`�ZCJ�B(�\��]�`��&�3ϝ}<�?#�^�"������vUjm}O���PMժ����6\Ej�C~�)���J�F��|��M~c�ou��Qo�e�)�a%6w���|G���8{���`�*��~"X�:k��+ӱ��9<�ge��h&~���H+��+C?�N>�~)���g��#>�p��"����O&�	;3�ۄw�ƎJ/���6h<?�-�-���<�w���K�M���V"ºd��k^B(1�Q���k|L��A�|t{�G�p;Y� T2� �>�m،�1���;z'��Y`I�n�_���v����\�t����=i!�Tz�0Ĵ�(����q�GgʒF2�w�@��H��$�fc�_�W�J�Hu�A��MC�	G�	n}č���|E��p"ot
?��"aF�E!m�[oZ�l��򖀡���u+ۄ4(�E�W8��E=7��]q�t�&?���qV�=	$C�*�i=M��2���'%Ԕ��b��uj�}���vBV&���*�&�;���0�5�oA� -f/8n� @��u�r0�T^;��A�� c����L�^�Z�Рa�
{�$�<l(�.�E\�(uL[�N�<�1Ԉ�yp�J�8�M:�G�kM��DmS�/z�Q����͈w���K?��^�)=��"ry��B����q���)ףV/^9y������nRX��-�B}�A�7�3��G�V'ة�9��X�#b��4��eC��yT��M�|J��|�7�c�]߫�!o����o9[?��K�")T���a��W9�D��3�P2��`=	8�"��fx�?h���I�H�I��+PTH�fk��g�� E�+M���>q�ڎ��//��7͋\�.�E���e؟���d/�2�<P0�cά��ٮ Gt�	�w[%>��o�Y+*���a`�E{B�Vm:T�gݝE:��_�n�a�8|��77KBjs�NY���r��_X��t��L5�"���_�	���!\9�!��yt6cf������S�2�L%b	S���\b?��J!�S͔Ľ�}-����k_�Q�L�.����D�nFU�\yI�@������%�����K��C�4��<�%UB��%�fn���WQ|~ [�����~B
@&|DЬ�M�R�TfEV��tX%8�&<��R��r	��S:���|�Ug���3Q\�hؗ��e�(�i��^�p
�V��3����Q$�N��JT����J�|"ġ顾�0<"C+��y���AG��a�8��2*A��-�E���
�ZAuc�	55��X�h�������1�	`��,R&���	���M^sԧ
�X���y�l<���[l��/����+e�hF��;o���}q��@.��u�!�����AH)�.�!�@��cG*��9%����@܈��g�����x�1S��]��=mk(���b ���p��jI���Ō��/X�;ͤ9��&�8p~{�0 \�,�ДIf���gU�%f�F�J�\���^��hX`�C�������Uq�zR��X�6i܄n{xN
�P+c�*�L����&!�4�5Ű=U�~�a�$��ng�׽�8�M[�7ܹ���`r�2�IϦ��p	.2��*9�B����x�$����'�d>�%�`\|G�:LZbh�0Es�<��q���P�鄨�����H�?e7aF!��x�*�A�rY���p?�:F&�e
�ؕ�fϘ22:�Q�]��ˬFC���)�yR�J���>'�U�D���D3AtJ���8�w����<�c7�K����XU���/��Q �G�v|���r\�P�FG=�Ć2�K&���ĩ��)�=�lz�9�L��]O�[��s΅���J�6�i�U���t%5��^^�Z�4q�/��s|N��Ϯ%Y7���i�;Ղ6�j�:�:�؂�o�m=�����q�Y��Y�Y���xfcI�,c8�f����xg�-xgrvǑ�Zi��6��,K�1�ҁ�y�����OiH`Q�"�ʇ�)���L��d��,�H��?Ď��<*p��v��+�\IN�ᡨ�ndd(�� +�,W�	�nV6��M�(���c�!��z	B꒹��c�X8�b�Xc�zU�`����	܄xi�n��0��>Q�nс��m��#��z�ty�6���k�	��m�:aJ��'CL�A��0� ۓ�Wޫ6�Ρo��k:�X>�PA;�ձ`W�-U̢��A�eX�@��ȑ�j(��[�/"l��{Qu��E���WS�^���B��:6�}��]�;�d
R�i���l�7m!Fɡ�Js�eʕ璳���^.��թ�)K)l%��z�����e퀸�~,yn�xR1����|��q�����mN�
���_���
�L���~�����-�	6iV [�i����n#���5�G�aU����p�\����)��hm�c%�T�bߓ��Y�x��Sxn��*�t*Ň<�V�2�/��0��G��>4�EU, ���9rY��Y_<��N�1yH��(;�x�X�l��<o�A��a�fm{2d�����ܜ�A��~�����v�Cۋmku�5�/X���-@Lh�ԯGA���uT�9t�X��>֕՘�]Gu�8��V���,^�<W?�.��yu����j�ҫ��|N��"��)��&����.�c���p�(�X|ҵכ[���=�<����"���fJ�UQ��#�#�2C��Z�]N�·�����mi&�|5$Eԟw���j�"�ǁ���G>4f�)�Ƞ�uאa�Yb���_k��j�o�m&U�ZE@�@���t��`%�(��#�贗8�8�\$oX�3y�E]J����0������eߺ��JV�1�*8�ˊ��[�*Gj�n�?^��+�<\}+�騸 ]�����������c��*��5B���5,z#�ȷ�0��&B�s+�s3K�?Χ�7��c�&�ۏ{�(��h���<�YC��إ����8;���	���b����wp�X@��a�H_�c[f:A�����6��=щ_D���e�m���W��5����a����!��@���o*F&�CX��R\y�8��&eٰipj�EϚ����M=,SB좻OV�6�F�W��.QB���Mc{0���ڵ�M[�"�W�ZpVq�uX�v�2�B��;~Jyҕ�qDB�Ŵ��di��u	����� �J��1*ሼqV�[=�>�ዕ��������{�c��� ��Ѷۅ�B�8C�/��,$�,cD@I�hC,�]��8�ٹ�X�2��4�v(s�1�s������R�{Ȇ��qE�b=w �z��|YP�5�)��0k���t��8�Ḥ�'H?�����T�kP���Ӗ�{��`z*M�O@eI�J�,�'3����Wg��Ve�e��N��^��uG-"$�Y�U-�E�]/�۝5��X�=���A77�6穭��Ŝց~��ht��^��Q*�4��6���n���|�w�Aӣ���h�#�֧��9`�eh$�g^�|�����n\ї�hȄ��(onC�mD;L�J:�u���=uJ�*�]�<f����h��Z���ژ>��R�2ٙ)�:M*?r�PM�r��۱�\��s�$	��=�H�Q�3l3xb���{�dNȂ�Pg�jHS�f�7�x���W\(�6`aQIn�!�׀�K��0i~�]-��SY�Bm7��xϷik�Ϙ��k�����4�}���ӆE���߯&�E��t��9�fˌX4 �/��zh �l
�{�����G�`�A觧:����xGNRY5�W�X�X�K@���0��P����M��ӣJx�����D-A�5��8ŀ9v�K\qe���'^:�M���qY�ӥ�Q�]��= T�-J�/��hu�m�Y8S�ifVa9S��߁�W�Mb �UZ�faz��/��?�61}��`�E�\Yk&�*C���v:���.Wt��!3}�Wsי�V�Z�����ZUf��Lk��&�쬼���ΐٖ]�~���C?���v�#f��T���p;��H�v�����7P���X�9]���ѥ0E����a�.�nS*���l�&w���$a^k�ǾU0�����}�:���-5�E̮n�]��� ���(vK��k��C��7�q:�d^�s�'���Cq�å�E�lR�W)"��ȥQ���*N����_����q��]o�^!Ư�����7��pJp�
#`���&�m"����-
�L�α�8��9�gg��-�������=v'�%J]"�������D��X��qbi����5��$H=�M�ψ��!\�KLg�7㒢�����U���	].��АI��N$,3˕�]� �w����F�sŸj��7./[»D�F����	�w4�)aB��vt45�T%&�c��vc6>���"\�)Yt]v}��x�ë1���z�7�5J�r��x�'#Z�3^O����i�G��d�Ԓ7@6����&��㆟�U���n;츚4��f%2�hk�����q\@{�3H�#��ݝPe?]%�[{�|��d���M��<k[��'�  W�?�l=�}GQ��ѐ�ڂ�_i�c]uSdU����w�*X����6k���[g۞<}:d�J�8}�v��24��p��Uq��9!ɼ� ��cB���#�O0ϱ��2�(�S#	�#����Z�j�R�o���H���"�b���{�R��rMӔv�"&Z����,`J��{aU+C��8�/�s�¢:�QvyX�){!�=�.y��w����b���E�Y��E��]��͖~��Rj�_�����.�惸������vK���Y�\
�	�R� ���u���0�����0�\+4�P��S6��n]r-��l����)�,�$ɚߋ���ys�\.�9 [N��4c����3��O2�a|~mVVp�n��mkl��z, �ǔL�.VCL�ȱ2�	��>b��V�B�G�?S?p� ,򃋷��y
b�|��R�R�.��6;,Du8����A�\��6C�
!�r�K�[x�@Ѻ����]g��&��ɴjr�"�/a�Ҧ1��6�ܬO�����@w��`�y�.��ϭ(F$YA<���&�@q��S��;J��X�E#?�l�F9]O�;/��+�"1���MY`X�k]�/A��M�pT�x�#�y�e�H��W�Y����F�C�E<�|���*�	-7���``]���0$֣�Up��������10���I]������W�å�]1ޕh��{���2��7z��]X�'����u���2G�Y�P�Pྋ] _zX�w�A_�E�y��o���~W���+Ee��'��5k��Ow���52z�ǈI%��t�/Pc��f��{C�4���@]Of	�~�V��O15��FH�j�zvI�&:{��q���e �<�sp��q��a��рw{��W�|��8vP��8WO2F��p{/�Sbf�톻1>35����uM��@��W�C 'J��Axf}+k>:�"�9����7��>�5�#f����Y�%�3Ķ�}iCԚBV�iU��)6����Ӌ ����[�_��eղV���fB2� ���E�c��l��K<rea�#�D"�;B��>q����������ru}��3c,�9}A�\�X+�ع��$UԌ0�ivOď�	����+�E��%S=T���ٖI�G~�����Aޔ�Z�^8i���	,�=���}��8���S��Ո��;�6tҲ��~�w�~�k3���$�\� :�	 5�܇��}�I{�F�t֠�mv�1z���Vf\�<��_."�MA,k4�iG��׆�z�߹$Pz�}xâsC�h��/�F�>�b&��|��0%5���ryp ��bF�v��㺒��jV�'�e�u�����uiI���8�����-B�$��}.��9��HJ\fT�Q��5�1����H������Y�Bڼ�	G�s)I���B#�Vn�nLT��U� �� /���{��B���g���<��R�B�S��̶E�O�>xק���yS��>��A�)��N���z/Ą�J�k����	��@��s9�}@^T@��/�6���~�N���I��.Ӿᴙ܆c,���� ��+�l�Vl��Mt��jss˦������]�]��9Y�I�N�#�����SƳR�F�ۨ���2w�H�jD#8p�wF�:�����Q��Σ̼��3?b=��"ysq$��ʹ5Փ�����O36�4-jV����O�O�&�5��d���� %�h�M\|�R黅���Bn:{M�#$��k�KN ��7w7�BF4��^U7�>�K'F�M�9OA��* ����,ڿaR���B�(a4����\�,��~����ZI�Z��?�xX;*&nV�'?�FHa	�Ɗ�j)G���0�埚�h
+]������ K�&[q�p�|�V���o��G��_��q��BaUa�_^�hw�c�>�pD3�?Mޤ$�c�=Xf@g��ӗ�{�Hu�(3㑋*�uNÍ�a�!����E��F���Z�%�VI���!��l��ы�L&�w�p��W�䃚U��I��fʸ��T����^}�|v30��g���b�3w�ŚCD|;2����"+m9��̊p.�Ŗo?\�\o��;�:Ҵ���~�.��[e���/�X�����G$!�^ғ��F1�ȰN\|U�r�fT�Ҡ�O5��"O[mr����t�4� ������btc�v��-x�"=���}��Q	��W��55�|�Ƭ���UMei
����~ܣ��x�>�4�t��&NEu���5��3~�������3l]Z�K]�~!�oF
Й�\�����_"����7a1��[�|*n2-��C^
\�(�����N��e��YX ��xb�_o��Cn=��ڈi��z;��.	��ɝ�||՗)��C�%*�"U�m��x���I��)L}�3�!�}
o]���	tI0����ϴE���ӭ�L=2j5�1:�.�Q�,���B3���ڬ���p�x�"�y��~��l�����_X�:����JG��W2#�b�JK�M�:���fE���7\�uvb-���1>� }K���K�XV�eS�j�s����5�Ӌ��C W�_є���2p�(u���؈Ş1�\����#�YJ{�G����98q���G�M�쇔��և|tZ+KL݄u����H�b�1��b�d�Ԃ���D�Π!|���ËjϏ�z�o�"�����]�"&��) V?C)׊Kѥ�R� ���(��bQc�\�hcʇ���iFk�R�'~w�Sk�����G��x8#iy<Os�7�����R�l��t�h`��W�@Ԩ >׷��
�P�,�bE@��!����߹��І�!��<l{,���Ϝ�cG�S��=�Tl/��!MD'#w;eRw�2T�!���)e�Q��T�۩�I�˝�H����X��HY�&qc;?f����;B�m��a���Y�@�?��?iͳ�ɨ���Yi��{o��ɓ��R��W���^�B��EW�y��x��q����n��m�֯�Pg���lռ��<�������B��O-/���� �fުk%���-����~�c#�W�������_�Ȗ�,��o.��/xe�����������U�pg/����H�Xɓ�"�r��@y�"gQk�}�$VW�3�FؕBcc��qP�0��H�ا(\ ��ȴ������� ��^���1�OԻ��@�'uWAH��\�QT�c�1�e�'j�M
<�o?r��(e�u���ڛ�fp��F���c�I���w���@�ԍu�,���E�	�C!�w���gFh��Q������<��V����OW�9G����o0I��N���lla]��Q��@R���`&x^�u3͜P�we�K xyg��&�]vfc^a�V��I����3�=;SnX�?|\��9��ƌT�Py	�ގo�Y�y4i�p 8V_������$H�]�n�Bj���J�Ƿ�`c�ӥS�epw+�^:�n�P�E��-�S����~��_r̴�Z�=K����>�P�T��h�!Я�q-yaа�G�&,3���.!�mƸ����V��C@`N����u����<s�;]8۔��m?|��x"0���-
���5��0���ϷfF�K{$EJ���y��nE���7�������r��7�"���.$[ز��>ǹQO��/��)G�͚>D�1Ӎ�_�G7�i�yQ���G��o,!�����r�q�_,��(�OS�9�c����@qi G��T\��ci'/���Q{�j��R�B�ٺ)?�I�����!fm�0�].�cq����cTP>�~����(�\�BX�t�P�&�f-L�Lx����@��cf�E�*�{XG� l��]i��{�_�I��o&|�׌��x!�,|mf�k*fT���=�P��8�@��1KU�����-���� .<��hL�:��-'�QA������|�W�������,R.嚳)�c���iR���L�9��\�,��u�[O/���e�Lء�ɏ����;�^�s����j�*�e̛�=~�;�X�6?����Yd�lН7)�2q*K,���3oΉ�X���2�q����e�M��8vd�9�p٦�lz��`L��j<`�#xi�`n`"�h��eL�����Sb?��'��
F������q�"�4�;]>OVV2{�,��;2��ip�������ـ0��,)��0���V���x�`���i���|+6P[W3��A�z�+`7ג3 ��a�F�5�a��Lq.�B���z�b��Ҹ��
����+��X��oH��G��f `Iw�Xo�p�$���Tz��a0U8[�ҿ>�uӮ!z���p("*z.�ݛ��x'U'��Ną$3��qrG�r�5N�v�[�͕hϑ���~�}x+�z����i������TFo�3������x`����"S �W�=-,d���d!U.���b#7AG$��A�qu�S)�������;^X3ƔH���`y�U���L�(a�&����#[XK�_����#�mdN���6�����\=�bJ��X�M��]/L��c�{������d<,6ФCv��&���I�<n��S���N����ѯ"����R����@�J�	|	��^���.|D��{B��hq�_��f{@&ǥ	���C^u�+0����<��M]��!M�0�S|�l���_hicb���S&/|	z�t�ͭ�q����=h��6��99��Pa����A��K��ܦ��O��MZ�!e?�F�:rȯ�6��mz��z-U`�	U����#ᶬ���'{�ijɊ������0��<D٨S��(��6<����1
�I�X(��(h��ğT�q�LF��ԍ�1��7���l�B��ث��,(��-yO�w��m,�/�gt*g�$]������z�4�ȂJp_��vlG�����E��&�B�(ε�Vq��zI&�_�q�.)^���U���(r~Qy�X�5���%#[\� ��G��1�5�4��A^��h��lD�uh<K;C֐�%���N�6{�E �B,2K��:pܖ�z��;��� �T�]���C�̨�#K9��(jWX�QP;!^V����{
٧Y!��G�e&�a��M���&i�8W4nѯ}w{VlŃ��Z)���A�H��A�������3H��a�� #�+�S4#V���KB����"Vj� KDz�l��#�}�+���=�<͝�_�S���B8�h-�XJ�
��[�<�����4��Қ}ȩݵ�B�Fjm��9�h� ��9Y���7���v-�:���by��l�X�lÍہ�$ �HAN�a�$�d�W ��[6���9)TR�2$��	�x��O�8��F���/�Uc����q��Pox0o��J�u��쪉��FlZ�L��f�8!���|5�P�֌ņ���9B*�>%D�9O`�s�!g�8t6�x�n���n�J�X��A,7���k,'��%�|04�ח ?�kp�/+�� �� AvU�=<�7Ŋ�6�:���o�9
�h��NdD�d���A�wf��)�@@&|w²�)̸�d�}��$ʚ6>竑�4�
������MDG�A�8-��'�H�E���v&E�q��H�_���.Dv!��xq0&d��'��b�I]��o2v
--Ų��\���S]^ٿe�n��&��1���QL���a�X�����Y���Q��U$� 5���	�\w���㐺@�^'�+� H��iq�R-���S��|2�:��7L+D(g1<(P���x�{B`7Eo�'b~�(p�q��)����K�-$O�-čQ��#���/��y��]�>%hi�(��'�M��e��K��������k��q_s@h4I@s%�OX��pv�p���C�v_͡wK�w�H�f�hcX,'͵+n8�
�IRټ�6&�ku3��]�
!b�%n�}�bV�R<���o�=�2� ��V�R	4��U_<ga
Ë$���:�0�����Z��l�����:�7���S���u����^�C ��{b:E���7����M��'�ӣ�w�l_�y�1��1��Uv5�O�,�2 ��+��/�\����&�J�%_�5`c�K�̝���Ͽ����:"��'\��,��$�<�!d:ȅ'j�� �(�D��Ad`�c�ۘ���I��Vi���7	^
��C|���;���R u�.����Ê�TwBڠ������ϒg�K�����τwAP�8v��<]�|��P�6���ڑG�3�{�����&�J�ǎagGKY��D���_��v�^t	��9�~A� z��D��3�#��q��)Ŀ�גţ��lC1���H^��2G�-�L���(Q���+[W�db�@�t+��.��
�Z��K�V0��\��^�Hxv��n5��dRE?��-I�8Eh���w��ct?R���m Gy�>TB�h�����"1֏ʁ� ۄ{�����1�i��|d����Ԉ)��l@
>)Rq*s��0�$�Z�&��*k����>�ɑ�C)��(g�=�7l"U+L��C�B�Ш�Y���@�݈��k]���&}-��>-u�9�N��$Y.���I
y�R�s�-��?Gs �ֶw���N%��H�]S�P�ے�䚢��k?r]Reo�Htzo]K(IS��w�&}�
v���Ϡ�Gz%���
��aj툣=�	ʙ틑XN�� ����֛Ⱦ�|97%Z����v��8��
�Q7"��`��~Po���!��s�s*�*l`
�~��sI��K�W�r⁾�QИE�dû�C�{б(�P-�kL�{Oq�W�iӱf 겕�[��cT8�m�;x�78Θ�,��e)cXU����/��u�m�6�Pn���wL�ߎWʲ0Jf�����Ĕ6��N|KI_�r���[��S-��<�.�c�ᨛ����3[�i���)���0��L7ˑW�#}�����Q�)J���\&QED�ɷ<�7��'̉���K������a�9��T���A!���+g�T���ab�<�J2�0I�E�>+���BX�O��ݸI�D+��l4����ߟ�����yb�V�<d��I������@������фJ�ZhS��_g�ZG���fD�������J��\l��1>�Ї+X�Ro�;�Z(²]-�( ��XМX0��] ���F^V�[�D']�A��q�]QH�0t��_�gh1K���P�}���V ���{�ó�*���>�����'��^^k��W�P�@��B�fH�ډ��b��ʫȻCW�_��Kð����_|Jq+ٌ�O1"0]\���m�cq��>3�A����0~�4�XH���?�#�QY�����4vB�����~�"׬�ޤ��^��%pܡ��B��1�Y|���.��G:�c���8 �RG!D�m����|�.ط�-�E�c�uT�cݻg���	<�E^���(����O���O]O��,��k���	|��2�;Ӈ��&y)��Ŕ^�쟹@fȹ��-���`��?�S3Jy�p2�+A�W�o���Y����ȋ�X4[�43�"F���d"�r�Mv�
v�R�fUU㳨X��z�T���� �= +tܡ�M`��UZ���ڀ��0v��lwE��Fw�(B�J_��\ʐ�)���Hc.�/�f�,�n:� ��;��a�Z���]��_I��%��͋���i �e�����-=�=�X'8��I5� J�/�y����#UE�/�բ����8txRE��E�ڢ�<����x�P�؜��@��,�B�`��!g�����d��BLq��Z�W\�Z�IϪ�_\܏-1K��C��k2�R��X�*�,�p����51��kiŢ?Y�zqA*;_�I[,6�?�V8��0�y��NT�52�=u�q������,jv��D1��@�[����;|8OD�`��jc�_�'Eh�f������\^h�LfP�J S-��	���F��W�yX������ ������%���>���H6�-A�	F�,�W�^
� ��u޾@�.�+J�*�G�,P[���	*¯��ѧp�m��'�Z6�vhФ���a�ffOtJ4�(7;;"��.�;"��S�gw�{�`�K�Q��g[ �1�MO'��}����l�@�����-/q=�(P��1�RA+s>��uRR%����`�a=t��8 i��	6o���}7%�����y�C祭�����p8��%K�}�[����Fe��~��9f��>.��6]>�U>�f���D�Z����I����`��DTN ���:��>UZ�|Q�|Atˏ� t��hh�>-�PK	1��g�ŧB��d�)ʸ�����7]W[F�͗*���Y>�����0"�!UQ��*�'�I��O��M�b�\�8ڥ,\���7�����8����<H�@��:[Z�+v:;�$.�� ���9B҉y��ƥ��L%��ڟDoV��H�Hgr��V���J�gt���8E�m�v}��!���N1M�#hڻ�N&�޹�.i����`�뚆b��Sm&`���)f�o���أ�mi���h|���c9]5������<7��[�Pc�QCg`1�%����h��-��'�5��y�3~4k��o�~�$�\B��%���u����M��X�t�y���@c�y�!���u�����b6��ެgy�,�C�H�xy�{8K�uPxd �pSI�.Ë~,�g�\��&;�)S��L%d�4�
ibE/)ĭ1K^-uR���߾�6]��u�v���3��,qƢ��[Y(J�F�.�ض�VV�\��n�i��L��2�a�HE��앀ˮ9�#�� E�M���	�qF�=9����L\�L�.��<`�iʊg��7Ug��QG@�� ��D�/ʹ�l&�Ο�onQ��i+�'�p9��Gʙ����,�z�c��8%"ͅ�/wD  _�$�A:(i���l�\��&�8/V(�녬6e��G�Ԩ_���0�����Ǌ�?} vy+`�H������7Э:�� �W�[zЦ�.mZ����~�e<��6k�wuj\_�l/Ѹ��fJ�Z����1�R�������tbu@
k�������'|c*�y�����"�p>qu}g�[���HzL!$RL ߣ��r��O��� z�Ȓ:z���r(U�j������p��gאg�s��R���:{��e!ܹ1��GY�`\W�(�S�I�/ߩ6EP� ^�KB-@]ܴcOQ��n�%Ί	�w���tIh�}��e���Ok:X.T|BVv9u�Ý3������ĵ��7{>�;sTg��p���#9;��\q:�0r*D�T�*|3�ᾒ���|I
���<g��.5�y��N<��MUAØ�w��	�ѲթK.� �q
�/5��2b�')\YcT�Yf�ux�v�\B����}��wu����(]�Mخ�����;��RU��;I��x��N�jh�9�I���\ ���������n��6�<2EW,��t�ۤ}%%��S��4�ɀ�%�n�8�w8!&8ٱ�)n(�Ԇϳ~>�tcڥ��������	?�Q���p�-?���{�?�U4�S����f����b yY�ix:C�%JL(a���B!uqmbF\8q�޶��8��*�89E4�Y1����{��O����[d,�0Ȃؘ��à\������rU�(t�x<"a��6��l���7���r�O2C�l�����X��*���&������v!�`	��_fC�5���TН��,�G�������ߑ��	h$3�����+�M?^��sj��y�.cDf5��{}���ϯ��6x�痩4	7�j.����곹��?��d��~�*R���SUc��Ȁʉ�۷�f��wvB��~�7�9��OZ��[R |��:#H�n���%ќ��W�^�Ÿ�X�Sw'C0�]�7Y�ˑ�Z�E��d�C�rs�~�L�F����7�KRָ�Z^�:f�bveOJ�冑�<+�P�Z>d>"�I��?�pH�ua�/W-�����O��Ra�RE���􂎛L���׏8�*m!� ��\�H�������H��,���NZ]�`٬�8�� C,d�^�`tBf�~��ceQ��)��Pp�Y�y�� ��Ԓb�B[
Üؾ� ")i��rNrw�n��j������^�zy`�P#D�q�=�1��>̿�1c��b�������@�������Z��R���s�A$�cZe�s���<B��7�@CjtA����ԳRp�)�qİL��4Cx��p�Q	��ޅ�*`�}����A�yN1gSx�H�D:��?m:t�R)��D$�yZ��VknMᬗ��b��)<v��WU�^��Ci%I��[�o~go=�*ݠ����A(�}���!����t�-�l/�Q��E��7]��U���Y�E�UR��s)_�c�ٸ��L�v�xt4�Әk�<>��3DB�7�)h�!y�����-�$�L�EBb�a�^���[���C^t �Uc��5wL�jWeE��6�5FV�τ>�"���Dܳ߰�X�~�������Â4�4��Cu�줤���"���(R��܌��dƦ���Xc
� ]h�|�T.`me��������V�\���i��z%�uԢ8��۫;6��	��������-�F@�"�yXV�P�m�:Ayxn�F46���(�\���z������:ڿ��N�7�5S����ס�,|�WN�*3��_�+`�>�����t~x����x޸�E_�InO�E!�ֹS}lfB�)]k_0�f���ڤƒ���
,3��]TU��^b�vS�����3y�Bd���H�����P#�X�I~N������L�F��ٽl�"ӨM���j�#�m��[ge19͚B{i"'�K/^�+� 3MV����S�I���7�L��U��H��!m�j���Z�5kV&����fw�x|1h����{��cȋ�����:4��[=������>O��i��*��a�����b7��[P�(ɼ�h�Ą������aieX&�]�Є��#Zu���O_�`
��M�IC�=��D;�8 <����u��
�����L@L,�����(-�{�����j4���A�ʄ���-9�HP�� ��Y�H�4�=},������ 9o�j8'��ƿ>�7��C�:���L�'7U`ղ����ݑ�r�$m�7�Fl�Nq��������Q�W�g,JB�o��ua���VA�X8�5a�J�'�� k����?K"�5�mG�ogIJ������	�CI5��~S'�3�@��ф��|��Q����'�~�݂�n�C�8�N��>H��׉ �ǞR�/�7��t��UBK��!h�12����k#;�]4���/l�����r���
��O��y]�eU%�`�|z�i������@d�M�u�L2�%pnJ�����mE̽�Z)�e���	Z�b����|nŊ�n$�Rh`k��;?��\Ɔ���L?x�3;��'�Y��.v�EUA�:"�m�1�������m,�2 7w�GFg�0��|]�U�G˂5�ř밍���u�74���يh����"MC"���t�,+���3|��Y��T5���Δ�e"w�y�X�g�p6���m���n͹��|T>���6�G0:��d4G�% �S��?�����ƒ�+�"!J`��)MK��� �!ͬ��zˌm��bx\y!�t{sh4m�6,w�������e[c*���̥qK�mr�M ��m����XU=PQ1�[��*}QD�����w�Q��c��}lVS��T��Mr���f\w$*p0/���v���?���;�t� �����k"���nwm�F4Mjr����ǆ��x
��fI�&_|���v�<�Z~u�ܫ�����;�����L��o�	N�y��k��F�Y�F�^��hnv�G������0��
�/VsYܤ=���m1����t,"�.^��;W]�����"�U�q��o�4��7VރV͎�h�!�t��"8×�Cp��V 6:g�hyE|�Pn/�,zs���u�a��?B�^���(�@�Az,v����>�ҿ�W��0n�o�\H�p^E'����m_��=z�v9ة-��q@��Q$�E�k�jk߸�S�I-d?	qY������w�֗�Q�9���� D�Hi�+��wH�|�L;�L����&���B]y}*�w�뛍$���@ 8��š?|W�ڂ5@�Y���ꀥJ�P���Y�L��*k����W�C���Ŝ���@��@qC�;s�m&6z�0��d���r{�ڗ������ܺX���?�l��1�QnY̧xK/�A��c��a0��6;�$��b�b��-�:g�2IQ�N~�lNxA��	cк�$�۸�.�Wƴ�L�\�/�Z��k�ո��<=#����_q"��Ȳ�d�AI�z��BY�<���_�0�
A�b+���L�E��Y���n�<��/D��2`�֯6��K�,�<������2.�9�ʖN�t
!��P+���*hcL��l�w�!�G�C�c%]k �6#��0o��<�?2���S���]�5�n���Fz������S���bXj1�����?t����m��j������'���U9�=�%��%����|���� v��R�T��߻�ί)���-`D�6}lg��b�[L�7�ps���K��,�C�͞���O$����ll��=�t<�U��X��x�Ώ|�N4@�^�2��9�J��3�I�6��ZvO5�L��
W[�����c��-zZ�tS<s�k6����Ar�dڛ>A�����)��))7A�0hL���ܷ�;mm�Ǟ��]V�b�;DÙ!��?�rx]|�Lm_Bda| ����]��u8-�O�}/FK̝j�p��=����-:!�%�X�~�oȳ\J�+��+�㦄�^��p�?�kFzQ�'=2���8��*f�VF��8(��@�	�:k6:YL�g��@�._�8$_�8�H�{9p��K�:�k���͹^j;EN6�U�ڿ0mW��BSq��Je�x�Cs\$�������&��0����v�J�q����`B�C���1�tM����T��>�\�9��؏X�~+�\���߬��6�� �ÔQX��t\��j�I��e4�"���O��[�b�C��r�­b�-�
�0��1�����Q���T uwʻ*�".���C	ɪ��� ��խ���K�b���db��(Dk[]9�J���
��<���{����t��W�?�&a���uw���P:�j��G>�K�6b@��A�
�G�ވ�]��)v��Ǥm%t��tH��h��ǌ��sv���|�jm��#j��(�>�ym��.����W��x!�k�QO>��-����y,r��E�*K���>=�-����:���m�&��4���tǑ�`/��V�خ��S��Q�#��6���QO��mYO-�oL��?f�н=��m�����E����k����3�^�tOSB�~Y�xv��l�y��u�aL���Uz�3M��:����;�Ci!���O���{�ą�:j�Pύ�a(1�]�z_	�3��;�v 6�!�M�m�����Bajo�x�X&o~��P{/#��Jm���8n����K#R"�d���1�cw��RO���t� k���M�s݌�����\;7�� �0�cq5/�H�k�D!�6�"�a��v���Ls�S��[������4�iD
З&�ߕ0�czr��=3��ᬘjfR��)u&S2�|nՎR<�I@�&S�T��	_��6�:�����q9r����*Ny��e{�� m�o���~Y�H�=��	Pn���f�o	�,nm�W����6�T�11�#,u2��C��1ѯ�NeGhA�Ј�L0�Y,;� �[��L#���	t� �������僀Ǭn���M�P��'�<�ziZ�ikZG{`�V�q��XP�1�"��F�h�M`)�]�_�	y�ho�6f����I�+7hЃ
��Q���h��a�O�
��1 l��Tb�f{E��bԺIQU�jXԖ�&3�V헱%s��ȇWJb��7�����/��g���ZP�%�SQ�KR��R�^�.V�R{#��y-�
R�3Lν��l�-+�$�����������)&�3��G�#��	I0��f�H�^��!�v(4f@Ř��'�yf!'��S��Я����k����N�������Y�F2�,h����)P����y2�(�Q3�T���C���L�2{�(ٮK�69�/	��U�~�5wb��L�։�r����RV��/�O���9�ҩ���X1�2�m����[�
�.ͫn�th-:f����_��34�%>�ͳ+E��&k���6y��%�.��胬"��vϖ#��͈o�@7<����siMiX-������9��ҟ^��׎�_� C��Z� m�B�2��k���@
��g��c�ҡ������?�d,���Q���g�k��i�,�`rh�7^?�N�u���Z��NW$%o�OlM���_�x�E?�Z��w�z��Kq�2����@�s�pu�_ ��Fҟa=�.Ѓ�e�C�ʣg��;:�I�j�5��_���ں��)��Ȉ݉�����EW��쎙[0!�D�kり���A��o��$m�浫g�^Z�9p�~�p�X�>E١2�&����	[�'�7M+eع%�8�*��Z�8�x�2c(�p�!=<f`gHi9R-�s��ߦ8����� ���ª�89���9��([�@�/OLS�#�pQS��b��j�|��̱�,�'6t~E�)�C���J�v�z��
j��y'��'L����{��y��P[�Z�[1wC���T;�t���"�>��G��T/�(&H-��a+E���T�htVY���[��K��:��dy5S�;���d�1w��F-\zq'�.a�ס밃8 �c��9tWƗ&�oxT�[R��1�Bn[X=~�e��� ���Ԃ ^�d���r��L1��+�SښF��C��c_5����}g���ײ�>5s�g���q��Z
?��[�����^����<""��X�����0QW)oP�2����H;�J0���:�S^wS��24�:�WonDi%7	p��=�6Cv��RgKg���x���ʻ�7�`�I����F:v;6�q����9#Q�v�Fx4��n+�A����C �� %0
�������{�d�Z��#W--���T�=�k�j�{&��0;�Y�I����%�{���O���Iu�g����|���T�L���R�W�_{�+�u��#t�kc�@=O�a��}7G��S��1K`e53Z��D�&�C������z�/e�|�̥�oі}<h*�������7/RПrr\��ʑ������w�a#G�k�(�?�"QA���c������w_��)������f���E��EeZ����ﻧ5�	+K��ZN�EJ��%��UD�h���{�%[��zx2G�`_�i����!��ԫ���������|�4C�\7����8�>�i�d���%�.�փs��#�w#�+�xd�&KJ�:��̿�+��Ɛ��Dj�л0ޗ�;Ib� �kҥ4�T��	�'_:��T�<B�(GD褯r�#>*%��
����/�EEL<���@V_z�2�`�Y��x�$n͝P��ٻw�N,�cΓvՔ��Zcs�s%�(�,�\-���	�� �����_��ҍp��,ץ�36�t�����I�"�Ay��F���fG�S�T�5K�K�������A������Q�7�k���I<�_�pS��B��(?��4��%
7Z*�6��k�g���=/��#j�,}6��C�H�x��My����M���U"�Cn��zo��J3$VV�����Җ�?�*�.�+	D�R6hĄ�R�fy�U�{�ܦ���Le��x��7�"�}�~�癅Ҡ��\��8�GG��x�ʂ�#��=4-�<��]�<*��w�@���pF�c�Y���l<:~�Z�-2"�C���@3@�N���Iofy��N<A����[`�^��=�q$�&��[�.4vM����`�_��!J�A��D��(�aN[�!���+ʬ��I_Q�蛺��,�P����f�¡Ok��x��R�DԖdw\,w����I������dʐc���c�ə���z�s�����A$�9�ޞm�ī+��U��~>�2��� ����Q�]�<�(-�`]L�����a��Mx�?;nk�	�LTٗ���SVu�6@�{"E����s��P�r\��A�3�ٴ$Ѕb��y-�@��-+M���P�0}d�Ba�wP5�{D�J���緐���6C~��U-j���S{=E� H&z�%�獽=AjH��<9���'Q@�uЁVR\6!e7D������O��1)�c��S�'�P�(�����jl~�Z�y����N�©1����o2��$/���mD��G^���V��W
�"��,&)Et=���!�UV뷡�,j�#�Ő-��1��p �n��]$�To6}*��`q����~.��xV��#)]�Gv��ޱ��2*��L��p�� �,B�31�G��b-L�̳ݘp���	qqF�\ƾy�W�^A���wz���������~�)��2ܺ�!Sc�
$w�:��F��i紺��T-��$k��>��\8wAi��ST�e���w�s��R'�Q�n�;aDf��.�M��+���)�:UU���{�#���`�qd���Ba��g�J�p�~�Z9�Қn`0�"L�6�'3�C9�{:�sA�;+�_�G��K��"	�0������Q<��?S�L���g�Fy�.%�v��$���B\��K:X�~l�b�t"6��������"l�!�J��u9Ox-?���7ܠ��k#$���R����*g��w��s��R%m�O7��٢����;��o�ʸ�:�o�g��K��-3:��vf���~���~ ��_�{\�)�t��v�ib��>[��@�^ 	g>����O1h����7��k��J�C��Wॿ�y���P��_�U6����9uS�A?�7�5�R���Z����=v�4�p_G�rv�ٍ�v����%&�b��ZU�r"��3{���z�O��-B֏n�����2��']�3|n���^�(Ũ��	:7�?	�e��*�7?�W�S�u�X[�8��|���S�������Ɂ�E 
�@�\ZG���Y��
��Ҧ���II�L��	��h�c 2�Jm)�rP5ט�Ì�Y(L\���\��O���(8�r�<	Q ��:�s3�+���s��A����1x��m�Ƨ�(!M?/~
�V����%Ƃ[X�Y�U��o�x�����u��c.�ۃu�݂�`9H������Y�N�е^_إW��,��r��oLVhXR	%|0�H~Nwn/p�J"g,��e~��k*4�׎w-
�tx� @��ͅ�2et���n�x]�,��*U��	 o�b��k�=��z��q1�٘������۫a�z�x��s��pH+�����t��Vh�ɮ#�����܂Rs�NNʀ���b�Tk��h OH���/5��}6��l����oC�h�N���J+62I�k}$�~ؤ�ex�Z$��n��4b�:�5g՚f�i��I%��9��T��5�\E2��ѩ}��"�6EW^�6��E�h�{0��G�p�ShqP��5�������;�0/I��z���f/�\Q5X�\P�VV"�@	F�z!]:�b&�D����p��S���k9�<t�bzp%	W�#@��d�6�4�)��Y�\5��Z��;�9�>g@~b����Rf/~`�{�I[iv�D�~���+܆݋E����d��͛�;���ۈU�1s�3":�z2M�;�[3�g �=�=�7(sҺ�A(��`��tFF�Cx�̸�-�CW$[C�������شy�!֙��nFw����"��Wh����@��@�'-Q?ME�X'�:UB�"��6�����:危d�?��`���®<$<�P ��='s3l�>��j֓%*��r�7�.�Ra�1ė����(�v�؇��l'�l�ߧ�	S����J?/D��ȣ7VJ�\d�E�0�q��Q�-T�u!)�N*pw�P���'���rtng*�\:��]R�0����j����W[�ǘ-Di7��s��vgh��fG�7��+L�.7�S�eԹH�t~�x)-�({�e�4Yq6����Z�11K���Q���e߱���Bʺl�-4@���Xl��
{H	��:��/l��i���A��>fg�^�Tle�D��&����@��=U��� <Y��tT��Ej�%�z��/�VYNu�x��zA�����L�S<"΁���)��T�c���>�ȼ<�#���a}��R��AH���*Fc��=>���I�,<Q#��?�#+�r�4�woV4b!�腱y��խ��z$��R��A荽C��fý�r-jU'�c�d�
�)�%�Zb��*�EH��:��f�h.T����O~�����g��hD)^���%�� Kt� ϖz*l
����:�w w?*L)v*�9ȞE'=b��'���i����ޘ�T�`r�� �f�D�XW��LߐD%�h$/eK��K+������I�A� ����M1����Ct� �k6�@]�l$�[4R��}��,]�,���Y,$L���]I���<�bRz�ԁm�Uf^:����o�	�qZ�,��f�'�Uk	p�R�Y�ED*҇�+�T�:V��?�Ca͇NPɋ�X�B�*�sYiu;����Wr3��27�s��� �+T�f��v�u������U�+a����	U�-��)�;�i� <J�Rی��l3D�pP%B�?&�?Q ���~��F[=��/��!o�	�2���;c��=�T���|��0M��E[TǶ9ք��3<Ge8���*~R� �
���ǆT�:u���/�xs�J�Д��w}�@�O-����xv�?��Y����G��'�Ց.�T+�Ѓ�y,�F��#A+#Â<(k�o�U:A��|��n��=���-A�I��f��W쨺�%v�;Mr��-^�{� �x<�;)J֕����3[k���&�Ӵ�0�}���4�T�,<��W�9���[sc��LY.!�G@v��sr!�CP�6�e���Qa̪9���	��ϲ^�.U�鼲L�U�SW�!	������_G%�l�,Z���C����_aF�L*��;�o^s��)��YĹ �=)�v�;Q�5������@m��L�#ʞ���d��Tߍ^h���*��\�"�[����GT�I+�9�<r=��%����t�kv�c����J�8��b�_�8�ZjZ<��e-��:��X�L[/�'֒ReL7*�Mf����n�����(l��r�Bod{'��k�ڶ�h���i`f��F��"Q�v�SD�����z|�I%Z�wE�ح�`[��}>h�b��d�Iܶ�����0��	%�'@�Oϧ��@9�2��0���Ī��f���a#nY5�k`ˎ?v����9v%;.�t��tË����e}�l��K�>�H�8����S��ưn6�cH�`�y�xC�d{vqF����T�qao/0XZ��)'�Y{�����iI�&�m�d��oZ��E�'�p �G6�>���`b�ƯU���M6�,�8Uc17����	�1ޝ�_e-����[��5��T�_q�T�e�e�u�,$tφ�*�XY7�]�b��`��&8�T�A�+v��E§�bV�2�V�������<.��5�]|4+ ��Q��"m���YSY���_�BY�A���򆺫�upr��ٻ�Ճ^ű���1�f�r��n$֏�˟���l��A[�ά�I���ȯ,��C��0�98XQ�����jՖ
@�=MS�ƿ����*���s����F��.�W����pi�	B4�ƀJqbP}�k�2�"�OX��mO",N{2oHd��K|$|:�ƵC*%�{�J�"B!��<}�o�O5j;�e)"`�0�rs��D4}C��M7gI�㺲c;^k�ԅ-��C�Z��}�QЩ8�pL��z�Q�K&g�s+��J��"��Z�y���A�+��e���b+��$4w&<�ӏ���:f��R�2�20��]�f�@\ko�D�3s�Pp?�%��:H�"�a��F���B���^k���9l'{�<A'lt���ʶ�V�p�}3�;d<a/US���k�
��E��[~����Z����9���t,� ��4m��ǼnG��r+�fS�'t�6��99�\����߄@���i�V�2�ό�|-���@��5�`�Co$��Ͼϊ�Ĺ� *�\�*����C���,�c�):�J/���TS���`�7���A�m=�[���e&���W����屫0N[���2��]V�1o�u_���~���jP�������XD+s��t���UY4��Z�lo�����,�-�St����Oŧ+r���ۓ�Z��tȮ�;p��XnK�ij/���v�R����6��q�ES)ď�۲�ͺ���l��Hx�6��po)���$�,����^��pl@O�D'�|���؍+w�m#~�lG$9K�N��"��#ʩ���1[Ș&�Οa�s]m2ru3Fc����с�R8�W!�+(F�<��|�n�u��a6�
���O�/��'�a�����|I��?y6;�Bl.�"b�I��u��v�@+ձC=���F����Q{U}a8�}��7%fM�⤏o��a�];�b����b��6lu���W2�$�G1P'�0}���� z�'�mZzX��a�Ǩ�J��X�E�;/�2ܓg�E6C��W+��>�K�/�E�6����$ϵ���o���O:1��O�����V���0��vP(ؒ"d���*1e�(%�Ǒ�$�[�X6�j`|�V���b�ju�v�Wp�R|M3%��{��m��������R�߄aJU��r]���M\#?}��ײ��8\^��|�q9� "ޏv� WT��g�v^��Dv��D�FiL+�&wn�&!��c�6001��BR�`$Fg�oR{���33�0��Y��� �/ M����bo�̸����<l^�^Ϫ��1�x��K�c�%|�<%jL�y8��L1�q&�˵�x�.�]a�R��jUD�vte#>u�>�i*`�m{4���=��4�!��O�ac�" ��B���I��`�9M��JV�'����׹�WjxU�VL��{o�<���I�r��Ew���jx���H]�4)K�k���}�8c���ݚ�t��>�������ҷ��C�k��0��Z���L�/�[s��2�V8�5Z��w��-4��8�`/n�� �ԙtL�I�/�&Z^�čr����%:xt�VΧ�%TJ#�&���)ӆ�����bf��z.)j�=,��������%�4y����̲�"�I��[��6�����7�umB�*�p��E*���U&؈�B�R��E�{ p�r��OC��Am'�޸��σ��,y��/8��$�r;��p
�r�t�|�&���v����9�¥K/�lC�LFdOIJK��o5�S��'fS�֦���}v�/^�	+��������w�׹uUU�^d*��gy�G����yϫ�=���ᛎvl�}��h�R�{Ɵ�����p}n%��$���}��B�����u#��롳�IՂ2��0����cr�{�;^r��ݢbI���cP���v=�x���ո@�-�����)��T�RFl]���M%�������'n#K�J�:R9��t��"B" ���Z���e�dZU�dDT$p�P�@^�/9���}�8}�7l��������5r)� ,�H�b3����b�0(�e 7ߑ�6����fz|���*��f�5ee��z�����2�6�
�?xm����(��h��,��U'I������"�fN3v�G���'�?<�ɗ>M�>	�����=�� [�R5����t��}�������"�m!'1�V�d���K�O�:,�A/.=���SR��ss�����+�0���$9c�[D��h�.�6�v��Kf�!�2�i�D��7���х���� kpq��������r�c!���\'����M��kؿ��	��`:�jȫBjр{tn10���=צ��t:7���_��3��kh�<)��R5+~b%���*�*Y��`o?��}���`C�m	�^;~=@G�E��o-�[`/�97S2%G�鬖ӗ`lڏ���W|�J: ��nQ8���XO<<V=f#��ᨭ�4�I���%�<��J��Qꋀ��ZF0��2�ÃoW��g=���΂l1/c;�y��]w7}�8[:�'����v�qQ�rҒ�[:�U\R3�¸���g5�W{�Z��cj��'�M��)��J����B%@�u9��_7Ќ��5�w���g�IFPZ�՘N������2Q��ҡCX�m��e�Z�h��z�Kj'��;�ĝZ�s9("��N�?��-M@W��GVt�{B� j_�$�5D��p�j�s1+qZj	��a�y;\�4Ͷ�Bs	�K+��SKQ=ۓ�y�[�4yX��D���4^�(Y��'���/��W������gp9r�?$�#�?)�	�J,&i�Z�� ���R���3����+�OЕ�E���fq��r�n=�$�{݈bW����qt�Ͷ�ꇜ���`5Y�h���J6�z;���#������3f�N�"�"fb�*�j�b�t0£Zz���&.�	C�#'밁���y���A����0%���0iH�����a�j�1����s\���e� �ЩUN��8:h�ݯ�g��{��Ry����.�>@y]�,�L��O'=�.b�0�	�u�3
���ָ��9�9g�lΤ��%D:գ[�pei��MQ���	�/_��WO1��z�Ġ�5��7�;��ũ����m��^��p��?�C�����bn\���ǥ4D��qz:J�*�k7�(V�X���\�yxm@�4�d��y�7��URF���zjl���q��cטu��Vm:���uZ���vGӶ'��7H��S�{8�g�{[��������%�����=<�N��J��+�&���j*f���ȋ� .o�{;+��AN�+͒v�$0�Y�D*�z�;o��Y�r׉ {\�>�,&-:�ֽ'�"����<�2��*#+]$o�#����M'�^�	��i��l�O�g^w<=�f���Z,X%eٷ�y���e��ɹ�XV<�r�y�JO��2٣�����c����XZшd�����F�;�y
K��Dڪ%��tT�&��߄PQ�p�]��,#7Z>��v�D���
��.�@ƤU2�m�T
[�^-m������P���f����ݗ�󰚎�����v#�S'�n��������xS���d;���D�50G�0�"��A�c��m��*�1���:!wpH�������,?:<�}�6�����so�;h[r�5<@��� lH���h�
������j�� ?ۤ��A����]�|�c�UȚ����N������w��l���Y��`��	K�|����Sǭ#OL3I-�+5o3�3�`�>z�*̍�%�ݡ�jo��ڔ1Nn�<�{ �|�?�ki��"�{��G�G;H�tإ?q���c9�d$��z��(���#�/�Ԡ��ڰ-�}|��U�I�|��.�D��؋\t����A�j��7q��.����
N�cE�J�g]&�;�����&�u�[>b��zK}n�&�*��9G�4�ρ�����Ooʐ�a�ӇF���y�I���UwF�ܾ���h�o-z�B3N��ǝי*ٞF�5w��*
?��]��t+��U@9���D�07�:�\\}
�1}B)o�����Yiu�ϷM0T60�t �{ls���x;�W�`/ߧ����X�D�!a�˷��6?L�+Aľ#��.ʮ�=dg�W�9��]D�O"cs5hf@�/�`;y�a����pG�w*��lyJg�%�l�� 8BJ\�#8��8,�S��B�nG�O�jL�\�\Z����WXh���5'I����5�a�������/�Z8��6KhEci}��o٥+�E_E>��j���R�����t���o��Lh�Q*ꬓv5r�ET}'��u#z_k��T������:<�J�L#��}��
'�c��P�q���Vs����R��L�p�hi`U��3e{ �߭�>��o����-�\��8��ℸl��B.�}�̹M�Y�k�l�����*�"��KKr2�Ay�y�5��N�#�o��k[�j2	W��%�8����P�G������a��6�F��V�:q0��<����D�G�O��#bf}S�ّ!�pDI�BE�vJ�V����w�w�1T��%��n# J�Q��&�"�o�"�K�Ԛ���6"4N:S��\M��Un���UiF�������3���_�Ǡ�Z����h+��S�L�FG���A���&�J�8��Is�-�~WB��)��1Xq�V�zw1N�@�)��>�#�ׂʨF�/PG�ޘ�z�j�N~w�Pmǻ�j�P��O$6Va�����Z`D��Q�����BI	�Ġ�������7긑KA\Z�`i8J]P��hB�"�q҄V��>��P(��lF@��i��n�\�=�+�C�?�:��;�3��N��^G#�:��V��,+��;%٫"�i����iϪ�*�
:+_\�y�zl
,���' �c��t�Ffė���3�8�t�H1�@8�_��t��	)[��%����]7:4Q����. ��K�O���#�<���qf�Gw��#�PAR_:6"��r��z���i\��`b��&�0�9�w��bj�:�\u �X�\���p��8r`	��(<�ؓ#�E��������N�b`
�C�o�0|cϮ<bǾßʀy�︁v=�7��|�5	��e�Q�Ӎ3�dq�а��l�'R�p2w�h~��6h���U�]*����Jg1�̑+k�C���y�O�Z%�t>Q�?��
�2x?���Ȇ��!�ê�p
)"��+��.��I����1}&��)��""�(���;�� ���+ڵ�	���۵JN���\�TI�)�l�9;�H�I���!욵~�c���c�~��`�%��^cy�il[��
�����'�o&�*6�dlGl��.#݋�}�} ����`�CX�3�6����1AKz���{�ά"]L�&v ��I��'��_��� D�}�6�����1gd@C]���##�gY��@������q?�Q��[�bU̘h�V��~���٢$L.BgѾ2}av�ޘ�AOL	3� q+���.)��ɔ�?h9�P��,��l��F�,g����%u�V�F#���R��$����덌)#�C��_!tO�2�sLrErDQ�d-f$�%5�s�v�܇�`W.�=b'|ʋ�H�e_xV��H��.{��c/����@����)����D9Ka`���T~%�ٸ JV1?��� ��S��YGGrEf� Vp�wJ���0��j����*U4��^Fg���M�;���1�~���o�� ���N�X��>�g.kS���[Q B.�VDU���ڍy7�H��6����Y_�ouֳ4)�6W�d+�a;�H&�;�i�s��&��2W��CYC*]U��$lN`WVQ��� y�7yR�2ҁ4��I�Xz]�� o����(�4s�&��;�VW+J� �Lҷz�^![��(ςr��Tk�����tI�_���P��z��mI��hN��܆��6sPsl�H'?S�f�!�A�@HP��C��q���������X��_s���ΔN�e�
*�P�����mܤý.8~"�bj/��D$W*�SaZ2-���wQs�{7����+J��-f�+[-���\���(�g��.��qKL_u��s3����!>��d���<93"?���ڢ8�DѾn�p 
���ֆ4�&ǈ��1]X�\�?�~�;V�q]
��B���3~@QV��L��uf��TB_я���"�rx,�9K]bҷA�H�P��|�3ݟ=��(,�̲�"���%�ĕo<�v6P�=�~�ѷ>'����Hf��D�0Y�#ua!}��e�q����r�`���M�
t��9��d�'���R`��v1�/O�=kO6#���Џ�W���P����R����~�d�#��2���5깝�ͫĜrPZzfs���P�zH7޻U����!_���g��n�.�ݿ���}�%�l1�,�=�5��>����i���jÿ��/8 U�C������Kų7�l�D��̝��p4S�^�ٗ��!��wm	c -�%k��'��&p�4Fۏ,2k���s���X����'��4�����7v_�e$��
r|�KO�� ����Ee��ܰK�ȫ}�jzn�O���1��3n�V���+��d;�>� ��YN�v����Կ�j�2�h���:KX_���*%�R�s�?Aϟ�M�cBKB�'�d�[S`I&���\�!$��F�1��y�B?�������^�v ���~�y�gm�� W�3�a��4��]d�=7�>co�W�	w�?�� �vk࿘Iп ��Q�;�b�g�.DOtC�m���-�?}��V��;e�"� ���L�>/��Y�B�_h�v�sE�^�j+溏�<[�c�8ୢ����L[��&�Vy�rKP^�2r]AI��`�o���⾺d|����WC���Y�
W��.�G�R.`ız��|�_Z�}8Ϳ�'X%�(Z�%���.�W��U_�M/H;�;eM���d�O�X��nt)V����á8iG�����m�#.ӝ�k����ϧ��䀤���)a���T߲	�������qQ���)Y���E_��j���cP�a��A�[Y��g������-����Z�b ���h�MW���=ݼ�����x��;e/f��{�b�H����ꢨ7�,�b`�`X ���LV`�)�l�t���7Kl�}�Ҫ�	WW�(�k:� J\�ƚ���s׃Sai��>�L�����\9^��FS��Oa���-QpN�.�s���oĊ?��h��yP,�G�*D��� 5�zY��K�>�;☳*嬭׿N��V�R�LΟ�^�]��B��5�B�n#�a1�z�*�T7�(�OR*zu&���]�Ly<5�
V��/��
S�>T���u��Q'*��]�l�*K��t�L�Kl(�-�x�S��t�v�r��tz��H=�w#�ۣ�ѤF�/�mQa��?*S@��U]�l@.>p��C�"A0�+;>�8`�d?A�����W�b���A���V�L�r�Z���=�d��jK�U �Y�w��r�qt76;���G|���ڵ1R� �0�X���&RO����95G��0�bޣ�?��?����~}V�N��S��i�r_扑a FӚH�i��m8+{ԉ{��s��8VA,]H��@h���`}_)���5��k�"�-�NSE`&��
��n������աF��(����D�][��E�]~����[�Z�nPe���JgOsJ�&�>ɝ9ɱ�ls�I�WT��e�	�ے�y�(�Ŭ��\j��1S�łl 3*ɨc
7�z�(뮣�C�l�[݈�D4Z_��v�sX[�@r��(+�u�o�����9���|/k�o�6(���u�
V���9|YH�!@�֤җ���"�Y9F%��i�x|�@��7[���f+T�,QU��i�hk���(}n���J�a16Z\�k��k��w$���@�$��r�)���ںVz|�2�s� �ї1S�E���-]#;;w2�l��mH�{5f^��IY�_�}+��찘	T��������K��q��MS�"��o�5���y.�\,���w[!���8��2��wm��=:f/镼=�o�����)��(�u6�&�~"'ɿ����?5�Z���v�o��LOK)V���b�$�a*�-+F�����{���17M�=�`J�����|�~�`�0(��Q��UC0_��C�$`����K3?�m��(PɌ#/JW~�7�f�%1��J^��^ޙ�z� a��wvs���>�<it	�۹l��G�D�!�rޓ�YKqFTĖ�_��%(�;1�u,{;`:{4ct������o*��+>F���e͔Jz�?���4qG���.�{�5������jl�(�ď���<��_�(!�����U	�0���<��Z�韂�"�l����|],24;GNNQ��b��m��������ߢ(���I9��$�����޸�p��N�H�Go�@D��@ j?/.��j|�j�4���F��3�c�E������R��S��Y:����*A;��a?*o�
(���mk:V�@�=�ҍJ$��9���{^��*�R�G�
�3�Hy��Z�����I�t�Y�y��ҋz�^����_;ЩVM�V�M4�և��H��������,�~����9`�t+��E{"����M|4��E����Y=��6�Ɯ��-���E��|�{�Miђ�hgL���o��5qv0qi��{4x�����+����W��k
A �_���spQ2Bm޶����5�i2�t	�;�L��&'��\P�`�ݰ�a�b��N����&ЩV���v�{��<֣�.u-5��`NY�gm�U�k�|��v)�Mu4$[刃,����V��+�������=��6�*u\['�����!����H�U�]�[d\�L2Ԡ����>4���
W��ƎsZ�x78H�~/gGor�HT-����8�tr	��ͣ�KD&�Qܪ�؇� WX���c̹H���=A��@&o���+��t(ώ0Z�+p���u�[e	M���;A�/e��h�XrK�|�*)_� 2Ԗ��M��3�'��7`��DV�@��k���vM�hu��U�FwI�$#�s����'���ao����P��"tbR�;Q��rK>?������W�����	ʬ5��k���3�7��"\����/�DS�M%eZMmٌ�'��bzQ;q��I��=x>���x���͌/h�F{���-Q���@�RT.J��6�I)ڗ`u%��h'U�k��$�	"x#���jq�~�����ը��t1�L��=����/���xH�'.i��Q���@68�t�R�-�BQ�3J �y#�.�C���� L)JK��hj�i���K�RC��Xef�����Q}|%���E�}���S
k�Ɨ��]_fl�sd@�w{�v*"f`yp�H��ĂO`l3�Úeǃ�ɻ�>A���{�ML;�R��(X���Ƭgf�;f21�kH�6�_�~0%�Ӽ=�	ڇ3�۷\������6]-�g,��d�#�w�����.y�XR����V	7'�A42\v���rW9�gK=�@_�U*׎|-���?��4��/�Q�]z��B2�N�U�ۂp�M�,t�O�����Zn��w��Q���p�R��t���G���R�@'���b1ܮ	 j8=�y!����������71�Xѧj��ȻІUp➊I�Ǔ:->�y֢eU|��MfEAE�R����qŒZ��u�6Di�v�
x��i^O[Lyt����^�Q��i��lLt��Bi��W �~��iε�WM��.{����_����!3S����Exսn�O���~����>����RM��x��,ff�'�G��ց�~m-(n߫}Ok�Ο� �!�X�R[K�Py�oLR�5���/<��`�ɠż�E�!��G̯�p�ݔ_{�X�Y���0?�f �{�^�.3I�E�/^6�[Ʋ�#�FPG:�5�#��Q{�����&4]4(Χі�T�<$��k�}��NB,�
٢�;���c,mx�G�)L늿|_�Q�Q��)�T�XH�n�7rZA��>	��>�xi�� ���%���4�תك�?.�O~N׾���3ǖ��7���ջ\bm_t�����b��1U"��r~>�F(�_ ��|�Z�Op�7�U2dG_�j�o��@M�>K7����Yd0����NZ�_(K�3}��n�6gb#�vm�P�t�=���qUP��*F*Y��iщ⋓�����ދ������ᕟ����Iʅ�S�����f_�E����R��W*U�eȖVI�?��,o<�K���a�ʭgS�{bmป^a�c��O4к�v��2@28v�e�;N�G�����A*�фt��[1te;�`O�u��>��c�i������L�N��(�)�a��7����jLIO��]�S���0Qϓ�c�����3�.��Sh�4lN�o w���r\=Q���٣�k؁��s 6^"
l�W�M;��%��6�)��;��C^'d�V�["�hpY�ڂ֒�240W��R�Ԓ��/��E��ιmH0�$'�h��\�
�+R����D;�/���Y��Y[����?LVZ��*&��a�-�fS��_a�~��>z�D�Xiw���x����fĽ�P)5��i���}�Z��ĻI��f����0�Y�R�K�B{��Ht$������|�P��~��"~q�s�K���gl�8և=(ϣ�Վ�>�J[do��OY�Υvp�ey"��lf!��j��Yޙ���D�c��,uvtg"ap��Q�ry)T��ۙFɔ~�"�[l�� l�dO���'��8aS�\�Hƴ�D:�q�����h�IeL����Q��-�+�H�+:#}�nM��_�m.�~�4{�U *�u�Њ���NῆT�d���=W6|�-җ1��;�����p9K��{W�p�Zxm�~/&\xn���4g�2���E y읬����M�4*~�C�J$"a�&3	�����5@��-�����F	�}���m(=�mlB��!v����C6�B'�1��>�;��?k����^�Ds��e�25�Yn�ݗ6��]-�`��l�&.�<A�-̊�����l�U�z�C�5��^Ԙ���c����$��'�?}%cp&!�\�2�(r� ���HL^��4�˻*��e���Y��H)�?��<�ͨ���.a�lP�4CپN�`X��7X|M��8`A�k"\��o2D�����Gxy�Omiep�,�r��N��p�q��kC���h%-��f�9%����n�� p�z���\�a�9eՁ	o,���ә�Ij7�������x�vD�(~û�k���i��v��@_,��/T�����+/��n!�$��lf	�%��;BHɗ�^Z|��K�Y>r\��Mr�0ŢkZ�Ч	b%��fS8���FC��^O}�K��0Z�"��]#n�/�B,�����⺆���,>���wPN{Jk�7�M$ꭅN�q_����˴x6�6�̾��S��1��$�b�]�q��$����Q�}�kS�����[%��e��@%f�>����
�(c������p(C�v,�/�A��1�\��/R#8��ڻ�^�f,T�d�K%�ɻ����QI|c�2�l�9�����\�jA;E5CyU�j]�|:h8CTm�u�= �i44�:a�9�m,Ȍ�U-l�5;k׵�s�կeL�&��h�E)��C��:<3�^�ܱ�4��O2v�J`C��
W��Ei�9�<��h.soP�m2���^G.�RN�ʷ`d4��S�z��[y�B�nڃ�sms���q��yu�p����I�������pP3�g��:7#�]ȉ�o�|����@�װ�ݑ۶@M#��!\�g@���W�QK=R�^
^Gۋ�P�U��~��	�x��w�ڣ���|y-E�eq�����#��=����L"�D�d߫��9���J�eO۟ٯ~���û>���4Z��~��&}ۢ�AH⪱��_���:H��`1|(h��4fZ�zM�َ�	���f��}1���?q*�� P7���%Nј��nd�46|��}d��P{�����(_+QQX�h|7��UQ�I�{l)/k�����/BϏ����d��������g��'�$q%SCPZ��Fg�\>��L���V�.����C#�@�<�)*�+�p!���z�Bv�4�V�IWW��GE�nk�"�\C�!|87�<�W4� B �Dݲ82�#_���]�c�5t�o������;��#Y�m�#y
�}�x0k�4bd���&&�v� _���ȁ�XıV�?��`c �(��-���K�7��V���˟��a�B47�7Ĝ��b18��U/WiO���c^G�\f��+>Q(3aK���9�����(�".�/����-#��`����������*Pc�R���754/rY�ƭ�_���)D.���"���(-@��f�|fa]��J�fq �W�J�R�
�a=arlh�Bn��s���.Yp��Q��g���#�օ�5k�9�-#�����@���.L�
-}A���	�r�at"����~���p#�P�܄
�`x^U��Lč1��:)b�P�:V��������$���΢�w�)��Dd^�q����L+�̘s!�-x��DA63��b�;���g.�'�=�_�A�ODa	:���쑘!����84t:�P�y4�9��n5$��.y!fV����������Gͷ�8�/�j=t_�v 3Zǈ|m��Lo*nF"�*�1S��E��D�{Yu�4�Y��w�$� Ċ��³�E3m�(����~�e�bcW
J�~�֏���d	g��^�9Z1�bD�g"��G,�a��O�{�\��x�� ��'^�*v�yV1|�o�� �5s2�j6x[�Gb!��`%W�4�?��:��J�b_1�4�9��2����Oog�d�ի�¹�>�����s<������`�X��*�����J���F���wT-Y�s����3Eڕ([�|��.9�O����}����^?|��W�ΰ��!��3�X���,݇��,�q��ou���r��t��%>d=�~ue����.��E��얱��4E�3"���~�Cʲ�෤R�t��+�;a&��n��%�n����g�Y|�Y𽚨�����'3�eJ�����S�WӾg/��3z�v�8G���w)\M_�ذ�ݜ\>��w����&�H-
�G5	*�[Vw��T�w��Ah���Վ\���q�dŎ(F�LV̧�JN&$eN�t�,��퓸��!�22?���Q�٘�0;�y2��0�%�z��U:7����eh'e��[�B+�w��>F�	�[�$�0qQ��<E�l�VB��rApL�v���(H,�{Z��q��w�f-��w�K{١�lG�k�#�~/!bu���R#߃�Y����!_�s�[W);P��ۖ��q�\�ϙ��T�4/��k����738q韽Pc���꯹sZ���bG�o��03W2(�����?F��n"�M�AC'��R}�9��fٝ��P�]����9��~n��ä���m9�eAm� ��rT`Oٽ��e8w�'ӫ!��t��bX8=�	�if0������`�o�@��2�g���p�R�L��}j;�<�%�̷��Յ�����g���a�q�}���.�1�n������Z=��չ�^��!,)�-z�F�4~���������~�)<�Ukj�Q�ͅ��[>���wmJ��q��)���͸�,LY�	�$�g�S�|�P��ǈ:/j�:��"�_H��$���Ɵx�*Pj� �xa�j���h��-�>�'��0 3���@��c/����s�v'����E�%A6������Jɵ!�c�`�(3�V\Si�y�1�/�!��, ��Fҋ���n$�żH7��u	I7 �DN�ϔ{UT*A�̎�����>/)�鏰���D���{x�QC��#ծ�P��Ŝ>T����U�kږl�����a����;_:bo��%spR@��ĭ���I�����9����W�7�˹�V�j�����ztHҾi�K�,���d�tRY��>��(�5�KǟtQr���3jI����r�5Z�q q߰���ӂ�1~�Ђ( _�S�v�کؖ�u�zhx(�w�@��0��4lT���
�ʊT������^k�]K�^��M���ٚ� �P�V������*<�G��_\�|�ք�ƁP�NHL=�(�z�&���|�P�<j��	{f_�.$�q���c�S�㇥W��C��a�p:��L@�u��vn�Pgߡ���r�H��OW��8��5�Ů�� &}�1KV��%6����8�s����EZp����s<��|<�AU|��ۍH��x_��j��
q%��Њ�t��59���'�GEA�u�=��w�SK���BH7��CE����;m.��^�&���{iə�0����G[���G�^ $�_�g��Y��~�o�',~6�91��4Ɛ��{�bJ�V
)��H^�;�s�.E��ek�)�$d�,A�Z�	��?�E.��	ńɷ �)Z�eX��g�"����
��M6�^_��G�w�!��/q�[��B�@�Ҝ�oq�Tn}
��0a�J�w_$RL�)���G��O�Vo%�p���<H��[��9%1#X0�^��&�T:��@�\?cO	J<yQ_u���/��t���S�n@���H�	+���/$���Ä��e��7�}�H�ƀ?z/i���7�+ܶ�q�I��z�`� ;}ءS�`O��C�d��{�V�iH���X���NV���W�]p�qd�ϣ.��c<=�@��r�}��G�j8�T�͈�F$V��/5�N��qa�q��[ ��VH��w��a6.�$�i>T�����	��j**�ڮ�q%��4L��)
�u��k51	��Â�RLTj=�G�O�&��A	r��4�ѳ:�6��-0�q.0��)*��U9��_�A��	��~>��T�@��~�~���|�Q?�l�]p�P��_�u��'֖���Cc���f�Aj����N���:�4FBc�,��!�w?���(4xs)�rh�Ȏ(VX~��cv�虛�T���4O[����"ǉs�)y2:��l2��s	fY���W�@�9k8�W_)�x�dL���1��"L���z����"T�f�z�5���pаָ8���Y9}*��c�,�Қ���8�����bU�����oM����FikY(bY��NEjΩ��N,=�:.>��0+���߼U�"x�3���F��p��~~���� ��rɉ�����fNH\eFJf'LXo�K2ˬM9��3>�؂};<��9���f�����B-/�����٨��e	�c��-��E��"���D9#�@���O|�?*�r�/����I �*J����L=����M�x-�.x �����!HY�z9����k��֪,��eY}!(�,��dH�k�P8�gھ�}�O�ӛ(��q˷�IT���:5w��|�_*6r�n�~#���Lc)&�Fع�m�P��ߌ�V�ͭCk���o����k�&����Zj�Z����R����&ɉP�e��.����פ^��d��k�vRq�Q�i2\՞	���z��^��܀B1钷�o��'��c'��+q��b�0����i:p��1������,EB�k2�`�Oǯ)X�!E�2���
[Q;��t4�4��g��c�i%����':��H���	� ����Mp��Ծ����&����Q&T*��cx� C���q��\�>"�:�}������ V����@;y�5p����eA�������dLa�w=G�G:�wõ}p̍e~�����I�w���l�N�xD��O���PMp,�H��������m��)���,Y��C��GG]#x���@Vn_&Zf^�ɦ5��Z<8^4��-ì����ߢ{A���T*ݟ/�l���Co�8�P^bG2�+�D��ҡ�0`����,?xS(k��6���=���0U�>"E;~���Nd��ֲʴ���$���.56�mI1�9�3��Y!�.ήK��T���Z�N�Щ���l�n��]t��O�;8��la �jC�#i�^0���(�k�8���A*�P���%jf�Ȋ��!b<S��0����ͅ��N�~:��(Id�꒧��a>�(��7s��jp�c����w��KG�,<I�ȹލ�W��X��Ƈ?�E���f��nC%�IF~�'p�A ���{�_��˃�1F�`��鳌�Ȝ�nޫ��:��Ƞ~��ʻ��OlG�W��S+���m�w����z��ll@��|C�d�1.e�s�i��+�W�xN)�!d��v�	��}>��@v��#���,D�{�lD��?:6&���$�32����V��Q�KD���Q&20!�ũ�N���7Y�8�P�#���0»�.�l�/Xq��?_��[d.���+������%�-|"���ט��u�B|�
�8�����8ys�1��ӳ-,�nkH����G��i�p�p,���fo(�]v�����(KO�B��ȗ�*�o���@�R'�S�S�n�
�����Df2���"hT���c�n����5��ʳ�xDJx�k~��4��2������\U@2�f�_iF�I���'J��eY�`־�/6�S��;�� /�ך�$�t�cC�q�^�rq�]��nv�>j�����jb�"1�:�e ��f���1��c��`hŜ�Z������on�޶k8~��e���E{�c'����b�+�^?R,џ%�9Ȃ�O("���8n����#K�G-��10'lb�U?�Px)�|z��#U٘�9�Cm}�y|�Ǎo�	1t���=��2-0��<o����4�b�Zosz����� ���9�]bO�
ų2xM�@񙿃}�O�If`~�]�m��+�PnHӍ��QV���V��u�&R�����_t� ��}iX/��f腏�#�7��������/����]�@m�G��
��+9q/�Nϋ�&���e����!�P�!*��r~'@!�|2�r�;�J��eTh|_<��X��
�]~�k+\����,Q������;�!������-r#�m���l��.3m+c������>����~�#��mMw�6u����S���hk'��QHDS���@��"B۟ǖڗj��+�9i!� k�sO��i��1�'U
q�qV_�CjDXb+rxX]ϱ[J��#2��ǃ����" �&a:u�vJjq�)��fs.���u~ gn���.;Lw����\�����1;P����9 .��N��@����v��z�������g������E20��
��ԛf�A���_,�����r;���a��C�lJl�����7�-Ů-�ZMjjP���:D��h�~.��Ԗ��ۗ��4Oᕈp��H�Z�K7�#�V+[�U)[E��lh���[�?W�b�#mZ�=Jm��[�/�o?�H_�"Ri7������߬:�XZO�j�I'��=x
gA�'e(d��"��/�Ϗ�ť[�oY�Qsf���+%��!T[r�����y�<���?\�m��1��Qo��5�� ��#�I5�wY��:�B���_h�F�'�lʉaFK
�[��C���8|	w��ɨ\iN�K#hL�P�?V���
'~sr8��/HpQ����T�=�ߴ�=�L�������n��ө[%P�jQ�,��X�i�T���r��R�йM}��7��Rc��N*�`n͎�@���Ǧ�L_]�&#T�X�`��;Un0�Da`���c�t��6�����Ħ��xg�?�?ⴚ(Rm�D�%��z*z@=�e&U�`�\.(p^M\���P�����v��؍3�6xz�XN(�-��/�=XA�(<��is�0h
>��_�&<�ԃ�5R<������V���5�d��#�X#Jp4;��6ĝR �JX��-)��r�-�%�Ɩ�ycc���D��emF�/�$]f�Ί�}��Y���Tb|�r�8��ߖ^Q�Տ�S��-8�1�I����$�W���be� B�/Z'�鳢��RvmdV�?W����m��L�'^+/֏�k��W�ř����gS���ZI�k�0��v����n?�Δ�}w(ф:a�:�<�6��h<�j|�c�A����v w�̀h)�,�N�]-��3#����J�^�J9��0��ܹrÕ���{+���CiWQz�ԝ! ����M�T�~�g0�Sx�Ii\�b8ZA}?�1#W�Xޫ`����"�'�&G<,�1`��,�p��aH�^Cԯ�
Fkq�c�
EK����{ۇh�X�����<��� ��U/Z{��q�'����y��'�x9�����3��0Š�-e�C`p�h�heP=z�U[NƊ%��Я]��{���g�~@������tÀ���c/�n��>�2���}w���c�t�t`�G�jϞJ�l-ݻ�]�ݪF1�^��Owz�ĭ����+�O������x�&}P˵B���*��?`wG楟���r�Q��Y��k`C�Fz��P�5#��4�d���ǰ�!${�ߞ�u=F[�r�!�Z��.P��ɪ;C�]WO���!��p
t�52ˬ�z+'K�Ha$�Z��֧����}3U��ɇL��b{ح�Ѹ�y�(�c��9fH���c�(l�ؽ��Y��G�B;���.2e����.y�}���5���o�Pq�j9tP݁�@ю.��w)�F�u�Ы��{�6����ν<��^icOjTqAF���b3�l�*��d1�R����j�R7���q������MցN�%H�F��q0�	����L��G&Ru��a���y�����nMB�C5�00�Rg�jLa���\�p������ѿ[T�bC̒��BTu)��2���9(8oQ�j`�ӑlz&��$X|�ē�/^�-[>�o��C-?�V��
O�y�ŕ��`c׈��#��i"�U`&�)��4����'���/��A����}&��q!k��t��p��LSBᶵ�wc�gӃ��&��T�\�MY�FF~�>Rw_.��o�z߫((Trџ����n�Ε�9�*�U)e� z7 ��9Кl�LW]�b$��?js��P�ku���k53&���Z �bX ��&W�|)$�m�G��fQ	zv=v}�9u�dXV�v��a�#3���L���<��SR�xқ�^��% ��I��P� �("�wx�)W h�� ;�j��l���6��&v��Ȉ�g���5�^Q�xF�e-�g���ŕ�<���?BA�V�NfV2�=Ѫ��>
�����DY�5�?Ȗ�Rt��tG0�y�qWL$�x�HS�\�KYO) =�3���r�Z@AVa���٥w1�	m��7(U/>�ۤ������n#+׃]��������(8|�JŒR�O��
�f�sߋr�I��)��
x���+0tj�?�@�0�A�[y&����E?��D��
�%&O�q�^,̩��o����Ú�����Q���Pn����=���~�H��{��ˏ�湆�w�d~η����`<�\KU�/;��R�g��)�":S�X�	����u�|1�>�a5�K���� Tb��2��CC�y�ڵ�|���J���A1� 8�a�����f��h���c��C��D ��_�}DN`�1�i�Qń����tr��k�n�q�������?5cq��8�HWJq\�G����:ѫ&���{6���"�m��P^�C��[}#��OHt:̆����3e���t��6'ȹsq�`l�*S���^�~+�'ۼ��]2k�3C&}y�U��w��X���8�TEiQ�+1���M<q<�Rnry��}�^��r�`,OaJ
����WT���H���+�A�Z5_c谗�ptu�(��sћC!�`ys{������r��Ef%��jւ�76l&�Y�1S������md��d���2g���*ј�?mI�"x譇܍�tZHj�oM2AYN=ρ,(�W��$�_�Tp��uŚ=Z B�N�d����U��XBl����v�)f��1aacHh��w��@kwB#Y;V�8��%�f�ͤ7AdeX�L���	��w$-{��@!I�*E!�+P��#&��m�WM	��Ȫ|��@v�;8�:iO6�/Hz�0�+�}�_��~m=M{����uJ���k����{r�v��i-U/�0���hG�{#;�9�`y�����-��P�8R��<��&_&<[��E�����d��D��8���7�M�M���-�/e�B�a���:x�������G&�=I��K�����R7��Yf�N.8��rY=~�X����c'gp�J�tLt���3��F��K��yo��\a��:�V�<��g���<//˫�(�g�7e�QU+c�0�E2��y�>sG�Dt���=9�]�U�q����1:�T����X*y�X�zʬZ)�!|��hoN�x1u�O�. �ˡ�oTs�̌�r�4�ؔ4\�^���K5�|0嗢��lJ�TЙ�&�"�h���m�}ޭ��C��۳�;?����-�M�y}:�U����-�,��Ж`�x�].^����NPC�e�XD�f�d�g���\i.��)Miv �,�e�^�����3��az%��F�t0�ex�rɁqL�J�������`j0�>�0n�:�	,�4 ���C��o� rW�eߵq7 o{J�(����	���ǈ��h������q �8��ɞ�}���\��Y6����P�O7]�a��z= �ͺG�� �ߋ�Z�[�E�q���T�8�KH�%��!΃=�>�1 /S�ZEr�!�a��*锌��tt�IE?��y�0��w�@�����(��t���֖|�2c�f���[ �]���$���8�XZ|��vffP����������RM���C ��o*�WR����>_��,����'p��BM���II��4Ïn1�@�&+-K�'c�-��Zzk��>���������� ��<���JM�aΚ��5�<� ����vnsR�`N�P�5I�DN��֡Јw��S��I���A�x�,���=n�Y��{�� x'��5\X��ü�V�-i���G��5H0�r�+!(��]s��ST-�%Q*�8^:����O&�ݤ���]�n���C/*M���v�@�ܡ���m٭@5����c���m@���6�b�32UK�vH��Dab	�3��_�@���� 搒9g<����ileǵ��:�n� �Z��*U�w��&��"�%"�(��;!��'e+(6�:�[~y��$�eK��Oh��x�sk'�����]e��&��'Y>/B׃yr!ȤO��(��)9R������15��� K�V�t�K�_a->�����q�e����u'@Er�ͫ�v���g���A�i�����rmm;��h��JyN֊������'�>���!",Ƅ��g�қ��Gl��0�~68و�n8�(����������[#7�hՔx��:� ���ܰ���h#׹5��8
�i|�; \�u�R���eT������������S��*L#�^USf�d/Me�/���UA){��<}���!��a��(o�K;lE:��"xp����$O1sOY�΀����#�v�/u� ��K���2�z�V�.�F\�ݑ�?6�!��Rٟ�Q��+�E���~�G4�?!�:��������n�)*��c
ݣ��mx����B����=��N�'Ua+����[L{P����U~�L�ɘ���ű+���`���J^�d�<df<��	V#@sã(��6�p�{ZM�,}¬^�o�8��@����!�uߛ�ɗ��o�g6�������p�4��H/^�	wvyn�x������M��厯Ϥs��t�[��P�&e�g��^���8>�.b/�T��Lfz�&eU,Q��J�G��j�[7<����CVŖ�b���g���9���x"ۼ�ac%�:���g�3�fl+�)�n����͚c��i���<�MNz����	�^N�72�;==|�{�"��/�hO;4���,� �I`$I?�4~���F#E�ּn��ľ(�~��{�x�!Ly��s�H���z)5k����Q|\��b�����8TZq��3GG�$�LYh<$]A4%0$��N��}������l��5���e�h7��}e0ϐ-{=��-:�n�����+@ء �7�\9�f���8_9�u�±X8���W�HH�V[�E;�ظcX�q�xS�c!3 ���s��?���6�
�ƨ4F��^��&�C� �Ը���}���E�>L,l��v����Ĝh}Ʈ!u}a���̽���a�Q��wV���4*�QAiu1刞�&aժ\𰶕/*�p��*�d��q��;r\�R�I������sc%�ѦM��+[����me��ݘ�X"WEx�-��>������	���������d�G�����ُ�Ψ��3��{Խ�t��_
5��A�iR�P��fz�O�#�ڑ�����m� DP��;��}֟�u�9�",�&z+�p�3)�ɘ�wH9 ��+�Y�xSo5�S7x���z�#�_�Ax�����x�0X.���һ�`�!�b�#�5���Vx�\!�)�kSQ~m�d��U푟}����4n�~���ٻ���d0�s.,P�7�(�Y�ʣ�-
���XS[tpS����K?���/J*a����տL��X�c���4O����Q~J00�8g<�S�\�[��PW}Ǟ����������e{X�Y���J`X ��sV��:�$�`�ˏf牅S?jd���+J�ܰ���r�����D}$nȪn�:�_����ģ`:�8N�M�I$4���wQ����I=�r����O7�9GO_Z8�#pf~bԈWB-K�t,�b�ԑ�?Xv`�w���Cg��42���5����	G��N����d�(PI��ϕ��{�lM��>���#�㼡� �di�ʜ�nd����B}�K_P%3������9~��c�ˁ�(�1��b�+���݉v��;@z´fJ:��R�(��/�-��ݼ����u�~Z���1F>��~}�2��J�.Ю���NS.t�BSl��R���*K�o�'9���c� �n�?�}��T��2#9ci㹓TnVTz�L�����OPV�͚�P����gK�5&������U���݊Ѵ���
"v��'l���2�ܩ�)��-��89l��zI����wQjԵ1�ccbc/E^C��B��/��ȵTQ��ƍ="�J�F�����4���s��9�Z���C׏�b�$�6�T1�V�r���	��U��=�zr8�Z'���B� ���YmZ��/B���Kff�%GRG�w�����KZ�����F�=�PN�n�?K^ͬRI�;b�:����y��e����L{Q���2v�����-[=�3/��p3�-Ue���A:B�vCp܌vfC�hЄ$�KV)�Up�sԕ� ��"gZg+ƴ#�-��q���f7�?U].O)'=�
H^CQ�Xn1��^^ �H=>�#�+�Q=L#ޕ����$� Go��5"�=z87c=��� *�1�C�k=��(b^&�+�����yFg�p���q��=�r4��w�����G�LT�,�d���j<�C�u� <�ە��-���({G��25C� �VDd��X-�mik$ψ���+zA��p�[
�ᗤ����BOM ����#(�Xq�I��~r�C8�R�x�����>���~C8�D�%2����Qτ5 K�\�ޣ���o�=���,�T�-H?�A��7��IsM&%�O�n��{���}p�^τ_{���ʦ0q�oּ�+�w�4��`��Ni���*ƕ��|�G�R�VX9�	Lmk�3R��'�IQ;�N^ r[�V�БK�n9�ib�#�ں��p2xw����r �M϶�˵�E~&k=��l��M�hV�B:�s�Ì]��cbv�)V-�����M�Iv`��48���1���a5ux� 5�����~�- �l�o��V|ӵV�PBa/7�t�� )�׍�.�	��I���̶�E��ϖb�sM,�6�d�rP��o��:�n������ꏤ�7���N���^%�Q$ў�_�����񗌲&�Y����[���%��p�{n"&��r�_I�c�M��b�/4�x��T������j'�[J}֑��sC�݀�xގ E����?�:��n�	Pm���Ʀ32Z��ޙ�<`ײ��!���޴E>[�*�����%��������v��i��,e׊z����|oI;�@n껩��+[ ��x.ޗeҷ��Mͱj�w)!�O<_M�F�⤌�N{D0c�����Kξ�� �L�Y���$�<���q+�	>a~"}��SɆ�,�������D��}ڂEx�͌��+��B�3��Gs�t���C�T�1�j���Ygjbk�m鋏�w|��
R�Uchi��\�ɼI�-�.�A���(�Y�<��6�`;<���BW���}�j�Ы-%���	��8����N��-5�Տ��w*7����fć+t���E��b�&\7xr�@'�W�g�S�p=(s*�$톧� kp�L����Iu��v�=}���=
hwT��-�������<��&���N�:JM%�T�t E�<ֲ �)c <0�
a�9��'iP,�d�q�YY�|��X����U���?<k	*�����8�y��9�d.�]gH��6�`�����k׼����x\�����ڤ��>�c:�f4x�$�\[j��O���q��.�<����R����Y�����ؔ��������H�vFl�dk�:m7j����I����Q�/R w�%���ſ�^�j���:ϫ�F�Z�yf����v|�+ք1�6e̙m�k���=0����bY�z|��c�e����[�s;#�/&��UE�i����`"�v�����<��ݞ�z��n#K�fQ����|ͨ�l1��Eʮ�� =v���%�j���� �Iҽ�W�����2�
Lq@�\�eG���~�5�f�e�����-McӅ����O�m(��s�>�-i6��s�E�!�ڦt�R�	�ʭہ4�s����?y��_1'� ��0w��?�Hyk	k�8�Ь�Pu=!y�v�3e-��e-4��q�Dv=����9
�c�F�Ȼ$�sF�{�;�IW~�f3����u�j��jşT�Etp�[7�����R/��c�P(�����k6:�*&�6}c��UY�-�b.�V�TC����������]Q�C��Ǫ^cŜ�����|��I9���KUG^�gI$��3y�V�zF�DdJؗ;��N�C��������T�ۣ�۝����cA�h ��wc=#w_$�l��\���K��}0�}s�B<ڕl7��g��ԃ��>D�9-$��O��o ��ޚ9�f���[�B�K[~7U,Q�E�n���G�"�G��A����Sf)�?�a .@�W_i=��{�>�ĢՃzX~J,K��0�.���P�D��=	�z.Wp�jHb�2]R�&��J4���3`G|��4{mi}��z��fO��"�A���q��������̴�-:��|�8���}�Q㇕J�Y�T�A߇��+.�SY�굉�J�����������g�m��Wgs���6��^� �ӵ�Пl�6�Tm�Bš��|ER5��,^��`�sm6��8�Ms�N��~�
!��Y�13�ͮy8.���<���%D*)7����&�r��* ����F�Ji'�]�o�ڞ��r� 9�0��I��Q�Wɲx���D=�I���#���"� ކV�@���c���^�<���1|�L��LS((%K1�����])�Pm�#-y�5�v��������w���FkBŻs����1R���e_�B.L�:�U���ʁ�B,+���c�����܇F�9�_�&�zq���v�4�}�rM*�k�B��M+�d s���rs��j�D��#�G:g릉0�����U$�o��*+�Q��6�qR�i��[�OQ����)�Nnp�@s�N�֡��@[�P�l/����o����|�WV��I,>�=��l��"y	�����E�n�_cMH ;KP�V'o�b����'<�Og�� nr1�Q�3Q%{�ʘ��Jp��K�{�F7S�R
EUv(\�@B_D�$:�x�@Ơ9�Ů��ՓYͅb�Oݥ�s�X��rC>ҫ��J��g�b���ܘ&��)���9��)ᆃ\5bt#h;n��V�P��k)?ay�\ğ)B�>ZueH�Bc��9�m�c	��^��K?�Y�;z4���@���개���6��͕z`�U��\�^�����b�D��f�P�%v8 �qI^��a�Z���\RY	aJ�?#�Z�� ��U�)E��̃��Dx�dڢ�:�h�&���G
U�X������ �+cuf0�ՙ��8��;��-�����e�IcB�L�?x�ֺٙ� ����2t'��!q0�֚yV�L�w����R��n�H�	=�@2�w��L�kC�M�k�����5�8�?Y�-�t'�G?��Tș[&��4D{մ.����YƓ��2tkOos�cbgwNJX������mE]�4��'UG�J�ڊ@:��i�Kې2��{�1���~��������1����0߫qM��:[`�+I�^�#�Q�����ɊʾQ��:8�!W>j���ӆ_�K�O��,�9���꨿c��(�q�������	���U`Sj��F
�+���(9����^AH�*�ziz���M�6&��~uy��c�zOަ��쓆�Z���W{E�-�_��tη7�L�PR��% �I7R&>¶\�k�G�K+}�%����-Hl���^��gt��X��+�H�6�X�A��$�:
E!��?����Ġ,�F]�e���{�f:c6��n�hJ��Z��3���T�@lF��a��M�RA^�A,nP#�3�M{$$D��K�Z )��#������{�r��ϨA���p\��]Y<b�FO�|rMu>��n�M*�t��S�2�#�AÆ����0�&��S��d2X&莍����Z,	�nvn/�b`����g���u:�b�5c���jo��k�b�e]�Yc�09�^�n�[��x^?/�)�ۑ����Z�ͨz8<u�)h�.�(��L��F°�]6;cd�'���J�y�p*�6.X��iU�C��O�0^+�/1L>��:aF������SG�1Ǜj��p���jNi]����t�����)0�jt^�9�r@����{QO �on����o���F[�'f��?�zm�!MQ��Y_���/�����������px#uj8Ѡ�Č�������d#�<��,�d
���j���c4��b[v� ��\�A����<�a��aGU��cc�$�ߍ5�T�^�/��P��@�d+a�@UB�>��������dk:���+Y>��D4b��BVG`�:M��bl���6½o�ܻ������`�)� ���ű˫�d��e�tRr{JkW��Oa���E�8o��+2���#�53WiB��}�w��;��m�)y BcJν02��+xx�R*��;@��x8ɕg�V�K^�Wpߙ�jo��+�8$��sV�͘��9(�L�DT�29��]g�2�̯�fU�>���: �6dk:�5� ��������F�#A�H�?'�;q�
�z�U?>���
����CR��T�[�s��K��r����q�e/V(EU+$���~_D� D��v��P:Շ���;�l��K���a�,\����G�\R���9����抱�n���a"��T�㷖�d�xq�;�|U�*�7�iП�ٶP��k��;M��2�E>�f�t�,��V�1���}�s�ab�aR�B��D&ZγD��y�zLdO�8�uG� �&�Ȫ��H�;Nd��������F2q�}[��9��W�������x�EE]e��̾MO�
�����H�G�z����d	
�c�QpuLO2�Qt5�����%|�� � v��`E��zt����Z3��l�	��Ġ����R!�ef��j 7�������9襨�α6حihY�Ε氢�{��kz�)7pY����%�-�K%����:�!�:�y1-H��KˈR�	����O,*x{گ�(���5��'R�Ѩ���nGmW��C㚀����D�%��������"e�2��l�_�J�u�Z*��l���8
�F|a�[��$te�� #)�3_����L9Q!(��{���殐59�J�z`υkjҷ�����(i��
�O��"�2?w�5݆Q�o�T��U3Or�s��[QE���Ø��9o��*�Xmø��b$���izc������ ��B��p�wx0,�Q>ڏ;빢�/�Ɛ�����������N�ɤ��ї`;]�ӬA��"~ޖʨ��׷
�П=�(Kv}CyW�I��z� ��-򧉞�<O@��RE- ݸ"	�~�@����A]F�t��Έ�On���������?;��!T��q�|�[���Q����0<y�+��ͫ2B�?1p��qh�q���,��J��E�Ԩ_�IwT8%��?BE�}��M'��?.}Z[��3�3"q�%k�)�;��)4ы�?Bʔ�Ɇ<�ѫ`f#�8������~��P&�$�2�&�7��?���%��f�����Io>��7��}�:�6r�s�������ǃ �m-I����kig)��vCu�������JU�b65�J[
��̺��w�ܽ�HKg��}bb�����h������u
������ʚ�2>7H^�,�;H­�)�����[v�ZS~|�uh��J/�l��9�-s��xB�:��T���0mg��C��9�<�u��L����P�]$��u�"��
�|�Y�S��N?��;ˍ�����u��7�>	Wb�Cx���{'Bsa��/)�S�Kv�d�Q�T�<l��������3�Ÿ�#B,-�KY�8�4���L0����ܰ"Ԛ�����u��,k�:Z�-��ُb���3r�{ 43�C2��»A�����:�¨��I沃{��e��\\mj�0�������_�.k�69rt�S¯Q"��w��J�L�m#3����i���O�����͑��XcaԤ�z�*�זǙ�Zr�9d-us͌�;U����<G�y+/:{��-��`+��LiE�V�X���SX�CE��o/��3e�Ou=��)�kܲ��>SL�
�=QHmH���4�eg�:���*�tܛy	�w-.Z$W��*��Ks�'�+�)�(��L���4���9ٛbt� ���|� ŐI�
d8]~┆26A������j�ɕ~���%�e'�5��ND�5���J]A/iG�@�lS?1�G�d[싷�u��Z�i"91~�ڹ8n�R}
<�5tIn���㷂%����fVj��U���ww�5�{��/mU�ڙ����GE�K��]�)meNϋ�-��L�+�BͬR��A�C��u�Į5��@$6=�]��X�I�
�[�}=$�)	nntw��P��>4w��K��ozv\���pG@���5,�$��V��D ܒ�ݝ^������Km&��;ũ��Z��Q��l�������W*:�G�������/LY'� �:Wk�
/m����UO�hY������7��(�bX�0����*��wŜ��EPh���Z����4#\��b1��GRS��qFl�k��Z�0�����/p*���Z������� 몳_�2� ��������t'��E�wfc��,�õ6G�y�c��!�oUyVF@�xу�����>��R��	\V�d'��]h���=�kN����p�,ְ̺̈)����G�IA�hUX����_�ȡ�|����jH�T_� O��E1�@����=��&��p��̘��/���f+�1�կ]��D&UJ��0$������ĵ=r�3Y�I=����J_���_V�jR�@ܟb�uQM/Q�x�ow�;l9l�h;C+h�#F��b�ǌ�r�f@�β�7�R�/�=R2�v������*�O��`x�9�4��Q���HQ�&~ʆU�^����:^�eY�r0�7q�� -�g�=�����i�u���)^��Q��K�ʻ��s�#�X�X3mx��3Ͳ����yLYk+��7��z�^��drV9:}k���K�Zb@��b6t	�r�����f#�U���J�3��a(�P�� j�g�)-e.`�:�lE�����f���8�{�T3�>0x<�W�>"�PƊ�����
K��� =��2J�|�e8@Ⱦ������o[��$��~H9��ȑl���e��B�����ۧz�L
f�*՟@�ZDϵi�ˇ�A_���N9D�7)>Ug�;X���6�0�D�K���ݚF�sݛŋ �3%Ҏ�dǌI���Q�9Z�ڇB8�n��� �n=�8� ��%���i"�A�����j	��J�O¬U�}�-��).��Û�>M'�"��%7J"��{���� J�[��L��K&�I�]t��/�N��5���ѕZk�0����پ�!g��SU��c���V���a���+�É�b��⹥�����$4:�!>�(�y��"*�/@�E�5��������efB��	Udm�1q�`�XK&[ǳ�P����$�q9��)6�
9��aqW*뎪�k�%jQ|�䏔�����%�ϋ�Ǚ$yd�j�h�s\�AW���~G)Y��W�u�q���~	h�⑋a!r��ٯԹXnc�t �S��\��M\�Wެ-/�9��%��t:|&�\�� &�k+�R�.�����I��_EF�6 "K%��d�xؽ���5�+��Rk�L�����?��;��)�0]�5��eB�K�O�`�˖��R4��!��Bu� � W�֤2��i�d��U�{B�j�n�e޳���<���]�ha�U�WIN;P��Tj'\`���k`@�X%������@�xe�`E��R=(�"�5U����/���!��j��%���.ŝTR;s�!�H�Ƃ'�O���-eY����]j����_w��#V��S3��goY!��p�[��KU�y�[a�=�aw<���h+���{���� �yK�����ۓ�t���~G�q��&q)��k�V���A����9.�H�sA�z�F�~��=N.T�����<{��z�yX��� g-����)�{m��&$�:�>�A��]I
� ����R{!�cq%�����dň1i��8�U��J;%�S^"J���ʎQ��T� ޹3Jg�uЩ�x��������"؝M�3D�G�N�&�@�ogB��a�t�O��-L'�B؝'�l���8L7���;�MG�p�*TA[7���+�]�,��' ҐP@� ��<dOW����!�6���<um�����TC�.>蜘�`�y|��>���������Ԡ�1�*Z�=�"/o'���I3�甇���%�o�(
�W�h�	hO�P�n'�M�xYaD���4�*���Б'����'����z=Z㛏Җx��H.^��V��S�߳։��>B�L�q9��<FJ��b�Gr�Q��y0M��D)�1�����.�C�fBB�m�����1?XŎ oO����nc��3 R���Ru�EV�)ƞ�g,L��$6T%ђ����鍲����㌃`_�L����2��s���O.�6Mݱ��c�]s �FEE獷�8�k �C�9�I������A����ҹd������D/)���4�qL�G�͒\]b�Y����8��|������YV��|fL�S�76��pPoD�SIo�%aa��_e��Z��p�~�B�����/�ցy����G����@co�V���Vlޠ!�j�*�!�v�z�>�/�&�4!��5�v��P���M�U�ÃVwf��Yx�������9��ƀ�����s\�i�XR�)PBo�E׹�2����͝>�]��2V|Y�d��"�d��3�	6I�:�-���3w����o�!v�kt9wQ^ F�==XS�? j`����J���麅���W�_���&�rTj�,���h ;q\��\�U�5��z"�H�Q�$�[�E�rQa!��yH7�.���~�f@γ�ځ�)��}�vFVӶ�^n^��(fk��#�.�e��v����/��ڨ3F^��T�wXy�ʏ%T@��p�W!�~�_�3�S�1�I7)48T���_��rԵ+��r�b�(Y�f�pc8vƮ�.���RVd���"�N�:����~U��(�������4a��N��d:�n���@��y�S�0�&��)�5+�`�\�W�#:�t�w������ˡ���.ʵ���8?��Ѯ�.�Eh [���<��l�.���e��A�n�ey�XSڶr7�o%���+���[$�#g^RЎUqF3�r�����v~õK�a��>��8��
�fG��@Qn֟���k�Қ�zMt����^��@l�*o)�h@����\����G��y�B�#�a�W�ó��N�ٔ;�Ð��R���={�����9emy�ȋ�C�+�m�>�{��t�j��EG�Y��$|��y���3���Z�I,���I��ѲuT(0l�|#ֽ�A`5ӿ/>�.�F�� A������!ɺ������i-�`�O4�<��L	Tr�Ê��4R�7+�F���{���|R8��c=���Q��2�R@�8�#��H��7B���\����hMh'�����
Dh�#�%#5�O��
�Kx�:�Y�M[d��pD���(�:��l���+ϛ������홌A�-4d��Nׇ��8����<�[��`*��6c@�X��L�Z�dz���v��&�$�l v��C���%P (�c��U��}ͳ���/��<�b (�����Cn�%1Y}ˇE��܃�y��w�L�%{��&��g���3v��B��EϠ���8�?7X:�.y$����%���YM��T�QK����כ�T��p���i�*g�[S2�,0���-1h�NJL�@g�f@���Y(�Z��Q�J�k�?��5��a��ɲ5�ٔ�կ��B�?	n:>�[�
L���:4-�[����x������;݀w�w�
ǙY^i|�sR�� ��
W��/�'�I��c*#,a���ա���Di9�&w���7�����1C���}�0���VD�e�N���@��K��Yf-��i�
�eX��T]�z2�����&O�6�K̰ȹE�J�S4��@���'�8i��k �d7ŉ׫7����$���no�����W;>�!*(W�h ��eN�/���"�xl"\ ����&�s"�5�kC�Q).NK��:�D��@W�������F�,���i��:�|Z�u�]�y��ٰ[�aaYAl���E��s�n����x��<u�r_�ھݯL�&C���N�|�Q�I��;8��W�ŉP�n�-we��:1��-��v.>5�/`�Mͤ7��l����m"^c�������IF~���p+t��
�A�	�{��wS�Q���l	���'!.oW�����vz'�^a�Ѻ�Ddr�����{^���w�9BE����^�D�	[X��B��۩�=�_��>-��[b>�	�|��<��
{��=ۚ�B�
8�IH����(
�Mōu�����X��`�轢='klS�GWcE��8F��S{e#�|ǽhSk�G�A����:�����j-�0�8AV�O\�w�V�����b�w�kH�_�ͥ!�3(�c���~�T> J��W��sB��wO����D,qvTB��ӫ/����r�+��u@��n���k��U]��u�/w�>V����V�$�����=~���H����İ]ͅ���<&^ЎD��@#�r*o��ȁ8����koKi�|D{]~�\�'����\HX3!z�Y�i�*GzZx�6q�E�uz�M) �-y��p7�Հ�=���X�K�D�����yL�2y�H�&�\��z��#J�����xpS�SR�A�
Yi{�AWwy8z'*-��V�Ť%��n*���=�˧=-:�s8c7��T!(g��W՗5���K��!Ь�P�"cW�:U����q���'��С�
�ӫEW��Q�
քj��4�{ռ!�	
!��h�mzEpNe�=m�0ݬf��f�P��kn���	��k�/�Z�$K�k����vA��>قk��Ia��U�½*���Νs[����дa)�N�E\�qL}���=�j8����M���V�P���l�'`�fQJL7~�UE�$=��@��XR0wP���ˉ��)�D�x`�����2
���gƁ�길�[���»� T<�T�/�F!54;�PYOM�Z!;�W�Զa�E��`��B�'`�{��+	Y�´�a��^�6Jk���&�g�9/KA���*�bPͯ)�����A�������>g�m�F��R�{���y���Tá��O_r&CeW/(�.���j��7��{9[\Mug�_��U��<�m ��0�E7p���I��w#�E.�GЖ^���
9t)��V�O$�����W�B�2��X��nt>Ҷ	$C���e�h�^���������YM�T����b�D��D����B���Ț�����g���ũ�؇촭�/6�l�HQ@��}��x�%�6� �[
�U��s~�z�Y�թ��B����D�p��)5��j�o�iz._��������j�E��\>��s�A��]�Q�����z�ų����_���'���Y��}C:�d�|N�4�	}ìTw�0 �����M/Z��JZ�ͱ����HQg8|K�E�3}q[�lS�Xϛ�@��g^�5EQ���2�i���5j��zxl��ٲJ� S����� �<�R���Kx�7�[����^sy�s���P#��q���@?��~��Y�����x�/�킶�L��O';"��4�m�O7�$MN�ן�ሣYG�т�����\o�F����,7B~�^qf;p�dr���S`vHe^���E�z�5]xoO)xW���(@�ǳ��l�̯��Y(w�)�k״'��Y�
g��.��N݊%])�d��Cw�a �r�!WDH:����U����DWP05������ꇝ-�1��Ն�H�=�Y�C��8����-H���֪s��?	?}���M��Γ����T�0I������p2���	�z���檘�����z�c)��M;����w(����f@Mb��ݠ��<�D�C:{�9�⚡���r��)��	�1�y!���4c�_��$g�u�!��-�@K�a"͠����z	�)��
��<?$ ijg�-b�X�;zO~MY��JәR������&�t��;�?]��*_oP)�2��߹�>�$2����>����qO���Al�DY�ɢ6�{�q��_�6P��bk���<�&��lõo=���yI��M�n���lՙϞ�%�N7���2�)H����ٕ`��nx�hb������tH�Ɏi�fBc�Z�cp.Wv8�u˾n�������Vg��b�z��|����י��h���V}(�U�1�	sa�0r�nd�EfHY�o(�j�����_��B�a	V>���PV6䧢�Dz�z_���Ŋ�H]AЏ�Zᦩ}2��Q)�5����mX�|��o���;fުP��..QO��QW+��|]�V��W?�!�i��?<�+�T΄��6����Ã��9)@��񸠫�"t��f���Mo��+aNI :&�
xo�B��ǉ������!�;ԇ�pĻ��8�����������G�&\���YO���n����A<!z�۸�_���i:(��/�I��%���3c;��~i�-��](�V�W݉UC(��F3U*c
��a�E�;O'.��p@
��l�8%�b�ѻ����_��Գ�_�:[&� �(�h�/B��4#��b:C>WQ�{�0=���
�ֹ@8��P^���sH��P4�"�>���J�p��}th���y��)���_�ֶ���q�m��կ�~��1�=2]pH'�N��*��;R%TdA\��C*��4l�}����Q�k�.A��{��-��!�����8ܛ�*i�?�zj<+�!N���c�ܙ�%�S� ��M�x��8V���_�HJ�R�g=��?|��/>p�,.�H��ÁS*t���Ej�H0��@��M3��)��61�>�?4�Lu�E�\Hj�8BHhh���u�
�6�ճ_?�AG~�s�\q�*k�����}E�$�5�z~����E�
^о����^��~�}�d2���[c����+, ��B��EHy�����̭49��׮�wv0�JLz��aU]�����gp0 AU���M9��6rR�?�����ꋻ$�Aq���z�')�pȀ�"�a'٩	C�QU�.ƌ!|�/NV�rvo�7��M��f�H���~t�~T���Mk�%t��F�>@5M]b����8V��o��*�����WXd7B����`k?�'�2Y�S�2�-�5��q���g"師�40!��{x�qޡ����%AQ*������G:D^Y�����!j)��/��� �Ἒ4�Ęޑ�N�GE����|�~i����"�%q(�I��G�^{۔���o�]F���IY}iYu�Z)��O������op�0 Nsp�XA�l:�Ͼl����x��	�H���;�B퍫�\OH���2���c�<�d5����� ��m�8�A�pg��z��0�P���Ћ�,���e9b_�����x���M��J���{�)ns�C
R4��Y��E�K� 6��ԯ۔������ �_��՝>4�f�s��Y�̰�(:02�#���,����T�H����%x�ރ�B���G#Q\��&�+�~��i�H�s����]n��D<2��Qdd$�{H~��S���wIA��Y���D׫8����l�ݯ���yק7��|~F9�G��)�t�p��Ѕ�' $��ۊ+$:!�|�<��|:s���$T��5ԕ5Q�NP9%@;��oS,&9�t�nT�^��:��O�^6�-����/aƫ��Tz~"	@� ��6��N���dJZ��j10�����'���w�D���Qebڃ)�2����{�W�����Ɋ�_��ֱQ Q̪ ��(Ȓ��h�cq=1@i������m��2�k0i��=�Tu���G���V$��a�ޖ�o<'�k��"{�(��EYv8�]*Ɲ��L��]�]�[^S����&º�,X.��������q��w�k�Z��~BE�a��/�����ӦxYsx��;J�G�~ш���W'�#"���kbl���>&UB�}�����X~y�p)�����=yc/�ͥ~��a���A��c�*k�B�Fۊ<��~n4Iͮj�DN�,x�j婯v �G�\�xꈓ(ڟ�`7�V'�A�~�.�R�G�Q���	;ː>��};�:k��@V@��r����a����^ 볢�|k��P=��I�ءv��\�:���J�B���i0���ϒ�ՙ�vXe�O坿"����YJ����N<_�Vnӟ��Ԃ���r��*���R͖�R�S�
x�;�j4Z��5��C_ܶ�ݰ�2P��"�YT��HCRK��&>g��J��s����f���Pߒ%Y+^����2je?�����6�ܛ�4A�`Н�3]�R��GI�38P�u��Y�U+�#&�]iU�ޛ�y�PLe���İ��Sa.��=)|����ևaۓ����rY�ǘ�~Z���l��H'd�,���'ÿ@B��5啍{ �6�,�PS\���[LdI���.�
<4�ɪG��'�7�,�j7Vlƃ,ӱ4y㝙n�>���+>�X�FI��m�(�瓄L�>�/���]��6�`lx=\�~u��05KMG	2�!
]j�q���C��PD ��'�=k��6�������^73OjŻ����2D(u�سT�լݿgrh��`= ���y��1x:\	8"�M^H��_���F������7j�f��7��_`�i�U� F[ЖPU�X	si��P'��a)�~r�ZTR��A�����g��I�<P�#F��.�43V_nb^Zɟ
�W=���CrMږh�i�d+\������@!�xPF8�B�֛���}��>� �/���E9����y�ZB�p�Ik�u5C����� �^����Q�6���qM��n�r�H>eҪ,��(v:tM�1/@Kb� ��<q��W�m �Q�LWd��Rn�K͸X����W�d���lx�$���Y����Lj�R1�H�5Y�}�<�g�:[c��L}M�Z]����
t���~����6�u����̍Ϡ堕v`����M!�!�i�Gd
�3- zfO�M���"�T����x8�7kn/4/�Ք!����zAR�����43�yyO�8ug`{2��������e��Y2�1�� `(�!��p��8;�'�8�'N���j7�GS3���
r��:����C�/W��i²�C�k�z�%�i�ʃd��D��rs:B�o�Lx�hz�q�\���7�O�M'V�yt��.��� +�J�HA(�����0�os��p!�<+:h��i�+:���y���Ɲ��j���d6�_Wxͪ�?�&"�3:���d��S�Ӛ,@3�*���a�%�tZ��-5;���Qy�F���2�C��-{�fG�M� ��#�u7�c/iX#J�q�r(�(R����v�}�0k= �����ϕ�țhYix�T>n��Y��}������F���|!�o:='(�D3DXcE͵Jj��;�}P�V^���HՎ���r��Şa��� ���ha���L(�~�`9Ǯ몷(P��	�����i�����;x�o]���:HL	Q=u4B3Z�\H�8	�8V���6K
JMU��{-�i ��p�˴3�W�Qlo���<�7��@��8w���F$lʄ�,=���2ݩs�x{�0Y��9��Z�J=�Nz�d�M�2OF� O�]�T�>%˚n'0h��:c�)���Y9k͙W6x�d:
��Gz��������/5,�n:�n4o�/�+��h�RHx�����<��2���wޙ��6`5�@�x��S��=�g� ��?3���jUcm:�Qփ��#(W)3�39�WX`�	��h�v��ΉY6���ɔ�`�Zh��c'L�@
� ;!̈��M��?�P
�M��b�R�0�n�op��&η>C|��[Z:מ����͖ђ�)��#c�DB��	tg�;(�⃰��-,�K�R���U5gڕ�\7T�nM���un���?��� �s��b�vĎ�e��:�Z���sb֜|�ʁv� `'��Ih�#�9"�/౯I���kt�H�ݔ�;ೀ=M(�w�C-�J{��p���i\#�0��{�z����R&�����F�)�R�'"z��u��M��-�oZ�-`�&�D�a�V�[��O5��ܒm���-�������gMłx��#��K�'��	ާ�P�Q���IQ�e�ܕw�J�慪yn�r�ҷ*�_tY�(�[u���+��*��d�g����s�--y�A��[��˚��6׏쩈�ᑟ��"��1[�qq��� Ey�\����EG	�R�jn!�����:PW�i��썸���#x>�|���(\�9�?��O1����y{�>�dk�|��p�?YJ�E+^��I\q)!�Sj�GZ��+Z^�+%xx3�à�P9�ڈr���[1���ѐ9�'����ݟ���҇"G�=�H`2��/�wp֗�E�а�ͥdD.B5�����u$��l�A	��nc�sC["�`���ױm��68�ߝO"U��%/^��6�Z0�3�����(�aZ	��p8���V���?\m��n�g-W�s�i����L���
o`"
4 ��Gƒ���Gr&z���M��j$j�?eU�D;�k�H���)�]\��gQ6�*��nx C"��SB���6G�9��[�n/��+���9ɏ��;UY1˸�#M����(v����K���}�<�F;ڍ�zNMôw��|%�D�?"9z��) s�RL��4ċ��Wbt�?�`T�S��$g{u��@�a1(�1�2T�) �p�L���8��r'����Qۧ�����4�?��C8��K�[�}� �~���wH���_�PI�2�ܫ�Ʀd��`�\FF,���PC��T;/�
Q�Q�7�❱�j�Q��r@P�@�LKB8������u��Wf��+mW����(���s��Q�0�b�W�V$@m"�Ȝ�^u�i���@B���{�"�j}4����U�`���X\�u|���'�c^jҴ�;`z|���֯�n����x�O�-�я�|��J���yVᘺ�������jt�10�@3.�Ȃ��k�Κ+f-�G}�����ŭ���a��>����O��u�A�ƼH4EX�6����a�7�����sI_���� x����k�	�wz p��]��ȳ
,n��ZzS/��U0���U4��˛d�3t�k��^�Ī�Vuc ���8l����X�r��rwh��6,�� =�4��o�75����s�rQ�� ���Yq��a���,{�(?h�W��|-�p���,�o���G`�O�S)4B���@��������Riv���Q=I����~}+�̕�)b(b�<�L8=cy�k� �T����р��U�;���.cY�� ��q8G�O{��7&��JM�� �C)����;��m^�j���\�g/�������S,Q5P�ļ��_�g�h�U�p�\B�fW�ۮ�iC�>%cw;��뵓���[8�i*(��m\ ����ɈX4�O
���]f��:/�ک��R-�*�,�c3�RŇJ׊� ��Ē��ynB��4pJ	��%��OO^p��;rA`�0����4:�m��#�Q��7pH���r��a�f�X�z��s�wmYd����iB�BXѫ,J7��l���W��V�Қ��!��I���Q!{���|#S��߬���Xլ�R =c���o_�w5l+�,��-����5c�-�U�#��Xyo�k(��ŷ�f���{zN��L�۠�@Hd���w��Ge�ep6r������G��3m�7Fֻ��n ��FEkMڝ���U�1����!5��������3�k
{J��,���*M(T��)�u%ơ��K���g�\2�Ej�_����)�-	�W1���Xs ��"����	���p�и�a��i�s?���q!ht�T@�t9{�7�t�.8؜��̸L�d��\L[8��B|m�H	� ���Y�Xa�H�V��/�%�+[�{h͟cu�R���r���ȒǮ���,�AMj�8��>o0ͧ-�H9P,�贓������@դ1�'�}mUz혚/(A�,�Ӈ�nu@E��"�^�Ln����Ȑ�_�퀶k�R�rR���툺F�u��	�l��!]8B? ��F�"q
rO���碘^��=I�9���������� : ����xB�~Bg�-����R��jM\a�V_�]����L��|f ��xQ�X�2��&޶�/��@�hhx�u���k���8+��JZ�r��p97��Yր�g��p��D7>��l�k��]�A�5_a�wJ�r΃m2k��qĵ�5�O��-��a@���A9Q�.I��x���Ik�|ց\��g�SP��� ]�"����Y�Zj�w���˛"����
c�뤲'�bI|�(��ډ�M򏹉����@�f�_�a�.ґ�(T/2��W����^����(�{������N���k�t�{F�z<*<�Q(��<q2�c��=�P)�;���X횁�CY�l���[V? ����c�vh=�����N�e|�>UT��P���`8��a
orӐ(�EE�q �_7L�W�g�����ۄ1�������xp��7�~�����})!�N>�,�Kj�d$�>%B)��f"�T�M���)1E�;�D�^��>��J����3���A_��_��=�������tH]Fdj;��0.�D�un�AñJ�]�ç<���z2C�k5־qr�+�������x}����jN�f���2Ki��(���J�5q+�����N�j�ǔ?k�B~���a���|��E�8�L$~����U���l�J0E��j'�`�Qǩ�\��5�*ʜR�6�����I�$��N'��G�e�zUl��, 5��|�"��y��r\(��L����ks'�t%���O�ac<�8Q��|�\6ߪ1���y��?����!�
n�;t�R��殢I�;�.��;`#���E���繢��R��������W�d.Hj�x�]�%�!ԽJX%$;������|��3�O��jƠ��]����ƽ��� �*z宖���90�ad+�����w�Y����P�����*p\y�9�W�ɺư$(F�����V�G�oq@���[V����'0 c�K˵�Yf|B2���h̓��$ϮlfB��We��y�P#RG�&`B�r٘�͇<��k1�V����/��d>�҉��¼%�VݟK�ey���L?09[��6���Y�&�nˍ�j;�$,������9����R4��&�5����\gE��u)�v!]���?�}���R�
�f�e!J�ă7�Z���J!2�OY����~������|��U~ ��v��Wmqmx��Ӿ��A|)gѪ�����3Go�j<4.�&�J&Ԫ���u�I��(B�EUd�M�qYN��6ImI�uX;3K���/��[J1�a�����,�J[S��)�W� 5�X:�l�LW�)&����$��cq�<z�&@ˁGjtǮ� w��+d��>��=a�7�>��q�����2���R*�i��β[=������l�h��N��_�����O9��46%��;�DH�D�"ZJ��grp�����Q�U��C]'�_��]���j����)mZoV���0��O�'�^o����6V5�vq�[���F���X� �eD�o+�7#ժ$�����{Yo�mY[)ȁ "��M�Üm�O��cyR�y��7|ޤB��a��g���U~g�BKaY!w���;�<l�B��K;�S��C���?SXLfsR��p.�6�+_ �v'H+���*�w���#��ܼE��#�|����wH�,�q;���­�_6�17�~�u�S�g19�����P�{�5p�G� �r�~���qB��e�ꭊoS0-�	K�?�b�Eڟ�i�0�Ӹe0�F����o���z�u0�`Ӡ�������«�G����t�5ь��+`�(�=�R"a2�g3384$�\�y=Z5�JϚ���p|��29,v&4��/����HVT{���M��г�wnp8�D�O��4�A�af��������}:J�Lcu���#Uw�y��>C�.��j腦�
��`��wE,Uz3��
5�zav��Ĺ�{��}	0�ݑ��7J5$9~�G��b�uRg�eیW��tu<�yL���^Ѳٿ�aϨ3	�z�TP���5ݷ)�$����~��0�Z��N��*���8ׂ�n���>t��ΥJ#5�1���&,FE�%��Q���ڳMeM��[�x�W+�k_<1 ��h�>��,U�`7��`匴+F�W+"��%��l�_,�ol7$XW�\�:P�7wi���]EG�q�!�PJ#�9v|ځV�y�Z	+޲�q������/���-s�I�A�:�ڤ����9R&��k��7��.6 �G��M� �
�����i�UA�#�������J��@�! �!K�k�Ԍ�#�4�Jhdӆ��\���S�G л�$��]	T%���p�H#�G��Y����-e�����c�잁�o,4��N���[� ��co��.j��`	�!��z��H.(��[�!�j��5gv1N�%m�ֹ~�p��B�ǋְಢ����Ƕ���&��_/R�h$�7+I��)�('/��u�t>�<����K�(s���-�z����agp\����"r3JA_����V��24@�p	��E���Qs��������k�\���r
'
��'(wjհxK�9�L̊=�����r��c�&Nof%X���"�u@twV�T��(�zxW)JHH��h�jٳ)E}|�T���F��ty5e�D�#&��{M��c�
<F�6L]l<��!�r尰-8K	@T�;���o�t�����ӡI�Í���/]�"�Hт��,�W�]������daк����)�<����r�������M��d��݀�ڼ`����?�\�N�/�f�~��#��z�N���v(yr����<�������c�/y
L��/�ݵܘk���x��"�����d���}˥��uy���R鏍��[�T;j�G�"j�%?<��������+���Ǘ(�� .m���zmk��[�8w�yɒ�R������t,�����
�mr�^[�	����A�b�$�D]�r��6��� �+慄F�W�S�锑 Q�O�֖f���vD�o`�U4��'�ZB/�M�8�1����O�i6��d<��p�t�<vbl%'�տ&�sH�5�+�T�usү�aZ����Ņ}��Q�o������1ҕ�|ۆL5��X6�Ac�B���Ge�sdp�q��;�-����B,�l�	\5$���2�J��~8�
_��n9���\T�o��+� J;�7�����(NyC�.Ȥ�'� 0��^ݒ�W�A�1.'�w�Us��KrV�CB9	d_;��)��J��)��/��j�(&A��az�Q�%?�ٿ�zI4�+1�b�
_Y�N�asa'��lk�R��+�Vk˄������8)���AJ����!#$�����+y�_��>8�8q"r��9H�u���d^bQyo罋����4���r���EQ�}�}�~(��bc�p�hw�剚��X9l�	@�v��k�Q���I�La(�g�
���N�)$�$I���v�(�$��#����d�8���Ԝ��rU�	��: ��d,T��"&�f���0�)L��l��*Nm���2��d���m��
�3^mB�P�Q�Y�)5��5S���=v���X����R6!_-�r�/֬b5J�(���2��"]�,�w��[=vѽ�&o5��[/m�TFY��)���m`́�=WP�|�r*��6ii����5f�|��X@��F�6AQ&��b���?�2��Ij������z6�f����.��\[�� 4�T�6�/���'#y5�软��4�u-[/���S&�붏!]z=�ŒzMċr�KfY���h�[�%�=|ڥk���͆��q��R��(ݙ{� ���5��^S>�e\b1t7i��������o��m�	6��H��	�K�/UEW��\		.f�T�����3�aof_�sU?�����c���"���k@�)#^�P�m�_�z���#}��h�"uO���a��;l.�
	%�ȷ�]�w.:�����Vf=F�G�i�����"�ݷ��>}��]��@��}A��c��:@(��ō$�RQ��I[�Qu��(=��o��	���-,��M�0Ȋ�Q@)��|�Q;-)W�k�Lp�}��Ui�n�[�\�E�R6�y�-܁!�Z$60|GH��������X��3i{�o�=��n��D���+#�r�p��]�뻖�P�����%��@���X��v���ڌ���aw+[��.�T��8-aJ7M�3ɲ���xM�g�"y�b�t�H��EN�d��Go�¥�B��D��N�"��V��'7���
/Ԕh��ߦ�;Ep��7͋
���O��f[� -+a��{�M&YM��c�lۂ�<u��!n��?J���V:Δ�	T�9.�BE�V 1e��G��'tڋ&�������c8·��.�b��ⲹvx-X��적��c���)���f%��]��}4	��{�9"ȣg��\x�e2X�'K�����=�>��@O\��q~�8T��A�GǤ0z�r�\*�}y��B���>V��@k4X�vR9��{T�E����}E�1������F�77�pR�z�0��RP�..��[��%�e@��ۿ�����=�0����[/�R���$*�l��<���䋓�5�be�����Xw��Q�<����R��G%���A�:bX���_�2��NHJ{=ض�����޶����/�\T���a3e9�bx��X1���1��$�ɻ?in��$��n]'�
A�8&�5�Sk�K�	ϛ�'g�붡�icU���|Z�l/���7-�d�
�]v�T�}�x$��D=���y�yM�^Y�6��2��J�s�-ګ���=�s�n��,�H<X��K���i�n�hO#� ��
��؛8C������k}�\aɠ��OY��L���~���P��q����QL�b`�w�x���g=��̹}��]&R�-&(��T�适8B.d��7�n+�r�c}�8M0�ߵI�����6�h�9+zt�	&�C�4��:oM��ϨQ�~�B�� �f�y6D5K�� z�m�mzXv�Ys�h�x�� _iB����v	I�YkgQu��l`$��7l�d(-{�8W5�}�4�^��4����%�#��Yl�������yƠXQ�[UMI�[�R@�2�x���9i���[U�ӞVpZڙr�k��y��/�&�Q����Z_c�8pI�'8:cfO�TĘ�%�kn�b+�3���K�z8�W��au�K�*3��t��g�
�<��)Z�a���A�O9�|��P�����lZa����l�r��)
��X�m"?�^dKB��9��掿ۚo�Rm���PįO/~�����uU��:��!8cps���<����̥�hič8��:��h��@����>��ZB(����\�c+o��-���1J��cM��Y��t^1�?u�(᡾:��Ѯ�� �����e9Fj�C34�tw0�$v3�* S-m��<F�r�K)N������8%�_��$7���TH�ˏ@n� .�n�mWu�v&��I�獃��Nb�+Vt涏15Rv9&�Ͽ�wg޳�ӂZ�� ��~��Ӕ��?�IU�+3eˡD'��ٗAu�L{g0���Ђ���je��(��Ά���3n@Y_M��r��7`�p4*��|
,�[rzc�'˂�lZ���%��z@���|h��t��b�)�f��0��#���t��fQ��+���ت�.������1���5��A
�0[S�]���L�p�#� �XQ�"�\���H�&�ߝ���?p�Z�mO�Oכaq�S�;���x��3�Uo!��ܲʦ��ܻ#bD��l
wΟlP&�����W�`�)νa;M�cj�2��'��5Ǻ�+��q��F�,��4!	4�;�!��N�z}/;￭ع�݂A.GS�d��@�>[�xX�kC:�dǕxy��i�|�s�C�/5i <̒���b�3:XK]���ȉ#�e�@�s�G[Wb=���Aޔ9����3V�!	�p�@�V�59Q'��<�2C࡛L���ڼ��^͋�lJ�槼�"z�E\@H|�z������۰��YT\`}�����c�bx���\����l�fq�sv�?h��s�%���V�-�z"��/W�D�`Fd��-�.s�]��.���4�/���>D!�*Ӎ�b�|s�B��ɏ��8Ҟ��6/av%<l|y}�*�$��H��	��~]���^��B�j��8ȁQ=0ƯP�<3Z��m�%���
�	#<U���$2���:P���nnv<����L�ЏsӁg�������E����8����Dw���i�P�۵{2�`@ȷ`h0 ��#?� A��:ym䣾�7=��㹜oϗ̈́m�=��%��*�K!t�t�Z\͙�.U2C�Z�?~�(�ko���[�o�m|��Sғ9�rktV�@?�,���?�/����t�VM�:d95; ��綺\kA3�jg��r����r̐�EG>���a�"
]�:a6/o1^g�v<�$-�������~��|��t�X�ת�ˬ��~�g`]~��ODE����(�� ۙ�.^ ,J� ��CCA�>�:���ꙻ����B�nc�ð�b�S^q�i�n&�H?_Y�|��yO��B�损��X�v�J.s�X#n2�G�d��Ɍ�r$���_tx�|��<2�K(\Z3H�B��c�l,3�Np�̲iI XL*o����j�ˀM\�������pC���	j�J��YRS�t�I��ɨ����)x��������˱�@�t����Wˀ��@���H�G��!��1e��=�tŞ\��	�~h� 9�u��;1�B^e����d�s����*>mM��~���d��y�I��ͣrf���!��1���-X�ڥ>�wt*���$�gKiA�ŕ���Y�j�������Y�	*\GE��^�3�q�ՇpLh[��m�E�*�؊ .u�^�9�=T�L�������#���#�a4%&�\I�D�����W���ϰ�v��Z��.Fh�!��D�8b'pG�
[yu��?�?�.&�5�!�T���?�[+m���\���bus�� �����N�l1M������#^��(a#CМ-�3oV6(h�r��|�&��{�5�HJ�6E�Ĳ��d��`�a,D]�ġx,>B�
ز6c�牛}9Q�lJ�eM0_bv����m-�gO��x�Cl�;b�s���dBe�dؒ���8B�f�Ø~�[�w����G��7�
�fP�D���+9Ne{������ج���?�ɠ�h،�T�5�?�;a�����ڭ�+� �����C�I��'[��x]�.�<3�1�f6BZQ{�aA7
�9�n��ߗe��jc	ҠS�٪6��?N��I&�Y�:��uJ��1Z�b�3|�ӕDU{��
$"�x]�}�4cj�-6W'���?��mŅZl���9i�H)A���?:�A���7���Z,z����H�� 2�" ۶-��|<�]ko%�`N��,5�Q�4�ɿ�(�o�>7NP��>��G��G�	�M��q��`c=r/u�x}_����#� 0�ц2��3���0*�K�s1Q&��GI��+t�҃���������)��I�w��ش���b����L�l:��ag�%~m.FD��'r���Wʼ����kAE�*��lS����W������#<����Ǔ�}���>��R����RV�[X�ϸB��5��6N�2t���G�/~D��R@4��*�v�H�i|��@tV
pk�^wMB>5����T���BL�8l!��>�D�I��k}�u�״D�:�P��*�f{�]{�N&�F�9�޳C��O��<X�7��²�S �;�;Cx/x�W��q䁔��n�m��%m.h}ɿ�d��ާe_�';�pq 2�M%�r���^�x$ݙ�\�9s�#�$Zi`�\I ���ѧHo�n�@�iU�Ѕ�����-�s��p�����(�o>��y�X8kQ@��6�.�ǆ1�����XL�H$]�)���BV܄T�� ./� :�n��|��i(��^&{Ej�p7[��Q{Q%�|�]�����0O������բ=Yk�y�3�İ�����T�5fSz��ɧF;��;;C.���������HT��MB�ޤ]-
u^��i����#M�Z4�m)2�S�V��fF�U��יI�L��@���{~��xo�}�����P�۽cCx
�t����/������t��ĮKfB�ݘ��#	�oXU����J\Ŝ��?W�n�DRb1eE� ;1[�;��δj��Ĩ���@K�Z��"Z��� �	��?���N��{.��&Tl*��K��j~#��}Rg�z|�$Ko��i�yM���|Ms�``U�g��A�o`̊��e���z�i�c�"��.�	.�����(]G5����N��i�FZ�x��A��d,~Q�dz�B�c�p2,y�90>/ ���K��4* ����a9`�KƘ�JG�a��Q$�g!Ϗ&J�����d �]c���!�-�=����P[��3"GFC�F�]5:U�����҆&6�%�i�(��/bDxYs�Soy��:���҇b���cZ"cX��n���L#�ӄ�Wd���_(��p��P㠲~?M���AU�IiT�u��s�{n�����ua�����������~�
��WƱ.|w ���?Tu�$��Wʳy�}�"��R������~��·El�U��Dq�Y�bM|�)MxA*��m�\�[��w%�q���J!��CS]���I��.�����������N+`��z�S��2�*=L�xN'��iI�M���`1»F ���Ȳ �%�E�KQ�>�����:���8��5�S�|M��#�H���Z�⧛8�hU��sD���a5/������2�俜�lk�/�����gFj�)s��.Y��z!I��HD�Ħ��kvM��sy�逍E�;X`��Q�eӧ%�7�jfPa��0�{�
Њ��&X�ve v7S��2ƊY�Qm�=�-+m�j$m�w��A�ƿ��O
O�+7�2Z�����?��ey�g0t����O�O�"�-xYQ j��-8�M�;���c1u<=�6�lU6�����?�럪)0�_ʉ�Y�&�u'[X�߰&Y�D�;���L�����Au�A܋��r3�*ݳ��"-��.*� D�v;��㦢c�.��i�3n��� 7�_~<n������*�G@?r��Ǻ
%�S����0�r�^pnƘ[��������9AC]D�e�:�V�Q���\p��x�5��,�j�?;���Qe�{#X|����5-���+�Δ���ad�ϖ�52��7�\��M_4�>zI���bp���5$�������@� ���(W�x[K�>*Ei.>[����<��
U�g!jFD(-���G�;��Bļ��"�,=�;��L�1ȋJ�o��C���%��n%&����݌�/.�j��A�\���x��*w���o��:
[�%����v3]2f���h�N���E?p�ٰ�'&��Yƾ�Ђշ��7�Tw�5�@H��so^ �.���u?V��1�M_/��<'�3wc@�0�rf&Į��2,' �X�����i1<��Y=�ypڇ�GU2���mʨ2$cZ�^
�{��dm����Lm�=�Y�80���M� �%|S���|��a��ۏ����!s��6qʗ���SdB~e�l���c��sa0�L9�i��Ǧ��MVχ?Pr�՝�z~y�<a�e^
�qG.e�>6@XM�ꪂV|=x/� <�E�Rv�f�%Ln�ذ�0��O�0���@_�q��_���G�	9D�d�md��:
��
O�t |�W��GR�R�i�\QZ�b+���S��bx*��;?8�}/��?�ڜ��"���w������#G�fpI�[��M�a�i�,i;���b`J�M���nS������Ѭ3 U�^������,�B�[CQ/K+���Àveܘ�!E�i�֍���\�:+�����{��n��b���FV9��Y|�1`���a���O�h���	9��a��k�v��*`\�Q������~P&��<�s]��=NϤ*��H!?�5v�>f�*�����]�c���ꭡ�������:�s�,��_0��p�S�2�ߚ���\�Y��t]�g��c�"���Cn���SeY��
sN.���,�s%�r�١����;_�5:Y���}+t�h?ꫨ���e.wNR��,\��
GOu�� �%V�Pw����`y_-���Q��}?_�)��Ա*	1Yg��G��g���|��
CS�XB����I�5�Hd8T�O���>��Ab�ß8qL��<n���.I�2�mv6|����a[�=� �;����!�Hc)Z���E�)�e�(� �y'"2pl#����Xǎc�J�CV�*>���Og����d��z�t��o*U��|L�\�Of47+� �2�G�>�1���!m"6�#A�����|�߉�(_�f�4Ob=�;�5�<���ł�s�	T��k|u�Nj�Wr�v��A��gDD=�c���sg���2����P��V
��2a���;^��>��'�7�P0�?AM��b=s>���&
�%�a?��&c����ĊlA�M�Q���� �o�C����4���h!�h����
{m]㤐R9{EEض���X,����3�ҁ��ɭ�QJqؚ��@_c���� <_�+!||E�v8?YM�TS�"M�M�c�$c9a`�\����<x+~7+��p�g_a���/�{�9�f<C��z��*�;=5�5;؅�h�9�~}�_؝<дI��d��qc��~���M�Ḿ"�|1�}F8I�����������.xc�"5�N�%	3z�r���i<�S��T��q�F���1 ���$Ә��D=
�������ohO3L�O���>k���e��w��%	���dR[L��9��m�y�����+Xv̯��;pA��ވ;��X9p�Ms��zc�b���pqn��(Ӻ1��`��t4��5�\崬�y�1+ dj�*�3��+��y�?ֲ�k�^��%�nr�F;s(l��!J��-tΤ:�y��{y���%%��c�o��qu7���C�7vb�GCόi�@F�$,�z���6Y�d�s@yl��sS`lG�����6�]���u�.��=FsO=Q���2�4��u����tg��z�{����4��em��n�J&w�Y���u�����i�|�S��P����a�c�L�q�
��Ǔ���@qW34�G���@M%�1�����#�ѳ����m߮�l�c�s|���f�4-��z�o���X�{�&��`�{_N�5���8Et��Fԅ%Ŷ[b��Ql�Fd|[�J
���w
8+D�9��yo�o/WB�3��٣C5C���r�Ř̆�.�`���!��%��C�-�W.��`l���m}�M)l�u[������U�T�=�����7�q�s*~����ppI�&�Z.P���f���!s�𜮿��}�!⢇�R:�J3�8���r��Bi���~�)�L��P6�J�Hq��*J�� ���or�]�|�I�U�&�O�x�cT�a�dqI����~V�C�Ynv0J�_H���_w��β=/�L�3����=�ܜh�/΃v#��OTC��f3c�s��5�a��}]d���zWB!F���g�g��@�-��۔���d�w2Ck����@��CM+a�9����
�O����q"��<m+�> ;�UR��VU.�=�7��pz�""J:N(e�@P��Q� GL�(�8N�p2Z�(��?��(�^C�(����^R-��cHk�!�N������%h���cg�e�4��|�����J2{�gx����wSޕ��,%��\51�!�b�����j�@�q�����f����:�I��c	�6V�8$���`	B ��Z�U��F��C�8%���,e�9��-0(��EQ;q��ܬ`�%���?�p���v{<�3F�֣�y����9��4��^�2�w�7�N��s>[E��lX@��PgS���7hׄ0��k�o�cR��ܔ��'W�mfi���Ľ���nk��-U�&�~e�OE���W��[�(�%[M�� �T
�n��<�9th�O:�����"@V��yK�E�+��ئ�UF��"���F��S�@��9��^م�E�&,b��Cv̙�_�Ok���p$Z������{����8����9�ܕ�F-�Y��f]=-E_��.D�g��Y����K��^�������jJ�
]�M*�r���Z�5�ي������fW�3���˽Y]�LM��O	���k��k�-%��w����E6,��o�L=�%�g)�J���B�����%�(D� -��3���Ğ}��U��e�yOM�0(�=����), ��p�`4�Pi�)�_���6�GkJm��K�����&¥'�/�Sa����Z
��?�"	���������<�߱����1���N\������,������6��9���m&������a��� |�D��MB���Ը�����0^��Il�V�F���=�a�,[a.%C�b�e���G?�a����g�	�j��������cQ1��A���^v�����J��&��Aı{ve�x���1pH�U��80��g�(��-�򸡏X&Dxx�˾�-$��Tm�t�j�:�F[,����b���	�X�9�w`�yܣ|���
�L�Q~��Xa�@��uQn��oe2��{p�
��S04))�͋��"�s��@]Ƥ��BF�:A�3Fց�7�Yşb��3=������@*���tj8f�4��cq�o�x����*�o�>tV��.��*��D��e�b�W"W�e��J���L�J�p�*�qF�Ϸ#Z{!{|�S@P)�Ǌ�X�p�^�&41�_�c.H=���$��­����I�Zk<�Hz���Z���MA��2#�����E"��>�8$!jc`|���A���R^��٘o�K�g����8�ry�Ž�4j:2�;���_�~�ʭ����?M^)z�f0��8�X輅�8�,�R*j�o��}ǉ��)�~��dK�F���Jj�c�$�>��� w	-WԺ����L\4��I'v|�U��5�8Pz>���xGch����iB�Y���_��	f��pȫf�$�gُE_y��H�;��E�[hs~�l|�0<GA���}�������Chel���nF�āf�L`��>+��D�فV�d�-v���./@̭���GP=XO)��S�Xǲ��'>B�fH��T�Xh��&~D�ei�Y�mO�H�Վ <��Su|困��i����ig2�"B\w�\X��$O�ɦ0���J�*>����_�o���F����Pf��CLb�1�9\�d)�g��]�]�HhUQ2$	��?�jH�Ʌ�$c���3�Z�7!!$/�q�]�( ��n����h��W�w������>��λ��T��{�áe��oj!03�3��-
6x�	|}~Oߦz�YD��ՒX	˓��L��HP欨c#�=X�O�f}�Ϣ�#уm%�����o��C������Q���9�ym4�D��8	R��y-=I<��m̹�aH�`?]/\5ğAÊ�ܷ���r3Ջ�����2ۜ��JU\�'%��?,Yk�b��i?�G[�U�������%�o,q<_P�J��U��W>��y�:4C�I�i����hQ!y���l�5I�
B���:;`�S���'̦�i��F2X��j삛x��g��%
�^�p�?j�f9�s���=�s"���<�>��'���E$�2k$�^����'����bX��v�=�|E��\��\ w+Vwɇ	��146_�'k���I��b�z�?���UPU�CkL�Me�*�@G� ��):�d��b���&pX2\�$�n��ǒV̈́" 4��V�wS�����@��u܊�1e�juc�DV�2�c͖ۆ�	ᘻ�Az�ɽ���S:ذ�?n*f�Ũl�~�+�W�nZ!�/�NހkE�����D��Z��Bw���d�E�*��쬷ǻ�F�\`ǌ�I��c��{���٦�M��6�ý�/����v��3�k�00��>D�$83v��ʩ:���d����p�-��$'p?�#-�N�EF�����e�Sx��@Z�H&��[�� z�MB��(���O�t<�^[l]N�L'����n��~Bc��t�_��t��jX�Q�w�m5|�l���JL�Q(�4�N8 �[�I�����b�?v�g?�����7
�m�HA������jGQO�2-P]4)�F%���u �k����òA g�棙<f|���4@VX��3�ף�7��e����i�j���Lȧ}������%|L·�5�I��!�ԙ^s�>\���&!lN�"�cb��ie�N�Z[O)�J�DF'Ѝ��K���K��g�� *R�ƁF�\��C3�������GnM����FP��:��b��9v(=)��$3��݌����y�"9/��
��{&��=
=�[��{3�YI4�ƈ���?ov>� }r�0UBv-W��gXY�8x�������h�i���|��R?`r*������Y�ʅ?\l�k6�y��0|�Q@�A��|A!͟Ox�p6��&�)�'��:��e�z�ܛr͔�8������"T�	࢒/���L8�\��-��t Z���[9�N���7�z�M>��9Gk��&a"�vv#�hp�M*���f��4'c��'qU�k����-�;ϕ�
��.�Z�ۧ���)v�y勵�SlN����-S,��;��bb����!2�"�iBV�� �6�_մ��c�%?�Ac�M�Og��c�Y��� �R� )Y��Ϙ�oe���?�z��q�N)R�Y~h3HU���Y9��]�Q-��*6�N1�D꒴�����o^e��A��m���05�J�c�+�cjW����m9��	F&*�U0������!BcX���Cĩ��M�EML���ׄ�Z�)2�[�"	j�[OԶ��"�� ����xcw�4ǿ���.�R��w�n��z�w>����yz�KU6�$�̛Ek~a�I�|'�.	�n�w,�8(2��`^_Mɤ���Nj�9�8����o�^("jW֫4�n���{ԭ�=_�F�l�M��!�Q�ˉʢHo
�L{[r��i��=A����K�ѰV3�r-�b�7�2%_�Y ���m�m�;��K�P	����H��� #��XwuSO
�U���>�ϭ�8��WS�hhx�:��fY����O�u[��n�~�Q��L���_(�E�Wy���'�\�l��%�^��[�^��>���������+���Z2� �%[ዽR�N�oތ��5��Jh�H��$qǶ���&�S���:[F�0�D�d���_Ɨ�J,q��w����x��<f�Od�vO�?���r�8f�6�4����Ģ?tζkf@���3Y��zo���۴}j7o�^�l�Jc�?�}r�=�o27�x�z�.��M� �����.ۈ�x��&'$U�t�cҘ���TT�ו�V��f�����������>]��]��T��B�l@�Ӏ>�mC�̴�ɍ�>O�gYޮ룟�)��15��OϏgA�>t���\���P
&�X���]*���X@�ж�G�`��Y��/G�ٹ*�JZW�[*��3�eZ|/�4�/Xy���P��֒Ӻ��f�+����.��CH?G�AM0�!�OEQ���S��jd0eїVҨ�o�Es ��	�B�Hq�(���J��]�6�����eh{O-#�?\��Ԥ#��o&�B��N�,}��E�2�����f��v�g�h��#�t��_�E����0?���onPa�y��i�6b�H�KE[��01��!b�W�,S�y
�rT�toZ+�e4�	��8Ẕ̌Th��ƕA�c�BN��B^4�w6�>;g��(s������;e	�>�ꎡ�מ$T
U	��<����=rg@��!�2��>n6��� zH�A��2QŊ��`�ȅ�`T���k������)���ᶓE��!zm+�R��F����YvH#��T��{G��O��$�������"[�k�YLv7DG����,`�8�U1Y��\,��<8�������������E}Idv����G���H���S�o�&��J�v�Nߓ9��U?JǞ��u�j#D&�ߵ2��˨�bφ}c�1��|(�\q�>�|v ��5�ɰS�Z#Q�4�l�ס���(���>	z��^�b�Q��j�k�]�g6�L���}67�i�հ�;VOf���;�v�t����̧��z�l"�7�Æ�l_����߄Sr�/������@��	����bf��f�$M�M�6���N�]p�6=[.M��NC���%����X�t�X��2�����Y����\�t	��k��eH�� �pp|~��Jnu|�BX�oJSoz]HBɌ8W&���MGN�T=9D�􂘒�Ч����`IJe�В��z�e�E��[��D��������ˠ�Z3���#3B����M�
��Ty돆Q\�e<����:���u���H�=��\p��Jd QWyȗ��2���bՔMAl����u Rf�q  ���ii�ZrI:0�_�Z��%Yoh�k9��[��5�$�r����5#;���Yy߮:n7��D��X?�>3h*�'s+ٍ�O��m��r�_j���b��p�W�!v��h_0Dh�%G��ܵʮ��Sxz�^^����?�x��l�5]B}�÷��| 3�6��XD:{��ȉ�[�l\�4+2� �����6p��;pƗ����aZQ=H��4拆V��}��$����l�	|��v����������;z�\��⺯YA�dEos�"��U���42�4Ư��ʓ����*�UaD�3I `��s���V��M�X#��]�#���ѕ�����8�2B3����Q�<�m��71�Eq��1�SŶr�9�a&o���sC�i��nvq��R.�B"K[j&0��PF*ći�{s��nZ�FV��o� oz��yL�E���J�~�������W
j�&��d��%��__G��$"3x�r�:-���#,�(����O�	��$�
���C�i��ި-�������Yw���YX!�1�.x@��Cw�ϲ���,�������=�4�>_�K7ʬw�i��_��?���u�2vZe{�I�b�K��G�hί��r�(� B*G�mM|�iMt����q�M���n�"�NB��x-|��!��zLşpYP�MT榦���5-�|x]i|�j�0fw�&Td�J�Li��(i��m�[c�w��TP����wrJ�(���_�3�����t!y��f>��im|��Z-��SZ��;YxM�8���k�n�X~�8�RH����4�k�u�c�L_hP=�ߛv��Enp�>����[�*���}��s�:�*���v5\u���Hĳ@��T�$�l�i:rVi�Ex�&?ښD��Y��㎸�~6�74��������4�XA�n��:�)�:ǐ��k!�>'Y���,�?lPϞ���(l���������\�*+�� �D���̦aί��.CEs��z=<�� tK\��є���ߛ�U�x#��_�����7�(���d`-6���_���N �b��"	�n1L}�U��/�(�)�N-���8��P����xBHLk�}ZWDgv8R�A�����v���e|{�T��Ӏ����l0��
˓���p55扑���U.CT�[P{�Dyb��B"�oa�}�s�:�ܺ�ݳ��V��Ì�p˟q��TBm�`��ǒG-d7r{ lP�p�������=ƻD�W%+�k��"�X�����rem"m��<�v�_�������f�wL3F����^��I"ݧ�H����y�qv3.�6�f	.�+Pd��qweq�i�Ǟ o�o��h��7���� ��F{=8���v��!Ɖ8$I�Y�34# ���(��Oh'2Xr����Q)�.�B�$�+٥K�y�]��ɣ����`��N�N]5´�y���m�,�S6��-�|�j�R�r��"��6��s�&�R_��U�#�.�Hf	PHE��QX���$�	�m��Zg�/�;�SE��N ^�ah�8�H�J�t���c�-ђ0a�H�7S�YS7$�2��2��]X4K�����p�?T���a�f����Bh��bv������A-!V��ٶ���U�`�Φ����`�w�@�I�������$Ð�4�]N���QN��[�n�'r�������x�E�nb���*-��L(��.JNt��)w�Xٓ�{��}���[/ב�5��/#C�F�/�h3*�qA��)��:Fr����;�c�$=�0�(�<�f�x�PC�<{���|pDv�%��ܫSQ��涷����CqL��n5���I_̛l���C�,���;�$]~v�al�M�rܨ���0tTU�3�WU���ڦ�`�0g��:<���/���r	��Mʚ���-��_��,)!��_�4�ۖ�Y:}H��^ş�NFX�������7��Z���z��X��VF�KD,p����]TP߽,��*7<g���y
E�n1�ȡ���A�clb�S4A��� ��9�ެ<�4�^�����U!fȩ�����;�=|�W���J���n���^15�Gsœ'�n��\֣j�g�p���m�t��q_<��sG9�]�/$�>(z��.�f9�r2�xBQ���:&�E��9�Bb��Y�[�:(i]EK>�3?�k%��v�k�J9�K.3p�M]��g�H��I"h������%�Yxc�*^r�STDF)���@��,Ř�W��۹u��L���8�|e�����k�b?ۂg���_�6}����A��ŕk'���u��I>.P7M�a�28"�ͣ�l>P�6�f�:`z����i�L,��\���-O�"t��H6��u�$~_N���M=抇���<���b�,�d-�^BS���11���%ۍq\�,�uR�Kao���ơ
;Բ��I�P�'��yy��jK;��H�b��6�lL�.� ���*���D�I֛V���,� ��k�\R��d�/���l���Y'��/P &�}�%Eo�W�������ح��[�Yo�����5cU��Dv��6ko^2r�A}�l�P��ѳ�p3v凇[z�5�y�xO-�^�y�n�aG ΍&9��~k�ً�&:���cu�Jf�Sd�05r묲�ϳ'\X���nXG`��&2�Iو�=�z됃`~��_����nt�Mx`Lh�Ց�Щ��O
󢶻�^Ld��}o	u��\�����'���4�J�Q̍��)Nt4��-��>�M�r�Hg�3���5W��1�(�g��?�$�dN�0�)k���ׁ�[Y����H�ĥ|L���30ϴ.Ua��i_�>�2�>�.���I���NP�/H��e�4���IW��a�K��	�f�� ��V�i�i!//�)�B|��j�}�����������1!܇3�\fc�{Ed ��H��V�c����� �<���lud�ɻ�����y>Ѷ�Q{wpU�B*�9!g��u�U��C��y�f��>�r40=�X�ȶ:�*����&�{����V��/N�@w����9U��C�ל�MQ�J�Lp��ǩ ޡ��Oe9I_4�&�)�1 H��/�1ԑ�Ѷ���rk�p�����t~����<'��e�t�����s8�=��DX#ٓ˛j��k������)�qЃM3��>��&{�4�'o2=�In�`:"(8F6sq���P7�f�=c���C%=(0�"I�J�z�,��Ebq��`Pߤ�4u
v��^o���kg����h�oɟ\��b���L���V�xJz�P6p8���S�� �Z�ٌ?���%X4Es������h��=H%��:c�<ɜ�����D��`7����ͨ���DP��M��F���nC�_���{
��}���E��)$��8<5C\`�*�C	�Jw����u>��0�X�H��A���fX�t���~@�0>Wk�c��J�H�G�;����$^�dV��b6�qv0�8�T3i��.���y���u���wɹ!�y��Ȃ�v�Ԙ��3�7��/�Dj7��S�W�̯��-�}��+�$w��-':\ͷ�\i�֊a���,���y��M���|"E�^���V6���o�Wy*fl�;��T��T���Q�m�����
�@3J"ޤ��9["N�����W^�۟ţ��C0�/_0F㢕�AB�v!ZĽ�&�4Wk�9��b�I6�p�0|R3	����v�)��hFbL7�)�������	0���H���`/��sr�RWq��������<�HO� �8�u�V)��62�>�W
2;�b�OrI������@���3 o���$ڥs[�^��]��J��l�P��YU��g���nUq�p����������A��P*�Izs��.�4nk��E,�D2���Q�y	v"�'�:Et#}@T0���K�'-\+מ�c���;���u1����ާ���["ex�Vc�߽n���#�h����6��X�6�zy+�H�}˳(Q�L�>�T@n���ԓxSz5iX�5l��"��K�U�uy+�W_�r���ZQ�:��с��7"�W�	,ee�'ri^��MNjZ���_��X]�p��wbI�T��4��dK�E��
O`���N��
Dmq�/-,,ZE�lPC0n�y$��!ā�o�#�Ů�/W[C��	M��@��'rΎ9�g4[B��yX���6���ok솊=	�ť�Qv�?`�ir؝�#N�[șA\�W�]��k΢�v{��J����d�_�+g�\-\߰�<�ax`��N]�t�(�2�5~1�H?��~����*�G]�;T���M }t��X,7$�ٻ�X���)�L�.�4���>�B�N�x8�� ��d  ^�T ~5�ԧ����)�i��/�a���"\nj�%�)ʵF%���$�gBN^��u�u���Wp�#%l%���1v1�*{�a�������cgEmRiE;��(���f�J���𩒼GΚ���
$4���e�y�x��4h����5�O̽ ѣ���R��C���	�9�,|tods�����o��.�%V������Yg�f���L��=�@�0<y��z� ��d8������c3�-/g)sk��J^��P@��h�T�]��!�G�3��.y��.0S(��n0��\��:P�n2"�Ev'ʖ;�s̸V-C��^�O`�~�X*��8��H,M4_$�r{�8�o��{�_��T�G�r5x���8[��O�o-�cL�!gJ��ǢLP������<�A���GԳ8�lM�O�Y���\�ӵ�!����Mߥh�T���3d��ߝ�ÃӖ"de��z�ZV�㐚�������A��a*�I=�-&���
���.v��w��qv��o�$2�L�d�:u��w��śJ�J��ի~[=���)������H��'�i�G�a�d���`��+2�K]ݵ�_�Ui��xԮ4 z�����3���MOw���@��D�R���=���hӅT�X 
�(�=��HG�5��9�8�;MB�i3�^�	��CX���Z?�����p�6����:�+�![�+���0y�K��9��=��|����1A���yD��t���޴�ł�2���711�@�sG�-1�ĺjI��q��%��F6����`�
��d�]Ɔ�VL�0���&g��Ĩ��d�^���f���������y�������:C�G�,�0.iK"ةt�X=�{���iDO�m�k4Z@��E�*���vOy
���i��Ɨ����B���\�A񰫙:6��	���$����_����%l��e���h-K_֯�L�D�$�((���v|�C�X�~�9�>�by$Cڡ���հ/�-b�ƴ��U��l�m�e���
.�/lJ������c��o�xGf��ga�����K2p\d׼n��L��	�؁Љ#Fr ?8�u��#�x��4Z��s_��f�~�7�g��f(���7q�$�5�I�v�-�8L�^%.ۢ�F�����1�|��`�Dg���J���"i
��l����+{���?*��=����u=�Q�p҃�^�!J����v�O������y�nr[ȟ��F6,9��F�����_y�OjѴ�*��\��zz�J��\�	�rV���� ��"1p�Y
������S�S練Y9�6F�{��x���� ��{�]ȫ���2 ����A��_J~ˠ�/�eyD���w�ȷ�*� <?s��PğP�2���?���`�ow3�L�+[�h$��Ty�ص��U&#$�ڭ[~���gc��K�,^�0BL�2m�qώri"w�H���?�B�����I�����j�~�8������	�~[uE�T����׼���+c�;n�;����r�x�3ܱwI�\ym,�`v⒐��8���Ƭg����5�/������uH�𸩏�$�����bYx�0��-���W�PA����-�����Y��˒J5�\��*�M�јX$��h�;tjy�+2%�`c��<�$֠>	�����g����>�bT��Qt��#�xV��J�l�H���!`�t��N@����o� ��⋕^1C�!�������\�&-�KzӼYʟ����%��5?2�vL@���*Q�33U�bM�W^�'�F�z�X8O�n��	W�}_n�����0$��>�ع_���1Xܴ�`����H'a�W%�^�yi�-x('����wd��8S(e3�ba�A�B!�T8|*��
,-7�[���R�D��e��=�	�m-��|Tk�K;Ӟ�Ȟc?��{��2���ҘI"T������t/Uk�d{�o�}۷K�_�Mn:�	�r�ͱ�p�%��Ǳ*��f׏�2ю���9����^(��� �l	���T����kW�p;���ǐ}��80_�����BNXMJ+&b��>��D`4L�W�\�Z5)PwهZ����<�xYv��-X��I"���C��
.ɣ�v������nc��C6��i��X��/U{^&C��ܬ����5�g7��p�Ps�&�W?�R
�t{�Xem��	k�����벫���:��la>Q�yC�>k��<��^̷aըʢ�ύS\���\7�@�Cj^�AwtAf��Oj��!���`M��ӧ��I�׼-x?�U5�[��X	�Fm�L�	I�7Jy,��� �P�wigͅ����K A�L�-` ڬ鷰@Ѻ���y���gk����T�d���'�M[�O.�����o9�f�|�}��G؎t��?:NVZ	��VQ�h/Ұ\$1R��{����@���0m3�=����a�>/��a;�..^~]?��Co�0��r��������!�1UGq 6q Krq�ai��'��4t?u��2���'w�\�"J��G�)����Q0o����>'�I%��R�CV��L�aиNy��]P����|��Z(��.>���K�7紎�c!	��0q��0�&�"H��^G��˼�se&A�XS��u��+���\s@-"�K3b��`����KFb��F_�!�!)��Ϋv����hHT��p~1����3 �:r
�?�G%�e0�X��C^Z�d� %F��-����f�����m�䡛����,����E���BEv�G�,�DN*E{�����x���˧���~���1�$dd�ߢ��  �R�:^�]�FCW�l]�������g��H־�}���l�9V �I7�	�.b��Yж=���&P��?n�����BN/!o��C7mZ?��x��iH��������g��'Ŝ[,��׼�a�``Y��G�"�J���Ӿ�=�D�a�����Jܾ7:��;�ܨ	m[[Q�1��qϰ�i�s�(W�:���pͮa
�4�qb;S�TZZ������㝻Q���{��ӕq���ҁW���g�0���c�~	.���^��<Kf��2ؒ1��i�꾫��/X�Z��)z��lf� ��
�^����mATI�l�I�5��B����;|��mRp#Uɒ�R�D
85E}R4��X�âf?؛�CkS ATڳ֋���{�`��z���[/%���YWᨕ��̺�� �ɘ(��+��dRr�nɜ1^D&Q�~w3���.�;�%����N��!]�a������Y�޳N�:#���L~��\�~l�He�	�cׇ��}����!�P�<�mi�$�y�)*~pmo�6H��5���i@��]��)�����m����K;��L�.4w��M/��	���r�Wr�*}��F�뎰�a�I�?��/����	r�5��M�,�d��m��7J����8כֿ���8��)�ߖ�=O|�G\s,�iu�_��(��#��4xqq�Ҁ2
8df*���!+%��}�|���Q�]Wn�Ws�)��d�ň��\�Kb���6z��fH������ hM��K�u�9?���&��W��_�&c��0��ty_���=��hS	�Ȟ�卷a��E}��񢳋:a1�/R�T��� >�A�KfD\|��y��WÞv��.-�l�nõ9���cBi�91G��Ş�d�^�A���{}�t1�׌<7-���s((����\r�a���u�������o+~F��`����Wx�q�ꯤ`(��rHH����*�^,�G�x��A�{���9�C�5�O}��u7��$�������w2,v�M(�A��9A�����{�e�(��td[a�d
)���q��/�B��]�9� RI����w-�d�q��/$�7yV1S��l�J~�/���bw?�^n�GP��DAË� ;7��� |���8��#PȽgoXV��3�9L)𸔌'��G�u�/Cb?	����R!3�l� !P�s���g��f3Hؿ0ﵨ��y���n�� �P��,�@��M�ES���a�<۷٥�7;�CV+�=�q"&%U�|�?�����	�֡����2�Pr��#�q��ո��HU��]-4ѶV��˱Çg U��ͫB=�q�*��`�W��^��J2Pp��i7�U���0#A�Z?����-RJ�?_��i�n�r pmw�A�?�k��V��Y�MB@j�I+Y�uM��Zx�$�������!_r��w����1�����
�?�)�h�����&��fL<�K\�"C&V��H�cRY�L��Pm<�xw�
��ܶ'��s����-9����ꨟ;��yv��Ie�O��*:8�v$i{�K���2�L�\ L#�����5J&<��ed㢻�إE�,a�`e������憆.�q��hR�xXu��C/`C��:i����e�%�7" E�t���Y�à�:��U�܋�y��챓����BB������4nʏk]'K���R��fH��AE��	lY��18�����b\x֞�3�}�g�M�:UO��o�"�R�t�^�;5� <�,��=���㫬̈����n^d��&y�h���S���-�z�}ҍiTx�����	bG��k���jq,O_�o���b�EK��'�U�y����ur9�!�;�����L���0I����U��Q�Hȉ�u�d,� z���P��

dU��Ӝ��6Ύu Jb�V%
F�E�E���A�'�  �O��'"�R�W�������RY����;� Td6|��mY����]&g�=�d���S�D���������w�/Ua�������٬Ơ��ʈ��`�����U�Xѻ�[��ܘ�G`WR�@N�E¤��ˡ���b�%��g�� ���pŉ��=A�Ju<X�|��f?�b =�I���c���0ܐ�;� o��������p�t�<�fB�+�Ì/���5�_��q.�SW��;j��v��������5��Q�/0~���ˮ�ISDG]t��*Z�vY�`wOԺv�@9�WX�'��܋s�2f�z\^X�>�S|d�b�IDu����ݢ��a��'E���ٗ�����{C^ ��xR���q7���#kVh���a%��'�D��oԠw:��׉�p��.W�+9��nj����g�r�E�'��1�Rs�Nq�n(�Ќ#�R`K�XcKM��LNu@�g�d˝�z+�w4.�yp��[�q,c��\VS�$š���>��ϝ������EG��һt
ы4���Z�#��:擾8��D�\�Dc��\�����[�J0>�\/6�YT�*�eY�W�6�_5�$m
�����h/tPlݬpp��Ǔ�����wO��j
y��r�k��Xpk;X�"�}�V��l�f�ke�S���h���+�]B��~�"�KGl����r��ĭ��:G��W���/)ǰj�]���Ooꖛp�*!24�.MĔ�p���p���
���ls�m�IT��zf��)�=�F\�p7'�_�gW�C�cC$S���(N�y�9�����w��!?P!Rߧ�.ۢ`���z�6~�}�b*JuX>=�����$������9:���V:>Im"d��T���^ALy5�g�}H��!:� vH��+� ��ͺ=�rH?�q.T 7�������*d���iݧrЯ�=	��;I�"�P9x���W�$��O>�8�Js{+��i����$��O�b��!�a�w[ƭ�2���k{���{�R�>n��X�ڛ��3��B����m|�(�fd� �<����఻��)�R�ݍtܴ�^
5D{ZrÒe��i�uD�'�b: ��4c�`P�L��eTK��?t\W�G��1e��M�S�W�!-"En�h��2t��� po����`�����s=�����f�d�^}��_�U��]6�a*ݏ,{���GɄ���PW�A���b+_�"��S۶���=�m%!�{�e
������>�� |v8$Px@Y�%�I��Q���r��t�(�vv�>����` �P�����M��B-V�1��x=�f�Ń�F�"�;�(fT��a�/ʩRMx�`��E��"����6Ͽ�{��Ǌ>�!]8�&�R.��)rL#�4�Ǎ�,F{���!V���y�^D�9W���i[>5��(��)��=��ۄ�I2��X���cE�lh�N��D,��Q��8�g��OMUPA��'�� X�{��;UL�t1�G�� M V��VFf�:LBu�Z�ҿ�6\�ۼI�E�ס "�#KEt`:,(���}iX]Kl���V�]RE_t�%�.�%N�鐆T6�9t��TW#!��������Y��Iߡ`I�qm��˂9�&�=�5�6��m��Vώˇ�/s�{%�dH�&���X<g���@%r9RX
{��xs		�*��sQ]�:f�Oӧw%��}�����%y�E
?�a�%�� k^�Au~���[���d��a�u+G�[]�{ i`x�Q+��C�@MC	3�8��@���5N_��*o��������M-�&�����Q�`�����G� 7~b�VT� N���p��9y��(����+�h�e�q���:е�׉89��÷�PB:N6�!ơb�����l�
������Z�{o˹� v�n�B��T�I�H%�39߬S�Vz����U�l@��dϑ]TI�񑥵{��Ԉp���A+����\�!qO�I�;����^m(���1�XSק��#�%���ԑ�G��7���B�0mc]_6���ͷ��:Eu�I�n�����՛����2�\u�˨����'���q�b�s\���"�Ҟ��� ��9����d��gY��`���զ0�$*f�vt����K$������*�|u%`ɀ +n�����<��)�l���ܧ�����8~0���-��$q�PO�·
:��Y���E~]�W*�A쵦��QxoC�
,W�L�,_[`N�%�헒t8��k$_��QB�m���p\~�S��|���"G+���������	��9�FoŔ��
8����Ы.nhN��C�=F6<i�'�OL�:���n������0$.�^�>K�0�䝿��wک[�V4���'9 ;�����~��\w$�����-�v��iC:�j�!�)8�r޲�m�<�-��}N&�#tX�=��6( ���o�އOt�*���o&��N��u���Vy%��g!V>5hX2S�@�<nR�Ԯ��G���|8;�fwcW� >ʾM�ۯ�����K��d�%K�q4m��nՙ
A��0�fa D���*�|t|�p�~L}��L'�Ш���� �;lY)�}���-��E�q|H9�p�X�<�당jdz_�r�l��������t{�՘Y���]l��Т޺�S��	:b�fVM�V�{���@�Nj�8�;�O!�g<���*3���sgnH/�����&�f`F��6�)�o��)�^u:m+Z8$��.P�ˉ����l�� ��ܤ�f=I��(du���@.�WIJ�B�>禳po|:\��$��a��s΋��Z�A>��[;��sԀ�A!�/�����+r����{��7`�(�= ��< �g��P���UW���jl��e���<�ҷ�n��;'!�Y��o��2�ۖ�{��n&\�F^ņSC��W�z��o�=�p-��p��"��w]:h��0���Q�o�T�8�"��ry��Q��?��*_2}%���÷�"(�][v7�n��Qs�.�~hW~�#g��7L$�L�HS<1���c���u� .66X�)LϢ
�[��*��c!U ԏ Pr�5���`�{FE8t`hsb@/U/i��e�Wz<����7&��t�0����R�#Ϣtf�(���E�|Ȩ�Pg��q���M�]����V�I�;bD���JPw�!����gh���|�x�[���hE�.�%��<Xu�dH\v�?@�x'6�I�V�e�J߀7s;X;x ܏c'T/�awr2����#� p�Ѿ ��"8�A~ Sb�Q�>½{�^!B{P�1��J�>�w3(��*"�u9H7�E�%`7(�_���]Yr�|T�u�L'�����Q*{�pa�0�ᇜ�V'� !~�!>�A�'o�_��j`��d	B�y|��nLR1i��&��j~pU�e`�'��L���Ʈ8��p�E����kY�1�����Єٔ;�O8�t��
wɗ��)��"]Q
4����8g�Z�@*�-�u��.}Q?�5��N���x�a1��t��� ,���gL,�mW��-I�r#[qJ��N�Wg�l\���zOo��)��<P`�u@^���q�a	�[�n�r�g�k�2�^���������3�B�A�B���:	#�����[�@G�'�����3�\��Ay�"nB ,�ep��M��aD̀���%)iH���{����R��Q�a���w�_��>`�+x��U�j��M�ך�J>�g����b}hB��Ȫ?x�lX���"H��X?�ǅ�
����Ѿ���S�����`ύ�[a�$7F�Z1tDM���i��|V��z�r-��[��`$/<$la?��үB����|���x�m�<�q�^�R_���75� �����ȟsd�'8h��B���m6�auњ�6��k�'mln����߲w����,�cb�~� x���[~�cHxZv���?x�;�]VB���gR�L��b&r�mj6��y�<�21�s��<:����藮%1oL��EL�KV)�y��1٥{5w�R�� ��4S�8+������3�f��
�zU�W�Wu\o��}$D�����>*�������OF3�X�%�MY��@%���X6R�L���2���+��?�h<n�]n~:a1������7��.p��P��n�Ty�N%����E�����yOV��,��g	6_@^����3n�-3#��s���� ��1�	�Y]qד�_]���Q[r
	9� 6����~e��H�TK4;p{[ԆQ��6Zn�'r9�_]��5��6�b�I�6���(Wj��~�S�vj�=���%O@M��G�Bsg���4�Gl�K�]X�w;�DQ/Q�k������q�t �TH|�5p&�}��(&G� ޯ���@��Q+�$ܞse�K?U�O�k�z��s7���}�Ԙ=HR�r?�k
���3���"_�/�x�	L�q�EXP<Y�d���4�H�J�"C��[�Ŷ�sK���� �,����+4�i��u�(����q���ڐ*b����̒�����`$�����A`��d�~�V��չ���2!���°VkA�F_��g��0�"q��R��e��yج�r�i��2�K�Wi�W �5sV�M�d�o��+Z�ǟ?�Mg �u�Yv\ab�4�Z��L���9�����B`��m�u��c�(x�Łc���Xg�U��p�8���|���!�R`(���� X/x�[��~�m@SF�ҔV�4����~�K���s�Ne2�M�*�|9�{�
�-�%�*v�.:hɗ��Ŷ�a �����r����>"\����$#M�wp$�o�HzC��r��ͅ
�
Ϙ�j���R��,��дk�:/[W*6����$�s��f!	�{v�U�=�)�p���b6�]��m3��3�co�boH��v[Ê�����N�HZW/����>��9� ��\}#��i��+z��Z�
�;�_��p�xf.�s#n�K�;Jry
FO�~7���vt��FH xG0�c"p���
�+&�Q�g�,�W�/yP?
�M2n����X��	�`տd��'�N�9�`�0N>i�\v����â�,����V���M;Ȟ�W�����.U�0��yAI�E��q�H;گ#u{1�W#��ig��L0��(��6�c^�ܞ)�It�Wq�6{N��m��|c�gĬ���I�5����
POyRN��^���,y�,�Zx���r��䩆��$:!K��4^�)�
�_�z"�1�$c�/��Z������+]��"sbѹָ	���d=\6	�ۯ�[��p����aY?������&�c�-�d�_��n��4��m/���k�!���W~Al�(���5>�M�~�q�oy�/f#G�C������BǼGqt|�!'���q�r�Sv�U<?V4Z�@Ŋ��kY�����{�Z��y;�����n]��<؍�`�u;�ljl7�Z�3�[�z3Qk�?��d�62?x�,�8{`]3H^_
��qydA��~���o�] ���OP�/��rK���#
�%W���uyݑuq����T�D��`���&TE��nÁ{�'���W�=�q%�j�
q��˛G}�B4��(������y�\���f7�w	2v=�\�mh��(����޾M%LI� (��7�5�f�*:��؂��)E��"ߜ,��)�L �E���եMrD�L�&�ڲ	o��Z�V�apllNnᕃO�©Xk�_��y剺�17�gkƚ�MG�Rc��RX73�ge��w>~���6���|���^RW�F�������)�m��|6�F���K
}�[����ry��G�K2}�XA���uo���yB�HS.*�%�� R�Y�5߾ �cH���.�z�����;̃�i��(�m�m˃	t��/T�����$H#ׂѕh��t���]�+jg�8��g��稾Ë����f���V ἐ>��i��U���g|�=upF?`&d��B�f�v��4[^�A��@�D|=$�ِɼ�g��]f��	{�seG�i	ʽ�K� dh���Ò�"�
 Q~�]��So��a*]H���U����F�]���%��Q�N���cCS������jTVU���MU��\W���*n"&rP�E����إ�9(/��S�$�P*ˣ&>+ӏjf9���?�oJ�ï�1�t��<!�5�_)��#�b��U"�e}k-�>z3i�%p��;d�� ,�F� �h����uv���z%9���C�㕰�xݲ�Z�]Q��h�8y���.	�U灅��%������4�yC��+V� J#��60pn�ǎ��D��'�("?��Բ��6�4�
/'�A����4��^���8����Z�=�x���/���46�}YF�M8z��\��1�V�|��JM��9i����N�FI<�����I�R>L��,��<�%H�U�hA�_�Vp��.Rm�ǰ��yKg��-o���;�$e�D=���&���w�W_�lƧ�RY賍���[f=���S�V�m&�	Y=���J)3����s����]�	���z���΅a\{0�I[�WX����t�a�}�
�~������p�6�Y����!=HZ�����rcp��(T?�S�/5 ��2����Y�9�8��˷�lf-@of<zXe�;���;����]Z��#��*wԗ����P8� {?�ӈo��Q�w���_���R��~���ə�i/��������������&1��5R��Z�ٜM`��W��L�hz��˜Cؗ��̇[ᰓ2�H<J��O�U*J>��J�2ʧ�Gp+~g=O�>_�����#��	��'��䥓4�]��U�߁����j�Q��ia�ID�
o�
�˫7�L
NRG�f�'��&^��N�R�!�%�n��#�e�x���{��f��
��	xя��h� ��jt\�F�ߥ~WW��EdufE��L�ޖ+�R"ʞP��_wKH�ր�I?Ӓl���U��y�ʁ�`��?9(=M�Ə�3�>=I����"�^�G(0La=�'�jײ��u~ʭg�kN��}�\uj
>��>��v����Z��D�&\��2J�ɗ$G�#\Q��5�w&�P��g��ts>�>����Uc��F5=���$nGډN��!� `�"���i	P ,�ǑȭP����,��̷S� !����VȐ22��� �q6Ց>���k�cL��9}�"+�d�|O���t�@j���'�P��Ò�\#�v��ۉ�!H�k�hݞ&�p�R d4@���nr��h=^�=Xz�I��O7+F�!2�.gٞ�sVWF�tIz����'��۪�J�f�:�^$/�=5B����V٤lծ�ۢ&���4x��w�'�ir�$��L�W@�z��)��q��K	���7�?y	�b5����B0�|3o�~ʰ;=B;����l恴ngM\b���a&�uD�A�VI���.T[���� ��Wɕ�|+18�+$��j��Ok�I�vꔠ�}��]���uo��v].�A�.��(�gl�9�����׉�zK��+����������Wk���p~���t-=8�l﫤%48�c���:��t���\֯+���zߕa�$>�U\�F���i+lA'��~�^�%8/p�Ԝ�k۠[�Hߞ�a[��ϳN��'�#ۥOg�G�U@-����[��f/H�������c���;[�]����QWyO.�tȉF�5��m~��^uu�F��L��s��7���]D�N4��GY�	'���P� Y�W"��6�Iqˡ���ڵ0���Tf��� �kD��#"뀿Ƙ�`$bD����~*>f������9�����#���졅�D9�ʹ��J��=p�Z��䕮c��`M�X�3o�e/p͖2ɝtz���M���Z�٧��"���Q���._���î�^�|I�q��Q�\�V.nv1"� ����ˑ�eL)GF�ܴw�������ħ���=� ��D&w�����U��#=�YJh�4��x�C����;�I��R�`I�3�0�u�j�\%ٿ�*B���[ܸ&��gÆ>{������H���˥ng-ZS�PN��P��oX(|�4S���:�^3e��Q+�p1��#~%%(�|�y�`
�4C�t���1`"�f9��1�<c﬊�A�
é�K���me��q�R�~���s���ăK�OS�ETq�pieS)��J�A.����Z�6�Ԁ�r�aS/\n����N
�W��1��&�d���ʢ��`8�ׄ�c.�w�{`�B�L�����9v\:��B�zUv��=6%3(F/�{�$��A53�-�)'-L���S�z�ͩ��&r����5@子x���<�9z8�*�w��k���,����A�ξ5�;��x���7d0���H�1\{�T⇢l�	иg���fd�Fs������5�U#�����z�z�����*�7n���)G�����י����~}�5BK/G[��ӔE�UO�d�/aτI��F��s_�*~�H��79� �<#{��
!�9)7���\�	M�-y\�h���p=PAF�<��Ar֘YT�N��M$���=�*#�� ��~�]�w�dp�6u���~�O�o�w����b�m߹ǃ��d_Pu8Ϥ�Dv��t$G��i�ȞH�9�>L5�5o�� ݑ�fYqpô�zu���d��$�E�ǩH�p���S��q:���������I���i���P�((Xzz�����ԸO�B�ޏ�>�HU��ôz���lE�z�1I�_ il�_Ћt�)�p�n�1@ᇷ��5Ҋ����yQ�����<0��3����T���ŷ�3&n�뮁�a~q~�Yv�%ya��lA�9��v꫺I��ܧ�̷͝��^:��-Ro\���A@JJ٥y�oQ*��]yN��C~�$��L#�E�(���5�Ŷݝ/x�U�Z��I�qֲOJ��� n�2$�����1�pm|�(���F�ݴxt��R�MlR���xqᎳ�2��ε�=�� l���H�&����U��9o7}�6"R�9��D�����q�	�9�nb,Vn��ɤ*��kK����o/��,�y1D�3��8��:���I���n|����tcn����4ԷBJ�Lܽ��߶{�{���L[E:S�YQ�6��#���ݩ:\`���nW�*;`Y	M�u* �������K�}�jҘ��I�Y@#��T'^#���*1h����������\��VDN�
�X�?���Tn��uR��oa>��K�V�&CY�+G��Z�fQݮlLl�R�I����D�"$~{g��B��w- !�/�9{�#*�/ ϭ�(�4���JbK�\)c��?9I��:�v>;�Ϭl���`��%��F��_���P�[j�s�S��������K��
D�ö�v_�1��)yz��� &�[�
�V�ڟH��dx����ٵm׆+��e0����~��	@� ����_㿇������ґ����>��ݼ+�x�-
#]�{`"���3K�0��N�xLw��<pa�7L@�5��,��bp�.��QǑ��������U�!>�\ˠM)����/^��&��L��#kW��v����J���q2�:���K�W^w�}e�O�ې:�*LK#�$��郞+�Du}�(Ɋ�7�n�K���b�M\��\��.�⪵!ZC�%�Cw{��x�F ��Õ���p����U�j��@�;TНU�c�����,]���4'��#nK���@������5��=��7��w ��m����L�Ү�*�7"P?q����ZX�'Z|G�u�_�7�%��6���˼O�6m�FR��9s�"�i4�V[�����*�9�u�q�E�)�4t�PU����b\C`
��e��1��A!,8�N����23Dq[�K������HW��]��#t��Tr���r��5I�w��M~$����ڽ�S��?F��C���#(��L�N�0�1#XV^��EZ����6V���[}HȚ���!��m`�?�4�<W:Tb�:��d5�΋h��[*�[��)"���kd�p�7��$�ZAE�+/��|#��ħ�1�d��������X�s�d�I�պͭ��&{R��Ɣ(�<������:m�^�p��r�����>�L8'��5������u#���9F��/��K��z�4,��R�W\��M��A*�h60�?t��Q鳡����@��y��9w�7ırEx�F�����֭u?)�^�|��I `W����8Q�)��j.�e����<%�%˽��ջ|��̺Yur�c,)�Ɨ�d�=�x���PN�xe���� >�
� s�H�ǽ���b�G+l%�ۙ�v�k��s|Z��v��2K+�3���e��OM?g��5�K�P�@
Zu�;K�аXnaj��x��5�i���֐q��t���"��_(�v�y�t�$fM�h�����3::9N>m��)��_{�P�($�Zd������vy�7e��<�W_��w�)ҁ��R�%ssJ���X��3V�V@�6�u+���GC���ɝ���`�qQY/g��&g�"k�'�o���x��[��u+��pa_%��9�,�j�"r��8��j(}���~�s���b�Ҍ��>�y"��'�Y����Y>�:�n�{��ڮK�Y8ht~��z��7�����띚��9�I$�k�(������>2��uϛ`|�]��K�d��Z�WKh��!�OI���+mX3��O�=��������i/�Њ�N
�7̳�[�@1�u{�ܢ�Z	#@kL��;35�V�f,fﮔ��'7��	����.�a�e�(8��2%���� +;j�+�����&C�čU���O;W��ϸ����h���ϑ�VI\��/������bX�<߸�-%ľ���C�'�#(`�k�"�1���f͵��smF�c,�1>�����]�g�ڎo�m�ǿ$x�U��Y��^�<D{�,��a��ɼ�C&zrr���� s�*S臞[և��
6+��%�\�ߦ��)��j�����I$��X�9���@���e
���t�j��T�b'����`���9v1���7�*���յ�앛�����fSG~
��8s��DoI�r��
�i�@
�^��j�� �� O��W[7�D~%`9PY�|T���w���������.|N@gqbgX_��4�i܄aO[V��g4�n0>�ۼY�}��QᔨYF�ŜO�#Q��[)c��.\F[6`6]��s���޳�Lć%���_�%<{�<���(���VKO@��̬�{5{[q�V�6�kW���� ����be�~?Gݑ�}1`���o��������QP7�x��n8Ǌ��	XQ��3˵�����'C�pҍ
�R���C���Q�&Ѝx$+u	9�p���j�Xr��g	wi���|���n�Я�Wp��M�Ӑ�S�'J@ݿi����5��^|����V��\�Q-z>�(��*v�ꔧA!�Mr�pAQ(�����;(�)�	{@|�Q���n��V�}�ߖe9`Hr������ԨGz�3�z��xC�xWI��I �f�E��Etu^�VXYQ���J`=���5�4:	0�ߌh��qX�@+���p�2u�L��a�ԣ�=���CHZ��?;q�d�mG\N���-�j�����_��,E{x)ICn��_T���{��E�SoK^I��s�eqRԮ��s�Y�lC��E�0�B-Cǘ?�h��5;�<z�v�����z�!G?zj�c�s�PdP֙� ������G���>Wʣ�W����0K�fb�����x�2���{����,����m�,� �0󓯠(a�b�Nc(FS���A>/1���1�B�#���{�Z�O���w�v������q�{پ:�������kx�l�ʏ�p9�[��2���6�=0�L� �C5��)��X\���
h��GwK/�\Y�UD������<�
!е����5���&����}��ʀ' �:`?�����a?/��־G��~��8�
���0�YmZsX����f����*ʒ�kU��t�H#�,���T	�c�lUU��Z�nv�8��j�&m�%��Ā�hͱ��,�Dv�W������L��v�Zr�.(\��d��yT��E��[�
 �,T��
	���	Z��NH��M�C�.����VD�M�s~�v�eΖ�I,	��*R����=6����N�������ͣ��.�%kd���X��ƌ��2��Z~���?�K��WfO�ޚC�g�
���0�'�EǺ�/������^�JT#����@:~��s��]��
!�J�+��;Q�7����+���� �5�� �c*����^�,ٓ�N��7:U��]1Bfu��<�M�ǬJv�4�˶�j�|Av�M�M:M{4i�Y�����H�_�pS��nq寪1����vCr�heߤ��_���c5�M"M�Th��t+
��f�\J�O��.(����4��hޏ,"���U��_�I��r��W��y����R�S�^vɉ�mK~�#���QX�L��;6��n��P,�����	8��nA�=%r@�uP��.������ u �W�Z^��q�}�q_��-@ߩث�%������HY������A	T�fBm���h$ˀ[ߑ�NWdm��5���#�;�&!tє_v��t D�����n?Ԍ�v�:�[r�>��80�G[�}�Ip�Х������[�+��~`/���U��G'��W����s,xB夣7��6jd��s�@��Y��(�T4�3���nU�
_� u3ǈ�� �Á��aYw'bS\�z�4�;��3�p�^������wW&
VD��e� �@���U�wӂ6�k�D�>L��	�\LV��6���ɗ�?�T:���"�8<�de��[3X�
A� H)�h>ک���L���.U�O&���Q�qu��pi��~�-��>���.��x��p�Lfh��/�ע������[�ӆ`��d��H�o��>����+t�Ze�<��Mm\��7�ϴ���a�l�|o���{�N���4�/}����Ɍ�74P
;��w�H�������&"�g!PV���dCt~v�']pZ�%p�O�žzv�zy 7
=?&��L��uZY��e����+|��0M@�ޅ�[7B�<o!���ޚ��){=��c�Z�������.Q[	0�c�%8d�9u�P���(fn���#��o��9 �HF��'	���&������q㧵d�33��I�+}�gL�M>����"i٭^�o����e1�Z����HV�J�7EhoQU����,�%��HnEϡj�x�����LI9�}��"�;{�&���q�;˫�C���-Ro8�Bi%�B;x^f��ݵ�{���$��t+r���\�Nթx����<���=7r��A���tٹN�2���WF;p�u�bm�k��Eӄ���խ�J�����C�?���f.�Xdr>Y��s�ѽ��8zõ�h }x��U���6h Di\wjPA�L�I���Ov�,�mָT|��l5Ig���&�����&��'��|]Y��|�N�}f��1���Ⱥrx������v#����d|���仃��1��a�-��D��KF�Y�&�,��龽Ze���ëo���[\��5�:=�ڍb��N .������R�y]�͆��=��O��̪"\;�T֘�L5�؎�1�e`�9��x,��T�3��L�����
�gª����,�c��eB2�ߍ��p���ۊ�iZ㺬6ii�E.&���|�<���AsF�������u݂��Ǘ>0���q1��Cȫ��;qA�i:o���|x,��%���A���f`ɋ%���J��s��(���'	��Z�7�Z·!���O;��М4��"���j�O˙X�B�*��/�@�m�v�w�ͦȦX���ڹ�� ����	Vk A�_kv*���d�m 2����V4�\�?��p".��+��+N��ί��+��3r�Q �J�
:�_�ۼv����8�}��j���5�S��Y���3�Pr~�Y.f�yÏ��^��D�F�]���� s�45�_���ҀC��ݬz������j���H��j<k~�`	U��%��Xt�¢ J�F��'ק"Së:w�a�,m{xs���|���^� LA���;a�][&aol�V�)�B]B����b�ǒ��
j�$��d���<�[}�f����l��U��Uz�rL��#ro&ݖ�jf�C=�e����ncO�h�2��q��Φ9f�?��7'����Ú�e/��oD�P/���S{s�諾����J�X~��i�dl��6�[��՚g�P�0��ʀ�^��G�S��O��VǢ�ͯ3�Y^�#��z�|��'|�ϼTQD!�2���
��1��
㑈�NµĤ�ˊ��2�������Ax��NY�	�p���
�2����Ғ���@�`ظ��2O��$u�S2!��� �ky�3YWȾ�͇ �#���ߨ}�P�a�����^�
--��~���u�^P�YS��dCr>ʦ�m�$d[�^~��٩���$Ty�l��k��\w^��PMT�A.�*ͧ�C�?�k+#�ƿJq������ �ĉTihq�o(HH�L���?ZϾS���l���;P�
k���F{&�H��˲�%����
��'?��H��� �9�S���Z���mh�C�p(!�_B����I&c}�>ZXk�Cb_�j]o$Fq\/<T��<��F�r�)2�P�e�I89¿*�d|�<YSZ��T�2�[Y`N�ÉR����Ђ�7wɊ�k9Tč��i�<�R�uAC��b���$�1׆�:�=�.}J���kw����禦i;�/�d9�ڷ�j��s��)%*�&aD�Jc^�Rx��Q7���_�~��Ҩ�N����Q7����<�>D ; �A�����ssjQ���BY̳j4��y�"�o���;��9߶x滩�3/�Y=�����P-�`r���JPN��[��l��B��DV.~�^���*�G�˹Y����������KN���7���QY��ͻ�̶�h@��]��|D����DN��E�`\B�W	+GG�1Ja�*R&?��G�Ν.�	*��W�\����@�Df=2
������wn>�>���RR>�,�{�p��E�I�m�^���>*�ԀG�:�M���L[$���&�C��o��$�����&��������Å2LB9�Y���R
�eqX����}n4�ľ� ���LN[+�CZ(Y�i��ۦ;�YU(�>�{�ѿ)�:��RçRT���b�,BT������Qd�H*�����$A	��]���I��L�`�TT�
��}�Yj�y��͆�vېH�a��� �g�<�����b}�~�I�*Tn	�2��&���Z�E�����EiM3@�Tp�u%�0��#��Ʈ&׷�U<��,��q� �>�].�Y�?rL�,S����~O=�s�I_���k`7Ur�TCj�/*S�fԙ`��p:�qD�\�Y`3v�oS5EF����t�Bw��Z=څ?.���NFC�c.��L�SϬ�|��a4�JL4�ҩ�5�!�I�ٝ�~'z*�5��Ee���#���5)fu��Z�d�d�ޥ�BOU���j��c��\��k���i;���΃d�fK�MD��!�/Yc��9���b?jF��*�^y˭44Y���So�BS�#8Yܒb���+5gl� ݙo�\*	�̗%����k���V׊���GZ�d�np�S%��Ά�;�i�����:���LwUww�P�B��tRY��<��7����׆��h�8�Q�ky1���mS u�ɀ�Kxo�k����/�
"c@��o�̵{U���E$�C�&Р�u���_����Q��W���6>��-�����t���W��gu�e�i��]\�%����0���k�gث����_�]8`�r�Yy�� Yg<�-Z�fc������_��F��vЇD�%=^k�s�L�PF�U� %��#Σ~ܧrJ	����b|O������$�����b��]�����٘W\v@�l�4op�C�%_�r"�2v
M���LFX3�.5N�f�.c��21|�^v�K!KB]���z�[[���T�$8$
+��B�#�XGj K�(�ş���L_q����mC�
�y�F=�QVHOj�>m�L��Cv
M��+�"��[J�
����p�k�F���Ƶ�B�6w�å��BӼ������)h���c�޽��06T
JM�H2ٹ`o$xK���'V���P>}�]v�9x٨E������G9�W�����1���3�5E����G`I�����8�����=�Gck�Q���?��l��Hs�����Lf�y>�HX�G
�r�<�YX6�C2?�~�����	��v�$ߩ*x�]߽Ĳx(ҭB�5�э䮅�38�>�ſ��J&ǋ�مK�-�̎ QOd�S��D g8�(E��/�G�}=�'~trkkO�(�yeh�����\E.�X�ym��i=u��+��v�/�W��oYwJ��p��r�x�)�IY\B4 �	�fdƊ(�&���`sr�vƗ|U�Z��Z|�{�Nnr�Mx��vLdT�����qBb�e���L"���[� (�A�ݜE���J��b��O1]��{O�����d�>x� l��2z�@�̢/�k�lÁ��)O/�C[k���k��d����|�ګy�"&��oM8*�s*ԿH�'N_x|)�YNY�r=�9<3d����H�'��Q/G��U����|F�V��+���n������:,�oVw�̺XYG��T��k��+F���*.�9;&��8�U˝�"3��.*�z�W�!c�s�M���88�Gv�9�2RG�яF�l���I�g��s�a�+�E������^�e`�/���=��#��Y	~WA��:��ءU��,R�����.@"��5 ��#%C�>���4B+4�N����;q��q]P��N7D�@�&@ހn��ᄯ�hgCW^��S���/i�%*�nJeBK��Cf�^�H}�d��1ym-�(Zm�ܦ�ޑna�w\-����Đ�:i�N�s̰]��e^J?�v��O��S�[��|���1�=�USE�t����o��Q+|��*G}=޿\�c��].�g)�'�(A��d!��kL�ѪA���/[��埇$�-2�L�ٛ��r�s������L�A�5d0� =���	�o��+��.��͢5c��=Z�ٹ��?8P�N�L�l)iH����!���寭��ϙ�<(����Fu_L��X�rB����ט�{]�\ő��.ơ�׫Y��=(�.�1�����0�p�#�1<��ۻ1���pRR��1b=�+E+s�+cL��;\�^�C���)�?�]V]|S�u�N3�B�lp�Nj�f�Nm��x&�w����0]��MMe�R�������-~3O�N�k��j�-c£x��P~o<~�m��*ޅ���Ώ4����Z�C/��揿i���չ>*�[0����V�v���|Ў�q����Q�5fގ��0��.�¤��Su���}�~�rB�͸K��3�!��������w ��%�ha�?MY�u?u��9�^�a�WS��|�Ҟ@΅�/B;4��ɯ^�0G+�l �X�x�)1�S"b��4Q�9��:j��_��J⣡�� [~�ހښ�͸g��[p���+œ�3���*�&3$.Y�)�
���a rI�gb����c���_�-t4(��D���+�cYyH�3�H�t�����EV&��+��͎=�G��6� F�����>;����p�*ď� �^+2Q����ٳ�R�h2E�@�&���ġ ݨ�!��*��%4)�)E����<HLA��qc%T��H6�b+9ezu�C�?�'��u��0����ho.-�j�V/�]ss����Wü�MI׍i�Ow cqR�Tط�3v��]-�Zf�yI���!�g.1��)��lI��;��?nͮ��O��p#8O�Q���q��{X��^�XjE��)�ݧ�!��ne���
�aq���t��tޗ�`�����������_2�v�C�V��O-rAoS �AAd)��U�[P��<�<���ܐ��3���W��������>G_6k+��2�w ���W�N�у�FeW���)����`Q*nf�(�!�sv�_&���W�K�69Aț���T��#WDU̓� �]���a<ʭ�%tt9}X�w��%���z�hW�(��tI�͜���-�1��3�Q�n��O�����n���nU����]�41F҉��'�����2�IU�S���J~&e�N�����(��ɏ~��E~%��")�/j��k}�(��1X�湭!��\F�7��7/]���k}~ڡ>�$u�cNgl�*����rk��3�q�7�d�|c� ��m_�k�d�Kۆ��	I��A?�V4���fT�jH
����y���J#v�S���ږ_���ѿׇ�(��B%������G~�}��E]����͓\� |?:�P����^mگ��.�eO�W/����#�);2@f��Ted���I�����.i$-S����B��aNk�4���B��dh�<�@�v����|d��4Yʦ��u:밥.6E"�ejv�ٖ5����vao��8�����=�LD�1o���&���	��',z
q��kU������S;4A��\T�Xܪ��#TtY}�<���*�g�h��u�c0C��Q�O��1��ĺOh���o��&��9<�g�Y��
9��;��譤AUif�V��Wc�%W"���|�;���h
�zm��\�!_$�:7 U����Úz2�~${���D�Fx22�l�f��鶖���ڪTEo��id{���W����x���԰'D�ܧ��ϱ�E�j�_��8��x����-{0Z�#��&Yʹ�a��o�cS��u
�+�uX����cl2;a�2���/�9��WT�9z8H31�%��?E.@�4�"�;� [�	�G�K���W�8*���� ����dHO~���>�O���ȫD?�1{Z���)�hW�JQq[^M��5�+�=��Y�ϵ�v���ҭ$���}\!=,����[2��EvP��=���/��Ym J�:fCS=�l�!@��OT ?=:�)��.ĕo����k<.p!�u���}�`9�m�0'�ʟ��fn(�ד�������+ć��+�4���ou���-�\���H�|Y����ֺ9�c��W{ε��"^���y�|����w���b��2^�j D!L��OpM�T�3��C�.?	����=������}:H�0������>=�s��6�`��z��Ȗ`y�㴏��9�MG"	K͉�"^$�?\�p;�b��ߧ�q��*v�W����&�r���n���EEyDȀ�d,�	q�7�{k�~Jk-T��jA�W��ab�s�`�_	�Dw�ps���h���E���'�X&��,R#�_�'h����zF1�]µ%�鉯���%�2}�>�lg�������φh�Kuq���J0������h�궍�
�'��5��%>�g������tH4�=�	�Q���;�v1s�h�+8%�	�(gmߧ�9�.����T�>v:n��XC�����:`hY���ڗ}c���*���,�i>5�.^1���� ��䅮�b��)_�*6;w����O8_�ԤkT�	(�*�J��<��H��i�P4��^Qd��\�p;"	��X��Z̱[�'�ߓ���>��->*$�j��UI_!=N:p�>�Q�n״
������f��6�|��nm�Efm�u�c4���*���VJ֓sb&  Oςpl� �"�2L���~pnR�����|І��d4V�N+����&���a���%FQ���Gƞ�
��]�
�K���h�TL���Bk�����<f]B�� ���YG#t@=*٤|�\ox�=oL�x�}�lʥQt��i�*I~=�VZ^�>��Gyf37�F��p�c!J5��Z��+wh�5�a������� c��<���Ҙ��
Ss���S.�Q���E`B�^r���u�|V�c��܈D$/hSr�]-�8���!��^BR���TleZ�vA�f)W8V>5��^`�����	������g깒o�e,]�GY�	���.ֲ�'����.x+Z$�uh/����"�_4����Z�k���z���0��p.V��J&��P22�<�m����	�����1E�۴�n$�����
)%�<tot_F뾴�4XR��0ZCz�� �����%`��>aj�Fń����>��kͽi��.Y/�,��n������e'����-a����y�Y?0���eh�Mz�1�űA�h�O�߆<���5Ei1JBdK#����
 �a��As%�N�*��~�l���о?H�?U���x�K�;g�gw+2��W�g��,�pO�"���A��_bp�k��;~f�A�b��$чq�_O�~��/��e��6y?�kV@���G5�B*�������f�~|���Yl�<����J\�m�sг��&�԰g��&!:��r
g�{jڡ�v6���3%ŵ�'��������N�G~���Z_�/R0d�le�����:���X�������q����ֵ�B�1y�w���X�|"U:b�-4�'�ݵӺ���ɻp�$�c�L=�g�5/�v����g��.t�c�~[K�����ͫS��%�3Dc2�w��`l���ޤL(*]�״ 	EKA��e����^�<��$
V��)ժUF����ٶ`3�x�0u���֐��D��|��s���w쑧I��O☧(�5Z�O��bvxӗ�b�)����@�K��l�Y�=�����nPb�3Zv�!k������	��c[�Er֜���Z�R��߿����?V��>�i�1��'��%<�e�J|�)4
��m\���$��U�X��)#��oT	��Yf����!Ѷ3צ$�)n(	ô���Z�Wx�&�bp9L����	!E����
+%d_�HK�d[#�ӉYn���c2����1l�l��ڈ _����N~���34BsM��LJ tVRi�H[����b��z�4��)�Z-ش���R��y����bF?m�!o�\$3��K�4|X_�$C����x���@C��5�/���yWؘca-%�&���es�fdO��"��{��xnI��W �i+]BS�62���e���_����c�Or��?��g��H�os��FZhW���)㍴	F�a{?�cѺ|�U��0�D��-z_��ZP�L���od;g���mƮ>f�Ѭ���(�Wى;2)��F;<�j� ���.�#ư�C)�s/��mK��:������e�/����\o?0꣧9n6���U��76t�s('����n'J����ҍ)E�c�ǉCgGh����e2��Ғ��֯��`����`��Ҵ.'��/���G�Kя�qj/�\9���ñ�������H��n �U�I��iPhS�\�iQ��+q�۠�>"P�Qٗ���f�+�*t��c݌[��mC�ˏ���WXT���ua{n�I����o^׈�[iT�i	�+K�t��ɦXG�/�~`=g!2}U$�J�ß��<�H�`ܖ�b������mXC�����-�`=Lz�	�y��3�zf��)�����aF&F� ~�f1�"��78O>e���ⰼ��j�{�䮮[��
���\CR�#TWJ�̀��fn��4���0�lK�\/}�[́�(p=��8>.;ƌ�s�w���:���ra��j;�A&�Ќ.0m��%�	��)3�5fj'���m���S���Sr�b�@����%��dC-s��M͞d �&x�}H�Vʂh9����z�iB�0\9��E~?��"�l�+s��R�2�D���BߕmQ�{,e>��E)[���Y�	p��P4yB��~��t;.������B_�`������q���o.Fo{u�u��U~2LS�9��(�����txR�uߒo�2o�A@ٖ(��{En̓�$�-R�j��ʷ��6��a���ވ�W�L�U��M�&F�{�莥rZ�E�/Zt��������PM��Hj&{? �=�� (�?�r��T�"��˦���DOR���e�|�<�ި,N�ƭ��6̦��r2V�?h�51|��j)�q����W��.�M_0��V�����1�'�`-z�0��^�6O�f���i����@!H�W!rщH��;��v��,�qo��RSbo���Y]�o1N+O+妋/��2�$[��tG�9B$Z@�'ڥ��/��oQ|�ؙ|�9I�*6�3�B�\A�� ���~5>KޠH6�J��pi�^mG����=� c0�J���G�?������gs˄����.
i/�u��n~B�K�ՅZ�?n3Tqk��8ßӇ�;���u�02AM�ߩcUH�Yv�R���q�qN�LP���Y'M"��M< Xj����;f���!J ���s����C�UtmE&���8`Q	 Na�amR+�j�6����[�)�9�tm���j���r��)V��(��j� �0����O=�q ?=�ٹ[.ڍ����s������˞�w�4O�q��y��i˴y�$�O�"� R�� �J��qu�����z��ަ<�p(��O!8�wtΩ��(��#�M�M?�f�=���V��R$0r�j�O96�0Fݥ�[h��#�%���6\Z?V��yuM�B��قA�mt\G5E|N�"����_if(:��1l��m�;k�B�x��yT�WW7��AȵN�����Y��\��O��T�X�Xg�h	��3�߶t��,�l�_aH7�3��N{�e���ԐS�fܻ.w���4)'?�����:�]��Y�����+��zmeTn9������BgI�a7͝&_$|�R��|��k@}g*C�u�<C�u���BY�:��	�31>xw��QO|y8v3�s��n�۷\d.�H�$��ͤņ2�9���cG}���F�<a��l���Y��?f r˧�`j}��=�F����3���t���͕L�!�2��?:)�7��� W��tG8��զ��FL�~8e~7��Bi��U� �7�ݾSG�O��o�
�L���Rc8�����U��,����<雨��^'��E�m����
�&Xb�J��̀�"كo��P�:'�o���{�|}$r������`�#-BӢѢK؍�GW�uZĸzc8X Q�"I�O6��v5��T9*3���A]�p`}�.�H��^h�st��q���k�����ɚW'~㈆�xx��%q��K��jj뺬Ѻ*U�T�H-] B)�m_��U���;��,��tȎ�&�z�t{\�*�)�x�O�<bm�C+�h�5�����p��)�����1��C�}�>�	��T��?�f�Jt�3@�SƔ�:��7�HM�*��4�5%Y�J~���q��~B>0We�mŽ��L� DkA�n-=����5;5�5�l7;G�:<!P±w��x[|�����9�gL<Z���A|��bڭ�a��3�n�1vGa��A����HN�k������J�= N�æ$�$��?�Gxk�*+K.J:�n�>��lAh��	cvΒ�������_̡�©Nm/yoz�}��]�E���v��n:�{8`~KA���N?��}���/�Za� ���>�Z�������]T�)�z�7�ըs�&*=�ݺ�G�r0h��	H�����ի�c��$h�G������Lltv8�^e�%6}���4ad�;��6@���zj���{/݅�T>u�磮7tNLTH9eI����_�������o�Q��)��l�#P��/\t+���\��r�z�Cr��\\�YjƤ�E��V- >B��!�]��*���}�ҹo���Ŗ��Ҷ��|��ɡo]E/W?0�Ҹt��w��-�ccf��.�Ԛ�ZN�%���Fr6��J�z�~�5�:�T߮Ps��ٙ�c ��:�x@�(�"牟#�q+�pO��ӵV.�Y�T��5;S�Z?�W�֟M5bL��r$�#N��9�;b�;���O6�@9;~�6\��=� ��2 ����+uߝ�Tm���4��*vq��X����*<C�9i�u
�����������-ȡU5#���8�Y������^���:3-� <����Rxz� 10�I5j��t:�7� o���M.$�R&@����apJ�Ipn�����C�Ex��^L�+�WN�yR��T�,b�#]Ʈ=�3O�0k�AOaͦr�w�BY /f���W�Ɂ��d�����r�7a��'[[^�����F �y0���V�����S�W��]�B�8&�����7a�lP��`�I� `w��F�'�5JJ 1y��#Ԕ��9�G�n)p�|�Ql��L�3p��*<'z,�MUo4U'�[��-} a�G}?�x���a��f��l�q1�ۊ�T S!(s��5��J�5$��%M���ӃH�E��"C���F˩���D�8��`_(��5�J|A�hZQ�(��%��i4�b�R��)����aM�+�IR���|x��իF4[֡���{bo5��	�8FJ�!�FxS%��%�8��*,��3���cm��eQ2��
7v��FE~
�P�v	؏��2}����p%fLܸ>� yM��2^ꪯ��1n
B��jՀ��7=��[����F�� z�����Ϙ>���G����~9�V�٠037.��|80#]}��t��j}�!��&]�*t���)���^�	���G{�1o��������픫�Ȥ�������;ӧ�r�Щ(���y���S��k�1�L�/ |�]^)i�VO�����/2�;_]�*�j�'hA��#�n�p�3�5��L3F�c��1v'D:M�Os�����t��C��A��8�>�]�r�����~�Hz�:�g���S��!@\Y.��T ����B N����R\���5&�kOi.��M'��L�-�Y�d��]~�;i4-[��P�=�/~<:��LYnřp�CǉW &x�Uæ.��N���[�z#Y��%i�юϛ5��1��qϩ �j����xR�LN�z^tTt&��9+����� 4�{e-��Y�2����U$@F�vW��mA�o/���t�m��R�g#���sh���t��(�[���m��Nr�f�����9~����Y�p�d%eE�zT������衍�{���R/��E'���$Z�T'������*�J����L�G�P/H��?�ܺ�i�^��fG���Sz	��'�\��rA�/Q �����!_Im�8ҍ�o%�?C+@�\�Ӆ$��k�f\�X���쇳)N2W�(�]ٯw�s#�����J����S�Ԃ�o-�j,�APkSau�kՑ)=��.nD�>�8����� [V�3ӤM��
� WR�����t&G�3YE\4�5�O{"C&�b�[��Ã"����5�@��{�҇6�n'��JV������5qB���$y��Jz$�eTaA��J��nυ|`�W$xi��vS	�w�xjO��nFÖq�<,��Q$���ĺ}i��7&\G�.U��,�����E��5�݆�!o/p�˘�%�C�9�~u�7�[�n^Nu��&D�pTk�Ҧ��L�l���M��X��hGu���U=��e���Ģ���p��H5I�4��pU�`���Y��js)fg�#ʏ���sB|��1�c�����Į[�xE�B�⾪���Eq���L&S!Z��e���apj�[�r���$�O����Fo[ϗ1���� ���,�_!�bz�_�r[�늾���{�iŊuR\+j�j\Hۯ�eG������[EL�Y�D���H���_�L�	�����?��uR�(�Ez�JCq?	]7yz�A�[�)N�� Ϣ9R��NlHZ�2����s9�Yw>�&*d�	�P?n`1p�4p�n��sWBcY0��߆�6��n����X⍌����<~L­��~��[��ƾ�K�̨x��J���}���d8;�hg�����گ&5D�:(���f�ޑ���J|�0��[��f�Yk�8�  �6��{�K���-���AяwQA#��.�ȷ�Ws�A�p��tfT�U�gG�}��ɸavy�W�
/gۅ������\UJ�X��$K�	�)x�Zp�}/T\x�5ơȱ9��&����?��5K�v����C�(���FrO��!�ʶ֝�w�ZGKpN$��nD������5q��=v��g��z6߸��V��Z�乭�ċ���۞sz9���oO�s�n��#ruL=�&�f|k6C�qx$Wj9D�=�nl[>' ���	�O��P��c1��R�-Lm�-i��L�ps4Uz<�k�D�L�0�'}��7�p|�N�~Tn?����L^��vS���h��(�����6�,hP4K�P��!S.�4�@Eno��X��TĿY0E�T4�6�Y	BM�� l�XJ�¬�I��Ux���������pF��_�u��J�Q�}R��qQK ip��޳�B�oG<!gG�]�����t��1�F�x-1�����l�*��n�[��!Is0�f��!9�@n����0�/K�x���a����^�N�}�I3����N1a��!��T���@�S�Յ�rv���A�"�,t�5����Ū�JA����~�j'��J�[���Y�!z��um�嘪��~�����}
_2ey*9���͚��M��x�P��nyO8���Q�/�l�������?;�J'�a{�t������R�[�R�4xb�vT�Ȟ��`�쬽5�z�#s\S_�t#c�O|�B���3�����*�'[w�3��t����5�V��$v1@��}5Lj��hr�$d(�(r��7<.�7�w�R���{�H�Z�������mi�k��VM�n�\2�-����`��w�B�F��(�
��suv\C2�_1�iI0�y�¦Xv)���9��O��`m���&����	���Ϥ��RO���-�vCP���>s��z�a���D6�<�w\O�-�u%�C��T[��1=-� {�`�dO%��̟��Q�8�#K�l�0,Zk�"/�{ 7p(���<���"�`8�D���!��ռ�)��^$��!(�@Yœ
a���� D�_�3�kA��Q���.�t�]/4Tf��}*�I���KpYڸbY�ۨxG�� :�b"V�u��:o�ƶE"r��7�v֗�T�������X�0X�3�5S�B]��{�>��H������
�ՠ)L���B�F(��6�z6�V8_�d~;
�l�jA��?$@T-��m�g!�����L��eu�\чz��֟)�4c12��u&T��®�|_5J)Y�:�i��f"a潫��CE�%�:(|rc>���sg%A��e{�񥲖Z��<ā<l��,)����k�f�}YS�L U��p�'�Dv.d� �ỿ����xP�Q2(	�9{�	����&�e�|�i�c��	\n�e��Y�S���傁�6�)W��un�~���k�p����kҮ��>��ӗ]���}������x<�VX�n�%	[��xi��jR�#BQ�݇6��Oj��wi=�Ĉ�m��b���xeV�Q`g��)�#�/��x]+�x4��񅻧�pz��~�9�0<w'yI{��(�,Z�;6Č.8;Aw��@G����y/�1(�<Q�~���GnM��-H�@*R��`c�C���!X��?�oCZ�;��#a)S�{wX�}roߚM?G��ݾ%�w:r�p-�������I�`�Z������t9b 8���/v�\��2�T�8Lh9�9TH��,��F�l���/aT��Ȉ
�@�7sY��Ոr���&o���*H����H��ʨ�����$�xc���?�At��)�CE��Ǡx �A�����!�%��#��7�Ŋ?Ԯ���n�����r���GQ�����"��H�sO>B��	��H�TmO�l�UBMV��F�%�8<��Ȭݍcs��N��?���W� ]w�Pj+c���`�O {���Ǥ]It.�p�ݟ{�m��(��"s@�aGX���� �����. g�0@P=:�U����]�A�͹Q�e��;� ��P��\���x��>�9����S�4*���Rmv Xѽ�~��G�l��+]�_0�)�M��6!	I_g�Y��O�ǧ��>��j*&Ҭ�ӵO��
���������;{�*2�����wB[mrv���=�e.��O9#��0�!!�3S��G �=}��: �H �?�6�Yh���+O�=i��pq֤�Sۢ��pR;w�Η/`��i�^�@x�z_'Ԑ.�@V���2��}l�ssOao�����x�,��_��aŬ�ՠ���9�{�V]&��n��S���gD��ǅ�� �*�|R���x�.or5Eo\�dp�Z�i��h�	�����/d����<�D�r5b���l�
�Cݒ�8�{�eă.:������)"�Q3�Q�$"V��BiMЦL�z������md8� ��g���u6�MDF�0౏?�O��	G��.�"�����c�,:�#�0f9�+���&�3�SF��s��>+�0��Q�Z�� �pO�l��o�_�~���2?|pTw�ݵ�#����*�d�_�}Im�>�t��0�?�k���eN�����9GAՑZ�p6�����4VBI|6I.��מ�e+�t^#ށ����M5�8��f�v\�h���![~������f��tAw�P��+/��9ۇ��ԢRך��E���ki�S0\��g[�ٳ�ޮi��b1Z�D*���f�;tS׼�epd`a��KC�#v�O��m�����l�s0��-^��F�ޙ��t����x~=UB瀲�qy��^�5W���+P�����/�4Ny�Y��)ʘ9 ����;R<��O�i2��({���τy,^�d�,���t�"܊Xoz����O���uk6�}MO�����A\��L���Yg���O%�)������6�-;���.���7�k=y�� ����>�9c\�����T+<M"i��9���� �y�\��c��	'�yHO��葛MXp���E���Jv��mT��4�J�2vݳ?�'z�?�(��s����]X���9��{u�^7���� ��o�}J~���t�+����������E���x�֔�}��D�)��+aj��?�e1zTx�o&D��͆�?���Gř-[w�ǯ���G�||ֱt~_��T�5%)c7+�0ޔ�!;P�`��(��ᶥk��]��b�\/ӧ@����ꉠ��Y#��`Ϙ��Aqr&h�K�:�Ntڷop�1t��J.V�Nj��fWhOu�pg�H���v�����ZR�PJ��yh��=�)�����j\{�	)�t�U�^�H�Րې	O�\��/����R�t�i�_o���3͝��� x ;��TH.<'�@�_pݘ�{o��߂�s,�g	���(n'�����'��Bv�@�Sx���R����ԫ!��u���c����gC�F@'����@oآ�2p]z�t�qx�~�P�t{�2cr��̅�0�Z�/j6]��fy��b������#W31����˸����G��ݯ/���eE����\��(L�(T���h�L��H��b<{�z��S�j�>���YX� T�jay�We�s9�o
J�ۇe|�hf�tG�DD� H^�\o��Պ�vYm��eO���3�ni��1
���m� �Y9�\����1_����p\c7D�O��ᕷO��@FKgƍx�#C�;��j���)��a���v,��~������m� �R%O����8	�+0N^e�/�X-�F߱f���;P�仏>���d-ɖj$N�Z��Ǚs�;X�Q�C�Ȃ,�ǩ��s�.��o�-��LI.|p�7B��l=ӳ}D� �9�L�1+^��[�)���u��X�r�=}��>'��؀z�AbG�1�Ђ@�t����͛sCCdS^���-�]�R�}��� /��~�{� Qn�M�`�u�$�ӭ��"H)�w�	�,a䂄}d��	��7L4n���9��a&.D��k{�)�P�7 ���.��(b��8�+����R8�%+��G��TҦ�^�C�ͽ�M\��=�Iw���6F���0E����C�n�6�Z"�E��R�]���)���~���`��F͈%W=PCq#؍��S��b����-p�q]1�Vt_���o�2�WI���њ�y����]?�:�����%G�E�+l}K7�B�(lҵ��\��A���%^n��cP�Ʈ?e;-��:���(�D�9j\fy�Q�v,�Ѝ,��o��U�|��jl}x�K�:��ŕ���'�\�ALB���LF��@��_�q�<��7v������0�!�J�'ކ��a�'I�c�K������j�57`���T�묧��I���ܕ !��"�+����^�̀b�:����$JC��n�P!�
N]B��F�
a{"r��tuZ%r�ab��7���n	���N�Yo.�TPu����m��m
vQ���^_B0Z�
����}S���Ѯ�����j�e5S��Ro��4�Z�)5��[3m*
��Ըi��=��A>����}L���l��������&�©__�a��c-{�)+1����9��g�w�s�{R��8�M.�W�ᔾ�~�4?E��j�Q�h��g�+̓G���nbM����	;�Vf�J#�eMQ�\�-���KXJ�Us������e]�x��Í�*_�\ֺ4�sF��Sy���_doM���X �nbm���j5�&)�n j�Yڜ��W�-Y;���m�Q�M*~����KF���~]R�c�.���\�R��B�l�%9����
X�p$�|�����4���V ͭ�����K��ޗ��\D�-y���*g��7���:#�*��Jb>������r���P��+,�s+f� UǷ����X��T=�&�����u�E�\���d3 ���4W���H��^�
���{|�`������+�AE��%x��L4MFeUۅ����F��z��{���>%�L@Y��'&��E�~�5Hu��l� 5������0@�V{����@�F$4j�]����Ι�a�b���8x�Vq����p)=�c,U�����I�AA'x� �gZu'a:���Ŝ�����9�FZNr�|����*�0x��w��b\��[���j�%*�e�0Z(y�X���������%/�$ l�����G������➡-G�*�|vW�F��ܮ��y�	C t�YbB���3��<.��� �B*J�2�S�Y�R��;S�H��Ƃrj��U�MGfa�:!g[���ȣ��
Ln�~~y�'�Vh��#�5a�k 0��.9B<3���g=�	�S@t�
�]P�E��������S�cd����%��d���־��KW�e��J�5����� =vYLL�n�g�9�{��W!#�t� �� �T���-�K���!�BX��k�/��4G�
P�8#�,��X���`gP3���6�Xs��~�F{_��v<���.�q��\�+l ��r��U��^f�y��5M�����ױ\Vڭ��p}�������mD�Hg�))��Y pH��i��23�����.b9`��&�j�4/�-=7H��@�ۚ>MDt0�>W�V�QL����O��icE���H݄��
�bm�|Gt�;�e�L��#����z
�/��̘#A�������Ʊ�d�K�~���e���X����#�#g)3�!�<���Ѡ��l���B�{N��dq0��iT��U����lv�k1^6��Kvb�}����B�OX/C'Ϯu����$p������A_��4�y���%7��I���Ƚ�k P�Dg�:��b�.�R;ǳ]���GG�����[A%�3�Zp�ץW�U���~�)�9�Y�0��J.���U���:��C4J6y�jC1�ȼ��F0cFE�C�"[�7�i�� Y,���ޖ~�	��GI�8�+�M������k|7Jd0�����)���6t�)@�m6af	�W��_!��/Bz��Z��b砤��/�(K�(�c��&$�:XnQoܱ�HLT���<��;�m�)�>k�Pd!��E������Fh����Yp#�G��}��ĵ#�j6� ��'�������,gL�/�՝�f�TB<n������D�Z�lx�}�|�:��Yh���8�H��p);�+P&����?l�����*b3�ڑ�-V�{ǻ跓 ��E�u(���7��Z�n� ��N����W���b����aX�O�Z���VLI��Y�,���j��&��~=��&�'<ײ0�;��a�S}���0r<����6m�O>^���Q!L�ˌ"�֌U��oz�U8��X"≺�jO�"4���0��h�lٺ�:2=�M����W3e�WV�����1& eu�CDkn �]��|
� �&ľŻ�����g"Y��"�g��
d��M��o2�S8��[�b�����-���}\���ML�$�Ɉ	nE �a��2(�d��9S��/B��6�������m�xB�l�?���>q�NA�Q��'�{|�<��.ӹ�fS���/ H�F
�[kQ�
�$��w_vm�lɛB�&"p��|�:N$[N�Z�h���x����5��t;������ޟ3W�`	�ݜ.���r�=����B#L�*��)H�έ�WK��Q�t���GU�ǩ�p}��v�Rb� M�P��[f�m���L����V��}#�IŐc`�'��ko�{�i��3d��R
���'��7���,k�vW���7��B]�C�"l���J��^l�*��cH��:6���6���"�1�1_�ʹ�.��bP;i�8���D�B�7W<A`�NM&�m������
�YnZ;�����Ȃ�7ޖ�3W\��p��B�E��T�Ov�Ӡ.⇒O�)2��<��F���OKb��,�su31U���un��RO�����S5`z��Շ�&n�e�ܤ>_�	�CW̲ω��f�q����-Wωt+�\��B���Jv����y�f�R��r_�pK���l�EF�CV׻ah��Yn���ĺ��؇Ip�q}h�f2���,�r˰��������	D8Zys���o~{�{]�@ �γPDGQşX��:�n����no��Ie����HVAx��������镐]��Ƚ���'��)��,6\r�N��R�x\ɺpǀ�����2}���-�Kcp�<�
�1��K�ϨD�!���I��CN����f<��[ǲ��|�)���g�|��s`8+�"��7���j�E��eE���2���E(�An�iÜ�l�ߜHQ��7�;T�Ie��b��^���%�_!�H�S~3��l�o4)3|-9��Oչs|�Y��ϙK��_��&{Ѡ���(������=���ɾ�[��ߖռ `:����}�F#��}��i���iB�i���Mh��hՋ���U7ss�ipM���V�aVi�OV³��}�df 6�k�	'G�$�Ƣ�;2�Tͨ�!Ұ�U�D���/ݱ1��K���9c�ץ	��me�4�"���X� �_6�e��J�3�"(��y-��ﷱe�h�0�����A.���+�A�N�U�D����}=��:̍��z�l��-X�A���-)8O����«?��H%ߵxQg႐������?�@��0��%F����}�ߐ���O�q'{�M�WN��$*V'i���E��U��Bx�Uᅔ��Z|���S0 ���8�I�����.�s��"
���
��InRm�Z����������;}��Nb�tIF�MVQ}��(g吏��U���@A6-�6M���Z^�u��K|�,��Tjĉj~���ٰ�U]�E�gJ���vw�6N;�|�G1ah]�G��x�χ�`�rKE�Ŏj����x鬍����½^��!:�"Λ�B@��d�ނ^$��#|.��y�;4�iz�RԎ�	��f��k�(8�7�n��<G3�!+�H~�h���J=��UO��)�J�H��5���?j�W'�y��϶Ke��Ą�Y�sK�ە���7���
�a`2랝(�t� �/Q�z���|a6�7ϣGWL��:A/��]� �i��:>A5U�Q��Qn�eN�u)��eR8(H��Ӑ�'�9Xd��]]���:��̴��(;~\4��s���Z?���Ϟ��
��<��P��kt�m߇�J��)��9��+�w��jvhEX�Txv��P�äFr4�yER��Ɠ�9)?�S�y�{lЅGI�W� ��S陎�^��DY�?;��ٶ ˲
�������Z�k����H7dS�T8Zpy��.� ��'&���%3�ED!Ona���E�r`cuۥ	r��㚭d�Օ�^�&���n�'ԇā�x�ǿ�kg�����p��TI���6�������,�j���B:�p� 9M��)�}�� �5���R��K����P*� ?s�]	��(�%X��A�T��ˣ/��2�����ԩH�W��\{���·��`"fn�2�
p�}�7���U?�TZx#����G���9ˡeKY�v���E��L�~��3O��W��F�Y�1ɎB�;�`�! *����/���k.�jCM�G� �}*x2��h7����5�ˬ=�:�8D�Ttˇ�$� kbj�	��Zl=���}z���FJyߧ��ޱN��=������wFM���<��!�9�oj��_?��1cӚW ꐘ�p��8���f~��\�G���u��G�X����)D����R2�Ȅx�'Dٚ���f����۪��MdK'k�e�7�>�Xƻ��~�H��qs.�����{]ެ<v.*1(H}Zv<�1����f#L_R��ǿ��''BN�n�1�n�a���:M��Z�S;i�2'�!W���,��@��G�^S��|R3jy�w�v'IE�K�W.)�~>�ߓ����ǎQ��ep"2B!�S:w��E����������ڟY\"��-1$F��/�+ŮH���H3�D87�j�w����ISY���9t���Ҫ�)N6�+2�k<H�Q�k}|N��f��vh�+_��#2�FcnCES�EY��:�ݢxvaL_7�����3�X}}>��/��3?�=W�Y�Lv37f0s��k���^bj�׸x.[t�ꠖ�����~���/ǣ��o]q.Vz��nm�B�d���<�4자�>D+���S������0N5�_�A̬)�Gh�ԃ؈�f�6sh��w�~�ֿ��_�?�D5^�����:0�iw�I�'��=�Z�L���<]G!�hsSVkB�{r�	QF��4ٚY ܋����4��X�Kޡ�»X �R�˚G(� �0O�w�2B��h=�&]"�[����6�f��?�9G�oV>�\��+�;�K{r��s��:�f��?�6�^���Բ�l����N�%�r��1�D��3I���e�T�0�16F��B��(c+��^��ѱ�6NAH��LU@���H* �̾i������L��WM�k�5�L��}�
�sW�|,������L����>��B����Ibb�7�.�U��|]/��QTה^'�}�#�	M]�цx0�y�0d|�m�-�b��t�B�&w��TU͇j��?�|ңC����7f�$l��A��>�M,�*���� �cm�����KQS�ԙ�┨z
y!�߱R�I7A������D)�n��\������".�Gj
���P��1�� ��aYh�-�XE�Ը�N��W�퉻�X�8��?�Ό��4+;a�0�Q@�rP�ն�/l�0�fV	�����E��62_ЎKl�O��$>.סv�)�7�XKl�@Ģ��ab.Os�MÐ{��AR^�������#X�/�6��BC�h�����/� �H���sص
����xF���B���%�8h.��>d ���{�F50N\�Ͷ�y��J���ۈx������J��Z���K��X�`/��H29���Kv�P��#�nr��lw|�n�lj�
��Be~B?P
����@�&ckT��%��<ao��Ӆn����|+�B��h�ZK����E wc��j�NinR�����ֻӰ;�c�a��2�z��X2bSCj��	�kL�y�BXz@ذy��0�ƴ��yr=io��Ew[evt�}�9ʸ$t���n	�T����8-jRkz�X�`p�HX���t����#����o��r����l��y�=8W
���:>!f�J �l�C�Zy�D��)�z˘�z���i�X�����P3���b��숡+ҧ����Uka�)^���$#�H�$�[Aœ�*8۴�i&(�V�g��q����'tk���}Y�v��`|}T3�Q�H1@���$�L c��j#��*R���}8�=1=�7��!��j�/�
5�����h�-�_�m��!7O�4q� �0	��ҽ��Rӭ��VKE�Z���F�B�����ϯ#��n%fC
���|D�{ۨ�Ҙ�]��B/�M���<��3'�㰑��04��D�Z�2���ً���_�n�}�V6�&(�J��������M���cU�ysN�~���o�*���S*��N��7�\��b&� 0Z2�V͢�A�il�F>^���ګ&D��W������պ_h���.�\H�8�����mt�YS�c�Ԇɍ�,�38���'̕�G��g�����^c���`ٙP������os6g-��H����0J��N�}��jɒS�vFF��	 1�k�n��/Y���}�H��� h��X�w�uezǰ5p��զ��]z��&y@4�'�@�E?:~(�J�{x��c��h=�!є���Fp��Z9�kt���V��Jl���Ⰺ��y���&��Rs���eG!�e�/��rX5�h�Ue�i�%%_��o��ȣ��Bnqj�1n��%��>>���ƿYd
V����k��T- �gT#�'f��/�Q�(k!�cg�2�_<��ưS�%oA�]�`�Ma� P�$�챀~������XNo�2���Ǐ�����$N;��~1�24 m�5��:�QZ�jU�M���3n�Y�R���, @�da6���)�x����+�� �O�)O����T�w���?��1v�iIr�q�[fϷ�_ -��y���.h�'��e�m��w6R��at�̜�W���ï�
�m1�j1 ����CR��vR֚<;��eW���Ñ���@�u_�V��~�f~GbZ�s��U����`��>Ȳz!�@W8�e��2>%S��^B$K�L~��-����d�Zr�,�?~�^�t�a? p��d��v��thٵsYu]�2�g,*}��0��?b�� !����]�P�yy��A�z|�ٳ6�ڀ�z�P�n�� �$(�"���k����(p�08��PgO
=>ULd�S�Ab�h�Èӈ ��ƁM{���A6����7�N#l�M
�&���챊�.�TOvY�.e�Og��4@+�ǫFT�A"L��lcj�&A�g����q��|?̈��X0������qƢ�ڷ��LES�߲��&u6��tB����+ƥ�VO�!qy��c)�XlT���r@�z�5)%������6(-����5�8A�����H%�j��0ě�}(
 n�eܵ�̋7�R0��Ǘg���夆���;�-s���G
��Ʉ.��v�a3�mcPx��$Lb��}W�S�T���G���aDE��%���_��h0ς}������H�fJ�=��0-� )�\�p&��P����Fz{o�4LpW޲_�=�q��8�[y��|��^�2��������NQ|� �c��Ɩ6,�\O�y�>r�&׶��$ljl?o�?}Jo f��^0Z�F�0x��vs��.P�ǁ��� �n{��ŏewjxp��^���as_Rd,h�����f��'�|���h��]�Ԇ��	�4\r�� )'f�A�@j�^'�jt$�5F�>�jԢ�}`��P�z0p�$$���C�S��N�-�0G���g����/�� Z3����A�L3��烠�Y <#z	�5��8f<+slB!

��?<��|���OK����)���w������d��ʄ��Җ}��3S��roH˄[���t��Ƴ�;JE��V�:v�C��a�畎�����N� ���&Hr؄��+����>b�T�i�r�,��x�
sB�5\�%��w\����<e��C��"k�#S��%j��a���HB�uf���YF�ۢN�?�24���҃�,Os����L��S ���gB%����?���j_T�^�ť_�����	�i<�` V�p|�Ng�ca����QI[^�W�$�����0-t�@�e�W�����[����P}��0�tdC��\��T(m?ۿ��$�h}�}�]�\t�L��O)cup�"�N���gԛ�%�WâO�nҤS���~pk퉜�_�x���.\(�/��9-�7a̩7q�Յ�!�_%Be��=Wn�K��5A�g���s�3.~>N��)������C�]2�laP��)�zn����9h6�"����] H�n����eI���;]ӎ��{�� �� H�q]V
�|�A�~�����ꯁ7̈J=��RA<]uN�w�������	4ShY����.bIt����s����9���̃�Mn���Ueo�����#�D�� ܢ/�p����vM>�ʑެ���{9V��T�܅h��u]3��g�o�1n�DO�S��Sv��tH	�d-�5�8�љW��<�L������/;����$���Aw��$�K����z�jy��/y�
α��Żv�༢��G�l��AIk�}Ab��O>� �0jY���,|��.�,bw��b%�}8�����>k}�T࿿iE|�mSތ�U�0�i�]��[���g���?���G���Q�u$�~����qAl�~߼*����ڼ�A^ɝ꽞�UO��Zs����ѽ�^�~O��*���VLMZ\$E!s�Δpo@�[�_vd3?*�{�X��d��`(]�hA�0$�@�w�99y��O�T�h�8�n琦!:�ƐT��=�sO3����'� a`�QA����l����������
���#��|���9�*Ƅ�����/h-H�7N��A�u�_�J`E�(R� ���3>p2�^�\��� �a���?��
eM��cbTóT`޲�x��Y�(��
��k.!���Jng_��2 P
��*S#qf�B,�x둵�q�)�m�҅�)?;S���z^�O^�~$#�=W2��7C�,�G��pB��{��!�Ǔ�ѣ�z�QW`¨��*P��u���{�;����q����c-Q�S��!����I��ԑ�e衷��~�t2�H������9�uZ�~��;����ۓ�z�Ϳ4ڡ)̆&xG�/�Z7���T�:��s�K�z{�&ʸ��l��h"�)m7�s>��@�B�4z�P�3�'���Tv���"o`]E����5��g�m���v����K���������$#ߺ"�fq�J���ъEϵ0�p�xц�����c޼�,�oRt	q��K��^�援�'T����xs���v^��	f
O���4���Z��DjE���/���Ⱥ��6mS>��irf~v�pͿ�F?$�*��/]�g��C���H׷��ɖ�"����[<PI�L_���8�{�b(�h�C�`�f�����g�s�ϓ���	�]R'�r}a�p�R���x`7l/�y�h�.�~h��r���/��V�;�c�^�юfG|N�~(q�	�~�Vȋ�"f��M��^��t�"�����x��2���]Ji�1zۥT^?05y��w����{}�/��M-��~Y����Kڽ��A�;��V�&\u��a4+�sQ�.�ؚGW�=�s�#i2q�@]�9� �C{Z�] gU�S��g��[(��?W.�!Y:_go}d��8�C0J?��
���s2z�46���j?0
������Ѿ�G�όx%�A�G���g0�d,+�/ce~�a�@���UFSXu�I��D�,�;�Eb�	�๓�r�ڨ�g�J�I*�6�r���t¿�>�'q1�8�&H��:����~W.EF��|�ҭrL�(,�R��w�Im&,Ӌ݁���Gx �s����}G�ö�C-�@$iB�����)^Q���/��ö�c����+�"pE�I^9�_������gm+��0 �8��y"Gf�����0�ڳ��5"�x�
�w��D5J�LdtFT�7
?�%�2���K�_���&~��2$��w >Ü�u3Ed�^C����jʪr ���""�/��Ǻ����W$׆�bt�^S���6�a/M3�W�z�>`�+�t��sl�^�����6
'�N�ۚ�>T�-*����ː�F����n۔%�9	Qx�%y2�H �A��j��q_�g�P���D�T#�����Z��?��d8oC��<_�v�̀�y[o<�ٜ|�%mad@�-
̿7�����?R���__FP0�IеR٩��xI����&Ƴ��4�䐛Z�H�?�F�zý�0+*��U��M����5[�A����i(D���n���^+�, ��\��s��Q��^OYD�o�m~�z�\��<dK����F� )���F>�\d�e1R�OsO�b2T���<J�+��njT��K���=	Q�����jfaxˮp�@����/�N{nA��G��Xu& N��=�:@r@��e�vO��hȁ
-��
�z�����Ǳ&���3�T������'��7@+��I?���1�2�g|��U��~�=�_q#�a�u��\�{-F h�=�X,�섨U�{AR<������0���@�n Ջշ�b������V�JZfi��yu�evp �ڵl�)�h,P_��CQ*�uɭO�C2���R�hޫu�L�1=9��nd��<�2b�
�,~���P�=<���u 6:�T�(��Kp�MU�ļ�"]
��-vu��o��]m|�������#��a��h���	>}����2h)��Fx�M�A��t a��{�^
�l���Zy#���̂(ai:t$���ߢ������#'x�4�00OyA�Є]����\sI�J___\U)���5����a|l��І�������gO��3��z
^�8����%�S �[ɺzp�=�;��@���Cc�����ٮ�ES�����`�<k㍖�<��n��|�Ȼu������F��3����:\��[�|����
������v=lu�,4����e
?.��`$1�V�Ke0�9�E�{������]�pȞ��rt�k���"������+ ���$����p�����c�8~�;�L!FA��{����@�����p�4�)ڛ���EO(��@*�T�w��HN�v_��n�6���-��N(9�]|��I�{3�Z/��%'�TQ����ՙ��4���O����Mޙ�uBIꈌ�����2�Oo�Р�7S�v׹�;��`�v���|n �3���߷��)����辒��o���V0�K�ʧ��Ѣ0^ �իC�:T��lpNt���I;�%�p�=���}���_�z� ���})��d5]��l��'�*��2�nݫ�����M[l$y��D� x7>1!���tm�eL�rrs�b���~l���o���z�y�+S�{X��%a�K�F5dJ�y��&�\���K���V��=����ݦ��9h�:��
��)Ԁ퍶:��[������a�g�!�j4��`3/�u�U��|wp
���0���8�#�vAr��ŨS�f������^;����F�<�X����K�G�Or�n@�$���_+TR�rA��/Y)��j�!rJ'<]�N 'skJ��|�BV�_��BMێ��>�˼%}t�ẑ�O��8P������Dw�VUԚU���O���X.�|�Q*�����2�?g�jyZ�-��|�E�Z4}�6 ��`BK�����an��9�w<F�*%�&�N)�s@�;����1Ɖ��F�ێP=d����ț$�U��� Z�Ij�;��L��͖�u罩���,'ۻ�<�]�����C�~H��M5=%�8S���8a!��h1�D\��&z "���@/���BO��E��g�܊]6����<�yTFʭ(^�iׄ��FX*d�z�D�M��2/�)�e�BT�JR=11�r�ȗ�5���}~sA%_Wʈ:�	���@D��2#�^v7�y��d�h��O��rR:�m�����f���r�
�M^]�iX��
í�{Z�S6�go"%���^eh+y�Y:S,���[�����N�x=��e�lN��m<���-�Y͡h��~�C��5(4B��z7���#�b�*�v���ӎ�-�፮Z�U�d?0nh,���t���[�Ea,���z��iWU��w-;-3��>O�Ȟ{��塉�2d�+��O6��m���6rT`z�,��2ڳ,��c��&�c�PN�?=��L�p�\˩� ���aC�M>�T%52�b�N�Z,E�*2(#�r�n$hu���k�Er<���ώ�vxd!��R3�>�}ơ���w�ωYqr��섄M��{͡�M�����i[�4�9���a�Y���3�G�i��K�3�e�#}��}��-!祢�r����r�"�YL�?{��[�kT���#�d����L�l(W�40.{��W��a�9���|��3M�<�n��4��xܯnxJd-7��xdX/�4�c�� I��md����F@�*��Ux��a�)$�<&Cb��l<A_ٻ�.�d��D���Y ��R��}��d�;�DˏJ��Ԋ~n���*��wy�к)�4`���P�s�*	���*�	�b���?!�'d��f�3�u�X���!�>?5�1H�4��n�5a�ʦw��sL*X�w���L���v�	,�WULm���֝�=y_ű=v"��GB:у�կ=�+�<������o�#_ۚ��ߜ���n��z�����;��h�� ���DP�կq�)aA��W�Ȱ@Uu���
#��T�6� �/�FB-���қgd�}�lD���n�V� ������$Z\� 8��./+@�s�e\�7晄QFV&H$c)"�M�I��Ω{<�9-X+�o
=�o�������'�������hRş}�"��=��-���BN�X�=^i�h�)�&Iה��0e>!�� X�X^�3�Q?���� 5�Q#G<<�W�v.�x
�,�����'�vH�:9��Z9���;&t1*'[��"H��p�`�\�Ǿ��N�Y��D<l?V�{9�e(��p�5~�۾�*�\��Q�&����V�K�=��(
�	)]����Iv��@�'�^'	E��Ȃ���z�[.5��`G��%p<�d'��R,,ԗ�F6��ܚK�n�N]�� �V�XPt�����y��X��T���StD���6�4L����'lR��<�H,���8�0=�?Q���=?2V���v�u��)�ѷi�L� ����B�ʝ>��g�X)���h��:	�'��X��c;��1l�2^l7��b>�6#��a.X���گ���Z{#�^�|61��#��O�Q2ӥsHI~�M/k_�P��dBra���&�3b<�"RƤ�`nU*�����!�#�d!�=k�Ψ��MH\k���־�o�k�)we���&��3*�P��A7%��D�3��6��G��yL��D�&�'�x�s0�}`�vd���U�W����yh��kI��J_�E��v �oL҆�����o����~���,��2��t��k6���h)��9󥹸���?�q���e�@�Hu@Y9n���3+���_��5�����
N,��c�q,�`�5sd�Q�L�L���m�Re6�~:��죉�NA���	Z�j�y%��r�z�j �dN"�G�~��b|l}QA4Px@��:y?�V��ڷ��Q�g ���o�SQ�f
4� ��|o����ebB�Ԗ�,�àc���1��>Ī�V�2?"Z�'8�3��X���zU��(:���w{L���������Ec�b���%�8�7]j�Nۄ��+%�@�]���!S�ܯ�4)9y�����Y�=���5s~������{��4�����{ڝ�	z�L�mWK�y��iu"
B�lA�x��!h�`��o�˄�6�+�L�D{CNMy{׊�$y"+ l�sl��y��C�y��7��E�A`+.�y���Y?ɗ_!
�%\�s_��u��RSk�3{��w
R�x)NH�ȋ�*�������@��A������/���i��ٱ_�K���I�m�b<�k�Dpе�Y7��UG�����Qf�k��:�QVtco ��\���굅0g%���1���������e�Ezٮp(��#��9�'��EW�I�}�v��&������W���iI���gy��F4SW7`���a�X����ybDzR@�K�������6e�G����E����oUM9S��K���l����\� 1����l�ex�=��@i�$,'��_J��vK�/���hr�nf��}>\�f5Z\k�*ے���Ja��Pf���q|�[jd'$ �;:�F��6�)\y����F�*r��:&�zm��)����`�V4h�����w��,� V%��tS��u�oO��[��~M�C�	�+�r��NfQ�:'*�� �n,��^���m�������f�^�Fm��Ԟ��Ǌ�ƫ�)u2����Ww7�`�G��	p�5�g�{1�}%�	\����aښߩ@�l��6�D�)�m�&������K��������S ע�.���d��s�м��oYhb/�}U]a���k "q��z��6�Y���ܰ�:D���ׯZ#���у^fa̔�|���Y�e2t���t��D�5���N;7�V��,�\՞&�}���F�O��oC�zdf?�0 ��|y+½�>���*P�ha�s�~��yM�D�JtiY�|_+P�]�KH6��@������N�(u���|G����~���@�
���0�(lB`<=|Gj=v\Ѥ��Ü���h2�$���N}&�	i���˲%�f��ߛ�ӕ#|�<݀�z��Xɏ��ǐ������¡�l�A����f�\$�A�R�'$5�gQ�=���Xd�\�[�A9 #�(���c��5ʩ���y��"דh��������\��U�GkK��._%y�u:i]��Cw
t}!�ip���ׁ]3�m�����P� H�>*8�>q��!O��6�_�S�jd�+F�����ϰCM�	2��ʁ�z�}��;��r��-����ݑ�`�L����k'�N�U6��
5������*m��	��յ����ta�v�d��|���M���ۏL�k�s�xu�����э�ǐγ<YAV���6"o�5���8�hT�yQ<�u�>���:��U�����]f��r)�y�T>�B�9pR���6J�rM�:�M�� �^�<�]��g��82x��m��>^��l���+ʁ8��(p���P�}ٓ˭��0k��$��{� Q�v�[���d)�^�(�����"��V.�L�o�BO
�F�h�X�.wQ����0#�/��rM���o�o�n�I��Vn!�m~������WU�Y#0��6k��$�L���qb�������wWĐ�W�ަh���)�������j��^D,le�I�{�����G̢���&2Vcˏ����a�[�.t6��fo0�\�@d1��P�Õ�2��J��0tw.�z���OxM���ޤ�6�_�CrKpl̷e93'����{E����G8��M�5q7#��ɭ�{b��X�Ňc5���*~V�~��z�7�߳]����ZYh�#U���WKQ�l�HW����l��E@��/��~c�K�y# AR8���W�'���[
;"�k�ktn�x ����RK6�����=�;8����I�Tl7��n�W�	y>k�,�,=壗�;r��3�+�r����`��cʪ�
ߴ��S P2��9EX�X���瘲��w۽6?�追td͊zc�h;�E�Z��}z��|�����vUZ@d`C@b�8@l<%��i18�����_��KK���cq���2���#�}�g�cH�6��ۧވ���ȇ��>Ҹ��F}_+/P�9����;�z�ȕ4�k�q( 3�������{6�`5�<�S��Oz9yDp�����x�Zz�<ccЍ��-|H�r�#�6����yx���2�H�}���dgk��IL��֯�_��}�)q�x�� 8j��9����e��;��ce��amc"Ǜ2+��ݸ)e��3����ch s��w	�������Jq�O=�Ơ���Ӳ.�9];&E�Pt͉S*Bn�J�qA4��eN�x���\����@��L�ӡ��V�ȡ����NHa`6�j_�kz�1�p�6U�6K���CXUG���iب�Q����Hkbo�'.��C���D�:�#��+rCR�G�#Ō� o�[�x���_`�X�+���۱*�Ҳm�sں�����]$A���q!;%��B�^f�TV�>Y3�`K��%%�� &^?�i�g5�l�Z7����ꍠ��n	k{b'L�H��;PW�HJ	k��[ `�h�����e2��~��2��mوX�-���1D�_�aa���x��1�W�<M��5� D��׸lOkv¨F��
��O��"�Kr�$�ág
dAy63��V�k澐
|�+˩��k�5���Վ9'�ٯ,�P�Y�{�wPp�$e�S���t�]�j������`K(��f�Ƹ\�H��;�VSF�]E'0�:��K7�X�C�<U6�����QI�p��;���+@�EJ����Y�J��} G�Xh�c�(hp�N��,U�hJ�L��yتG�`�C�;���ǒ��1Kƅ����t�y����u�G��sPW�X�wu}Dᳯ��!M�d鎼��&��8����#D��7�7�K�'[ .�Ѽ��@1�;�'l����L1IDZ�zv%�������U���+Vm4��?0�y����Fc�ѹ�e�0��4o���͐��S^��]t,���I4U��Pi���F���JT�͗��w�����;6��Vkeb��E��(p�E���5��XS�6�F0��QP״�t�/�`�p΅����@���@1
�X���vن�R&,�ͼ+傾b����*��/K&�ß�N�LdǱ�>5+9u&"��f_�5!��>�'6��Y�3g���T������K�}�Xn���w�����<�j����c+��S2�ڊ����M���a�鵜��,�ȉ����;���I�b���t�#6$�]� x3:hD!�W�P�:��$��m���lKϘo����`��(I��rܳ�s#"%tR��8D 6�&}4n���H�6�sS���o��0��dV:����n %{ߌ�Y�8Qۢ��dY��>�F���@�nz�`���oG�xR�u?Cͷ�D�� F{�����P�%�3L���+��h�q�ᡱj�p��ԓ�d���L<��wm͌�TY�$D:�UJ��
�ۼ�A�]sú�c��1��}�빚G��S���2q�`�n�u��Xd�����ٌ�C�X<���i���Hiw�&?�����6�h�ړP��>�;2^�$M`�,[�lY��;�qՑ��7��%��Dװr�$�����7;M4���d=p\���_2;�Nhe�iV�M45%ߥgdx�tP>�1/���}B��S��&��w����Un�ťg�q+Xϕ4z��ߵH�{�
�h��Z  ?7A�[@$o��D�䠓Mn�$��S\ץ'-pϮC3Dͅ���$�>zj@ED�0���k<�)Ԟ�Sa�\��ݐN�Ø)�	�q!��Tdv�jT�Z���b�J�#J~������.�MT�h�%�&~]t΍׳8��+>X���G['	͆F�XO�S���`'T�<'�}�!S�������K9���M���4�Dt���Z^yd}��l���=We���_IR�H��cB#�ꯟ�c��"9��@Fx7� g(�sE �;�w��Z<M5݅��o4vB�����K�����Fi��JG�2�~��j���j�e�(�W���/��f�M+�w �p� �>	{��9i�so؍g�j_��b�>����@���wz<�\%�"NַǼ���ǢV����_6�}�?.:)�����2#:�O��S$�@�Q�0�])�Q�G�Sǌ�bH�˵X!�v�jjHV�֢�J5I��MO̓�|���w,�q�2��gbX�Tלǩ��}^t7���f�Q�cI��%�H��t9�����O�@ �d�2�'�}���YC^i���:x�Q����Y�cDg��M���޼�$���\�H#Rj��1Fl#��	J�.�π�E{�:eX��|�~�)�Z�߬����@0���k!	��XnhS���3�)�v-zX��"�2�Ѝug�\�z������{M/� �C!q�����r�*��^�&;�頎qn��/Z&��w���;ʖ�n�ڑ�"Xj�}JZt��K�+�խub���A��LH�[[�� �5Ø�ni���{��〈!�NF;���{`æ�C5�'҉�X��w@�P"�O���bȭ!7씣��I��,�V�X�.���dP=�����ۨ�
��hu>c���qT�YY9-@��Kt�a3��QeՀ�wܹ�1���}`�jك5������h���s��4TvȮ��
��>2�ǧP9��G؃���BE/��-�}���Z{�r��G)�X�(�;NP=9/�tG�N8Όr�*rp0�n��<R�YX�'R̯SI�/ F<�*!{Ŗ��X�;W�X���]���cE���Z��I]�T�U��Z�G!6�r<Md�"�,������U>^=��꥽��p)����n�Q�\�'҄���ܵ�\�5��ۊ`�IX�o��Q��RON�l�>�b��ySi�B.VC�;�zѿdT���a۫�C@�K�'تo��ҹ=�EL^픐�i������׏Q`uG/PZB��iڍ��iʲ���<��5�}�`{��|�5�!��	�CR|�;��41��hsh�Lw��,�9�����F�)���]Z���52HM�G<P�"��$�;���r�?}�� �.�mO- �pV���2�	G�T���|��*���4��k�
���瀹�_�/��-pa���W��x��9�5�J'ds�����`	�����$^{�)!�1<�f�p�r��o���U��E^����ԅ'B�8�\˦=�spT(d0 �QwǾ0~�e!�w��'�"�_\Oo6�U᠗�]������I�� ��'��D���
Y/3���8�#/o�Y�^x������r:�[Μ�3�ȓ宱t^W�G�-��L�\TY箶n�<9�&��}��	|},�<���DmAM�U0�j��ƌ)4Bf��wu���6�X�f�KOI�J4'�us�����Ӝ5��N�N��� �xs^��d�C6Y��y3���l��JRS�kKs��3�#�6h [E&n�Yz
������S��O����R.k�p����� ��=[}����K�{Dv�d* �̕�q�3�7ϹP�mn`��p<����9���7]�Y�}9�,��FG��̫uʊV�0�f���Q������2_NT掋x~�y,4��r����,�&3_Vt^/Knk9��Z���z�����ᡎ��^p$P#��~��#Kv��>R�)�Mg�d\�w�FA�p��Pb��,� c��{k���L�`'�ō�I%�@�[�г��	?X?k-�Ӈr,曍���#i �V1�lw�"��v�zg����ߊ��UT�~`+�CH�{���P���sv����S�	K�F�k�~�}�<��;Ro��S?1�sm���NL��ѩ�ɏ@7�\�~��g���|V���]�-����-+��C�I8�W�`��0��;ڶzq�$�n��<|�;9G��7@�Quy���GsIC@�8���C���s��zG����.vkjJΟ��nò��`��:�f�V��o�+r[��^L ���Z-Ŧ����~L���TCzu�8C��'�3�K�Ώ��\���.8M�>[������1�p�J���t[�@����i}�AD�# ����1�H�g��	8���,U�uI�E��Q�Ϫ���kƚL��P���0�/��`�0�M����XX7��������-/RԌ�p��lM�U H\����V�v/U��a�x!~�U1�
)2Bϵ��&P��D&����5�c
!�\O6��F�t�� b�5P��.��c�#{B�d�,�i�[�__eaZ]����r\�^I�"�g��bL�Ic��Xk����߀��qC�<��>#0r`;F5ᗨ_˸�,CQ��ό�x��v�MO	 ˠ��a�ɚ��c��p��4��[!'�x�=�s��
����%��7�/[6�u��p�>���r�&��2n��{�ʮ�� ��]��)q�&�f'!o^kLg29�i���܆n�z�~v��@�I]���%
�b�c�~��z�2��3[�������J,'�"d���Kw��ò^��R��F	s��\�Y������~h{'���a_��5�v�F��9)�����f��)�
�U���Wm�v��E;�c�`0�C9O�S��YUrπE�!Q�,�n�[��#r�(3>���x�(����B�e2�y��ET�\���Z��̓lG�����Y �ؚ
#�W�iNӁͳ T	$�� �$���Yh^?�p:��;,����Ȕ�X�Y�7�ޅ�YR��Β2~�
�J1[�}7��K�4ҏ��u�?�
.[�t5��	�f�`q�ck�@�.�K��'�� ��$x���sA���Mo��1ɗ��9X�
%��j��^P�_���ͺ.�G]�'o��/F����|(/8<@��p�NVƖ�]��4"ʫ��F�E�i�ЫY�F�G�#9��'*�)|�=S���V&����m��]f/z�	�d��L�g����/v�l�p���)�
� �%����.�Q{.�G*�F�܈g-����텵dEk7Pqξ��&l�C}��|�4B�V,�c�:�P��by�٘L�C�ב�ڙ.�~C��r&Y���(�ɜ��o�Y�+�R�-�-G��qp��i^̐���6�и��q����MߡV����?|��-��GB�ffn�,J�R�6ߌyh|�esK���E�(�k���P��r��$�B �������OP_���Sw),����%�W'ɞ��:>�4������SU�EmK١wIB��i�v�{�J�]T��Q`
c����k2�#1��t�N�t��M�ߺC�q��o`�� �̯K��P�m4Bm���5.��"����L:9�a�{D�|��f?��)�k6�0߫}m��u�Ĭ�Y}���~���z!�&�ŹwM>�)ה��[-�g�����Eg���/�41�5_HѠ(�h�\��-7P���"���9�̃��s5��ކ�F���1��"������~�kʜ��J7�*θ��0�un���W1ƃ��d#�T���3&�m
W# �=�5~��"��@�V�-;��T��q��p�8�>�H\��F��a�S>�j�l'�4(�4_s��|}�d� ��0�A>ܭSM)��k�S�~���+��u��+�a��B`�v��X�s�Y[��X3dĥ�l������jx[Y|>�V�QkV#��4*��{�a�b��m��m�s�Ľ�Ը.U�\���y��C��r�W��=��d����D����Z��80��HJkxЎ��{�j%_Y���#��{� 8�m����5_��VG����c[3\������QgK��>5�֦�iܘre"��bѭ��ws��8���ع���PB�?�AA�X��z��uv�ntmg��	B���Ї�3�\��f���
��a�
�k"^�ڦ�6��A��j���B�62#h2�o��gboG���?Y������6�,�����L�a�긓���n�XS}E�
%��䎀�\Gt����d��	(��]����������,J:#���x��\;R��b	�0����0��٥��½m��um���0AB5��_�7�}<�C����Ca�s�d2;!�;&�#�@��#���f�=�v�%V�;Rݤo����Zڑ�v�����~�^������G�TDh�.���h��(��AN����g���wW�v/-�.��쾎�#�?��'��3"v �xk�	Ua�nإDbF2�tvө�`���~�)�h���&P�C`��Y�$�Ī�p���">�q Q��'������A�C' b�O�8�_�*���NB�{H�.p�^�k�9PǊ%��-��Sk
��p6�|і۟�
q~��㕧&
��Z6�6E٠_��Vv��>AP��\�l��-��!*8�j*��4kP)Ƌ�)AD�%��6���$��!��
:x2�x�N���\�w�9�1�,4	:��G�(���#�4�@�f����c������b.jʽ��[
 �tj*ҮL�h���`�����Q�&�'�<w��E�xxv"+����A7(���d�_;�1����難��#���?��|��A�]�4�p�}����~�$�}h�QJ�i�L�Ik؜e��K�t;����U� ofE���$/���� r��&�7Pf��U�V[ήRz�+-���=P����X#�,�H5$=�-��O�w<B��]�ΰ����	[����"Q�>�y����P0�x5|�2/�e+�8��U����'��䆌��A��bB�,��@�?�b*�/8qTM_�Y���m*��7����'����w�V��K?�os�G6��OA�H��~�7"~���[��"G�gS��W��Q��cF��׬��y�����0�F����wXf�ަ �=�{$�m�z���ʉ�1E���}̷���vU�#��<������S�w����<9��]	G�2\���V_pa>1�$@�A���E����A���[��)|.�`ɫ�S.�^�d�Ό*�
t+Jà�e�,����َn��'\��ptZ	���6X:�+USSn��ƫzX{��=��n��.8q KO�3UP�^&��w5g�/q�n�@�U׊��H�]Y��k�����FGs�x�����֟)q:����*_���gw&�2�>�G��X�y#���x���p`c�fG��L�7��B	Q|=�~UcSn�Z�������>�r^�%gmZ���W�{H��9,�z�䶧Z����5�g�X0����*�~��
��eЏ�An��0H�I8x��G6|�9	�41vp�Y�������6-V�C$��:����FC(�va2�r���H	A�u1��`��v\J��c`�,�2|�=#�<� ����V`S����V�Z�p4�fS�=I����6?bŒ������n�U�-�?e�hn��R�H�� ݒd6��}��_�"�dY(��>�!��/)�R��>1r��E�E6�c%��ڒ6�Q��:�"��-I��>���s]����P�|A�警� <��.�,��Ԭ���f�� ��!5�鵵�T;�ڧ~���*~�!i�.VSw���r��?�"Z{¾՝@�W",5'��=jSv��Q�*�4n�I��N���J�
����0���(��/�4�tW؀�ڮ�b���G�;'���x�q2pG�c��Tr.�4�\�m�Е�>��'���0��%�^{;i�Ѹ��/y5�ɫ�O�v{�g���L?�8qe���/j���v":���#^�AI��oVߝ���]����B�;hH���_Sa,���P�Q��T����"��Uқ���6��"6�O8���G\GSIM.�FwW��J�Z0W��:���;��v�������Ά��.H��~�����W0�oٍIo�+jLW�θ��Y$�S�`��/��I�C����)�R$W���."azX�y��J�bg���o������5�<�ʼ}�e���˃E������]�D��F����3�װhH�Q�3��_��
���VL�J�x�xp�(��P�+��`;��ћ�Sm������Ȅ��Ti2`�P���А'��mw=F9��@�e����2��hB�L�"%��6��链pm���X\�J��Ϧ�_ӧ �>��?��u �R(smd�Q��}m6��j�kr������9̈�O�E���t�h�b����C��;��@L����R��������O����V?�u��	��P؂�	��Nz���
�:�b���<�-}�жAS�׹����2���{P��*���_�M�Q`���a�������TO�@��p��:>pŉ_�٬�R6�p��S{<�I�E��{:Tk'�w�h��S����#+�~_\0��c��V'Tv,[N����{��� ͋��:`��⍛�����+��z!��!tDOG���7&:5h5��O�1K?K�����ই��[�%�
��*�$h��Š9���lw+��F�R:���Fq[��l&��W<�p��=�\¥�/��7����i�����3��>ç�K8��y������A���{݋%���O���"E� ���*��:J߂�^��� ��U8:t�^�`ryv�хCԃ���ղ�w��rP�����Ljmb���ǈ�x5nn��DR�7-�%�X���m(L���i����"Ʈ���������@�j�`+h��?�W��,<�$iq0��\���>d��Ⱥ��2�����{_v�f
����_�n�����,��o��r�P��4�����u���:Y���y=��7L�o������~�H����<N�2�ːߗW��U�����oL�X�}s�GΎ��8fGMm��jy�q����x����2��NN7Ӂ�����q:f�ȣ:���B�C?-�[�Z�n?˽k�:��zGyIAY����^�����b����X�y��[U>R��^�Hw����(�|b޴��"��N)I�hY�K� �3i]��b����A<\li��5�%���q)d�@]���m��e�n.A�%�<�"��h[���p�u)�-JK�{�
�'}a�[����I[=ݕJ^��+��n?��а�]��?&?�m�(�oK̗�[k%���U�4g��/y�
Q8,�9ߺy5���@Þ�nV9�Y��6���,��G�ڙ��[��k+[��Z1�,�����i	���+�3L��U��N������N'Z8��v�D���)0�M}���-�w�0U}�P���R�i��o��'�X�>ױ�Ñ@�#&|Cte�o=s�����d<y����;��XB�Y	��{��g��>�X�q5H�qyQ�(�H*R�rn�Ѧ��r��D!S`+Iuӕ��6�&�v�Ml�W=�2x1S�i{#GF����Y�����C�	f]s߆��&ܔ2W���������#^P@�3C��eR'��Ooq�+���4��Ƙ�����ѧ$b���b;��]�a3�9\���UD5
�HR�I�^�~�~��-޹/x�	qh��O�o1�8u^���4�پ5����.X#�qwψ5���	�<pJK�5�O��x�;�7����V�p��I�Z
��o���X�8�7B0$iSK�ng�9�iQ�6{�Q�1��:P�����?��K��/������T�S�ﺘ�*����* ��t�w��U�d�CB!3��� 2?�M�&�\k#1Ѵ��8�N�a5Ԡͱ�(�cwu�t�8��3ݵ����θ[c�g4I��򿀄Ttk��R�0Y�߰�?�r�s�$��c쓒��i4�@��g��Ƃ�o�+S��4��~D�a)��N1��V��F�^sI�LE�Z2��x�&�m� U�3�`M��H�C�O��O�@L�]�#"*��Bb�U�4q��/}��z����{V����5����FC���N!�O�-x��.H7�P�㸯�ǜ��N���#x�A�P� ^�����{��[B_\���&�-�K�C��o��m0o��Q�O���	M�}./	%���<&��E��b2��,�N+���?�s�w��-�5׽�Ά�i��yN 4.��b?eƦ��J�='�*�����p0sN��B��oul��R��� �d�=��^��'�{�߫�]�~�,�VsЅ(kDnIRx�;��}e � U5�F�![�xEe�)*�
�j,u����x�@���-\"=Q�"{�źa"�˒�������eV�
K���N�4�}W�7g�������!a�����@�J�a��@z�����1�|�������T���!r��!��`;,F��4įO�9Av(�$��DPyg����#�ц�� ��5�{�Y��Kf�?x.��*�d)����&1��]9ڰ����v�r=
�<!8�kn�<|��K�>�M~����$lO���cer�6`f^�d}}2���rj��5��({t>�ǰ�t��. �c�1k��S�J�"��*J+��NN�7&}��
Cb��,��{��;���c��~�6ˠ�k\����
	z<!�B���&֨s�����컒�{a�����1淪[>���W����Y&�^zL�s�8b� �}'3�^�0�p,����DH�~�7�¤c�>�G�p����a�-k!�6ۘ�?T7��Z�PI�H��&t�m'2p%`�BPu�"��6���3�j���.b�#hKQ�,��{�D9�Ѕ� ���d�V�5��L�1���Ռ�+wL�}�ĺ�A=GE#Wyc��0��H��I1VD#bJ~Q��M~�;���|%�� �3����Tk����c�����y�s3a�fR1�d*e���$,.K
�K���ۥ��wQ�%"���PO*^�"�i�nW�|�Ee��Sv�o=uI:�1m]����Z3q�0gb���
�m���2X��џ�7���X綔@~\z@v|1]�QNi�N|��a�X�u���"�3�M��.{�sDB����#�5(A��x�xZЋ���.t��3����_V-|��5���G�n\i�O�6�<=�M��ֿt4��;�/�X�	Lso0�Ê�Xo��)���DS�&K�Λ�?�m`�K�>[����Y�Ѣ*9x����*�},��s�T>.�HN�r����z���O�QpA��4ĲYg����`W��f5Cā��]
Ƚb�W����G�X�J�������W�,?>8�㩤С��k����K�Y]�C�N�K�#C:e�K&䬐Ͼ���M��f����,avX}C%�|�a��)#8l}��e�b�p�Otꛒ��Vo<z\����m�� ���םb�u$�b��J$�)ͪ'�� m�8p�*L�S��t�\8��q�|�kZL�[p��A�.�C?�`-D����Fk�=V](S� P�����F���ۭ򩭠�6�A��#��8�!G��f"�+vyG�/��<��[���_�py=Te<�x����(wl���	���t�$���������V2������l������W���+;��tt�S7/Ȁk{�|jŜ��"�&s�Z@p����e�>|K���KČX�C�G/�n,�˹EBt˹(���bg����I.����$�� !���� ��N���[k|�̺X
 'V̓
Or������������c��/�5���6r�%��Ɓ������&�o��p�=["�"�Wr��iv���8�ʁ ���4�p�%)�u��f� �����r��f�G8@ [����;*��ߧ���i������g9���*c�*3�,��5j��g��K)g9Ȅ{"���-?�t�)���)4�\��br���qCS�a<q�qXd�$��9d$�8�)�	&rا���u�a!A�3��ف bX�\4I&р�>��H�&\	Ɂ4E���Ә}p38�7�m�2o6�{�HS�$��V���^�?��m�8���G^_�jl]	2�Nh�Ǳ����W=("�6k�*=� 05���7��K��$���n�G�'˜���TnT~J�{����'�OEi�������Nz��kh._3=�=#������_��1ݘR�=�5�d>�A.^��;a6�����5�i�C� �����_�%����`��@"�7�(�%o��<㠎SyE���얨,�(`~]����p�E���U��[z~��൹ \::��A�w'��q��1 dE��~j9'��1�F�-����݄�h�����q�Xg1�:�15��^�AW�u�Du`�ƙY�l�r��+��{x��A�l��P R�AЗ9��U�t�[Y���Zr�y��� �lЋ�����%���!�S�'���J�	]��@�Y]���,5Ʒl��6Ŝ��[�3�<�P�װ�=f����W���6���a�LF�-5hx%i����M]�؎FO2�I������A܀�pSQ��e���l�O�:�L�FM�A�����wii�����Y��'��x�ЊSJ����r�����bҖ#92�%J�<���:�+�O��|\d��7�Kc+�b���wUt�B�O�q�te��?�J�v�>�zd��@�����S}���rA��+�Ϫzg*�c�9#�9[��jY^�6��>�=�d��zh��\�r�Kf~I�N����h�r�9@:�mP��dφ����g��%: �d�`*O>TB7�[���,�(�U�ީ�_a;���:�Ϙ��"�)��[���;Okep���.(��t4������O���OD��˹:N�<�ʕB/ޫمI���v"C�"���X-H��q����T̟N�p�V�W���L��|p�U�n�	P�*f�qW��}2��sm�_ߒ�t��sC!�K�rLRa��K�6
䃲Z�:bs��Ζ���K�TW�a-T�}��\�T�;9�?�?Me�������v� �L��\K��b�
�Y+��'�~S�cb0J+�
2����Y��]���71��>�K
��J�\��
Bl]B�/>\Rq�흤f�`~�n�?��=� ���4BG�X��[ߒ�'��gމ-��>��	��t7C�!�0#�ӌ�[���+d �4�G���yT� �&��Ln�ƸX�v��9J5�m�9���1��2�h�6�9�R�P�g7|���L��T;��x�N���r{�/�
s��C&;�b)�g?�Q_c볳�Z:-�V4O��%�#��W�V
l#J�,)�t/��p�N^-�E���g���V)ɦYՃS���R/�v1�E4_qi|T|oE<��.KHW��f���t�,:���Zl=.��£.\�Y� ���F!crXZ�a�X�8�|8l�����a�4��T��G.���n��!�ě-@9�Yp)��@*�%|S�	m�$�`(!M����1�;�tO�>_�V�'nTX]�!�c�o���qT����?�"�w�@(֯~�i?�aWX$d/���?~_4>��gJ�F�1�����M��=5�]9׹��W�v�� ��F@;��"0W�jqx�+}ͩ�^�R��J9Pl�/�e�~��EWZ�Ɍz*I��^<Ea�����.����CЀ���
���7\OĶD!U�9��=/�3��`'���z�(\�9 �v�WР�4Y�ŕ�?S)I7*`;Q~ڢ�lzW}��}���;oZ͂����S�P���gI�\t!�O}DO?�zv�@(���^ѵv�Ut�'�/g���<�8N�!�oK��8�L/�`"hZ��+��jg�棝@
+IxG�!e{t��dCu�N��t�v A����&���X������*�ޘg�iыK=&�e�Z�6?�{t�$�E���N�����<v���c�`�ᕺx'���X���ARo�I���ۆ7͐jT[b+���P��\��u]������'\�=|h���wlt�& ��í�6��aP�{7��:7|�ǝ԰������\}y��E'+��F�
�^�4�����E�p�bS�j�ۋj�FT䊘Pt��~��u�U&����rA�{�6�A�!w�k�1�dR(i�n�~�U�<�N��W�u�d2�5�%}�_3�/���$f� 	�C�~�d�o
୊ӫ�q�!�� f����mG�+9Cy�H$\r-�^�H�aD�Io�2:xW��,R�d{�Y���-/q����Z���L3$�v�B|���ݒ�����5Qs�@|3�F������:Oo��m<n��#�G�
��u����;O`����(N8 ܯ苉�/l�2;";��4ٳݤ�8��qX�w�@c>�	W����Ii춫W�\L�~��q$%�3:}��_�֥�����b�?$|G�ߦ���?11M�s9A��`s��w��r)M���l�Ιߴ��=�=��7�him�Ä��a�z�6
2���s���w28"�π�\��= ��'n�����J�!��8�B�1{�R�h�*[�p�F���8���b�p,䔷�=w�B�:� I��4az���
9��77�m� ���C�ԡ���`<Ҋ4���G���z~(LO��NA��*P�uH��.3��dW;ڳ��2���f�����di3��Q]\�_��.���!<���ѹ88U�����y���yN��'}NDV>a}�jaZdr��|g����=�� ��[�?����1�B���5�&�����=�� X��yR��Ӳ���6�Qjl�t�I֭2��Z��+�YY��k-Z�~x��C��sk���V�<���qb�x!���Wyw���$ϗ3�9nT#�s@�>N֑������`A��~��ݩ��^�wEߜ*m2H��<�U�K
Rcռep�%�g �G ��N�['o���q;#a8<rL��E��Seu���eQKW���A`��m`ߞG�x`I,{^#���W<k�`�6��ʫxB$f
Ǫ����s�"�^��b��sE�$J�BkȠ���>^"�O[s\,�ԫi�F@\��E�~�K�������!GT��D���m	�4v�	(���c��I�!�V�VWH�>�q�����&�5������@�2C�01WS�T�i�n~�����C�-��/D~�B�n�o���᨜+��M��0`�
s��,	�`���k�%��x����n�4Ι��H_"ex�]-�A�L���Qe@^�|�����dDt����,�S���9���}bӟ;��47�`~�3v0��d�Y���a[?;){jt�ݥp��/�*�dЏH�T2����X�Lg��w�<�壟4�ꉖ^�����Q�C����}2�\��L2(�-�N�u�o��X-I�9��%�=b���b��M*cc�V�/	c��tm'5���B�4�uһ.�� ���4i�F�kr���U�I�F���H܇4�������h��PȱD��JEaӡ��6�W��bt�qK����T7���/���ǏZ!��	w7X#CE����*�^	�݅J��#�Vi&�J���ɹ㾟�LF�lg��\x�6͌@��Нj��g19���K��`������%��|����b�J*EQ,f���ъr*8�� h�������[���F๎PmƳ�����	���ȃ�6����)9{���Ec�t��S��s6�����k���O7T�L�ԏ��-��k���O�T�39�1]�N�EU��W�+�2͑�o^�]�fD=j�R"eaY����g[d�y�}�i4�8�R��[⩅�D��'�E�A|�;:YCN�(�S:�j��� F�2�y�SR�Or2����v�p�!´.����, ��Qv/5mp��Y�����O����{jՄ�7_X�-�S����N���g�ҏ�Ĥ
a�s�0��$���mB��4�?Cr)������2�Ś��sN�����Ok
?�١���ֵ�.���z_&�x|?A7!��>�*������&~�u�J�ܾH�����M�%C�T���uێ�N��.A���*�m���`5�9��ԛS!�.��#�'��*�/~�$���8�4�n�B=[4�K�c��x�׀5��6}q0���D���$�	������=���]�N�d�E�f�6+�A(�3�Ӏp�I#AXС��r_ЖP:J�	p�3E�"͝L��t�=�ë�%d�ێ����|�<u���T�75;�s{L��O�4�I�!~U���U�ZN�Q����pk�f��Ƈ�{(�8�����}���v��a���X��?���kv�����'�~qF�C^��s	�qkT��l�z\��H.���*�w`M%���{j���	�e�BJ�a8G��;+!�̡�4{a�j��}���ʖ��į̀�{���R�Z�0V���]�Ȁ9N)�]9��a��`W~F�S�Ƽg�� S�NUKP���+Q���o:t����$X���5��$Ea��K!��Ь�̲A��-	�ٍ!�6.����ǈ~�*�3 *b���ʰ�^f�o��</��|Wل]"E�)Q'�\\�:�\��f���H��ww�m=��4��A��5�a��O=������]E1/�a�X���$�q�����QY��w���7���<��:0�ݬY�}}��d�mT� |̜֕�t��� H��R�P��&�U�4�L�er�'�D�:z@X��ϣڦT���S��&Y�������j�/[���ZD�6\��7�e��1
��i[�E��|��JK�JX���egt7>�-�t�E��k	���h�Z� ض��^���dcC�ȝ܏P��x����.��y�RZ���y[����EwX\+u�
&���d�<������4�(Y��ڡo#o�1�>��d�L�W���@̓L�'�c95#S�;Y�r�!�=����Gw���>�y����^uPኜ��<5��W�i$��l��&(0/�"�*ȩ�@͎D�ڛ�{�+Q�� ��7հZK`�iwi�f��b#�K(��?ч�+b`
��!z[��]v��Όd޷�K� mq�6�e%m��m\����� |��S��e�)I}b�2@�^ЃVy؏��ĉ�i._+���Q®��E�DjK�󀮖R�濶���I�*ȰD[V�@�R�M�a
�o^��$���FKDo�MkJ|K�f�k�;r6�����º�l�\R�l����-Է_N�����<���zD�k�+i� ��[�O����='�u�xc�Q� �����˪iP��U/y7��*��τxy�_)��"�/!k|��@��K�����{�68�ά�˨���Q��mF<Y�5As�Z��p��D����Ϊu����HY��ə+�l�7��|{e�(j���Ӆ�]���2��k���S�٢RM�8#"RS��g���9X�,�����)��4�٠���x�iߡ~-&MY��ӥ�:s����zSk���.�Q.Ŭ���Tk	M���MZ�g�����1���CKs�N�?��g&�|����R ����6�ҥ
4ǖ�`�h�q�4Q�x��.���w�"���гÖx�4���1"D���n<�+�ŧ���H(��s�kჟe�Ο���%ۃ��h<gmC��a�eu��
,b�T���i��4.��M�\��ͤԞ�;�Lڟ��iD�6}P����y'�bD�P5�˼��:FG��f��J�z��������06�����>��mG�T�^�֗�ف"������d��PS���X#���W~-��ޭ��-w��B0AEh������(ƌ�8!b
����T�w��.�aD�����J>�`�3䭌�)��WI�(��rNZ$^�U���Z��Ժi�֜.J�S1�Qu+�~���`~�-�^m�����p�N3�Ch�|�y9���ܴX&��������Y�\0�j �f=�L%��(�h��S�kr�c�w%�c���L^Z�+u��l:O؝����t얨�b��'�ѩG�B�奠��]G��臇��{�wJ��v>�D����R���8��f��B�}��KwڼV!+�"�:t���J��eh��К�*h�f/M-�������g�B���V��d�G���]�(|+�8�X2��W��}v}�țWs�)�hJ޳#d�5�GuHA�Tut5}��1<hop��((�ҷ��(fN�������>�8�l'@x����6�������Z��"��I�r��� u�Q�U���\S!�ޅ�����+�W�A��H�;��Ml�o1թ��!������aچ��F$ܚ�-;t��Ѷ���82�4P	C�,�A�T&���lܘ�ΤO�[�Ŝ�݀0����%5���bFğ�P��R�1����(q�	�����b�<Ϛ�!}�+��3mR�q�V��	5���t!W�x61X�-w|hxf�JZs&v-f�^�AT��A�[~�Es��]�sFbf�q�� *V$�[~�;���L��������J�	U��N�D�ѷ��F?��뤁_t�Њ��փ�~��N(2���VK���+.[-|�R��'��B�]�Qh�-��DL���ԋ$���޲�:F^� ĩ��:Kh�����Tm�3�-��SDWp%��X��y����Q�d�	/Ox�EoP ~�0Q�\.�X'm�6��ϻ�?H�1�i�~:M�'�Φrӆ�2$��> �f�4�1����!8��o�aY��o ]��dg�(�ĝHn.4�����P��*��WI3dz?Rv�Q�Q]K�-<���HYo��x�\�i���`d��]U �h�'=�b������c9*�~��Y	gϬ�u��H%���1�4�j9.��]�S�/
��g� �+}�Yw[�J��Kzz�-PP��hO�n�w���E̚�ָV^���፤z���T/�.&S�<���^<�'r�M�~��̿�"՟A:����=D����1���U�6{X�X\����)~�Q�#h�.i5�)�n���,I�:	�Z��P�6��~leD�o�4`��rЕ�O�9���t�l%�V�L��C��Ջ���I;�3�c5�i3�S���n)�L?�A��7��;:|�8FN�}��Ut_Z�_�B!�&M�dz��u�m8ͩ�sb��L:�����?�%$0��5{�DC~=2~ʬ�Q��t@�\e�etƞe�#x��E�V�1L�漢9wr�4�'��"ؙ{��I��C9��������|C��\���TK(,���E�@ �jf.�Y���F��_w���^I�dI����ֹ�y}��;��kO��7��6/8���?I���ώ���E��Vn�gK�Q������%-P; ��jgQ��E���Ћ�>)�Z=�4���+����V��v��X^��eZi����&r/^x�Ð���~����'�
?Ӹ�⌥X�/`Gd�,�g����!�x�B	w��ː�~���w�!b�g����!V� a0��&#^Eg�P��(N�4�����ߕ�k�="k>GA�>��5){'�pF�B���g��=~X�fF��61G˞�_&��ܱ�3b[ G�Ʈ2��(ȝ.��V�U���i���,ϫ�Elt�Ԋ0���花rd���2�,E0}?ɚ�,�[#�m��F��}'���\�W�:���Q�Cmd�e�}I&\�4��=�"L����n��?�b]2h9jP�  L��_�+�y��>�k�1����2�	W��O�����9�:���{����,9�uƲDc�6�+��W�˴ ��,!��J�z��/J��-˶�i<��r����mw�8!d��p�S��g,�ؾ�k̶����d�J�����.Qs+�ꚏk^��k���f��V[i��� by�n���cwMSЪ�m/�nv+Ig	 W+�	�U�@�cQ���h��$Z�p�hf��nr�[�f�+J�3��%�,�@����b}���0�^��j(�I۬�vf|�VA��u0=h�޲�tLc�K��M��խ!����� C:�	�$�7�1�4ź�%* q�M����	˲��5��+��7-�MI��Cv앬%�pH7��S���_Ⱥ��0����uKO�O��c���(O? *����%��v]e��!�m�B(l}�rl*iby�-���H��j'��X��>q��|=�J!�� �Z����fz�ȁ������0�"'�gy�����P�*�|�_�TIL�1�P����'Z�Ax��� Y�
P�A��j��I�e�!5�,_o(�=qn�w��|���Iϝolv�п�:D���d%�9<��ZDD�#N	�a��W
��3�p��+�_�������g���:	�l�˰p�l�����+���\����:z��{�4��,G���%����lьa0w������F�`�&C�<�~�lr���g�~{��:�^( _�=8c��s��*p��v}h$���G	�y�~�D�� ����ㆂ�Uy�0���_�E��P���/~�~x�`���&�#�_=�2Q��WvH蘌�>>���g(`-��������A⩜����;�Du�w7��p��Iz~8�Yg��j�� �hp��Ѷ}�N+��=G��A��F�C�i�%m>�ev�U��7F��C�T6ۥ $Ŧ�EqN��lm]��2Je��g���SbV���w���r��q�5�J½I��H��D��F��
\߶�u;���3����l���UZ�xڂ]�l�I�a*4{�m�����T־� �n�?��W�#�Zde���{��3?\��(J������h��C��N(tXJPf}Z��y;���~_t`��7��8�	g��M��N�6!�X���Zӕ4�� ����T�7��һZi���gN��ߎE�,��ɨoG�ݜ3�������?M�X]�SIId�
n�v^�m�� ��d������i��h��q��_O�3Bص�����\b�}R�z҂)����>ғB�{-v�o����M�aqɀ-W��>��LH�E��3Y �7�M,��2^ȟq����хt�Zz���m\`q\�r���z�Jj��G)�D�R��gHk�0
���)<�"���J`u�p,��b���[������.�T6�"R� Q2���O�x�Ål�C�bFi�F�ދ�N����B��9�"�jt?xQQ��{mj�𰱘��J�h���uD�5Fݱs��K�<����d1��ǐAdql���sE� Q�堨��,-���2�8<����y��N�E�[6Q��9i�m�9��i!�����L�i\�ӝc���ܺ�3�p����l͚#�?A	� ��]��q�-Ό%ț	���@�*���|QU�>�7DW��Y�[}κ�}S/+kص��%���S3�?��Z��//sph��Au+�>�4qU��g�q鄱��I���ۧ�?^4��[n�P[�<����D��F�*Xk�g�;7�g3MY@"�N�Ђ߂}�b�=��F�Q���q;�9,��%�L���|��56�Qze!�L���������W�b�q���_234��V�B�&�yʍy��3:3�����KQq���k%R�;��|��Ϻ�,EAt��Tب�2�U��| � f�$ݞ��s:�,9t�P��ƈ@��9��Xa�K"��Ls�ɔD\h���VK���3L�vu��4���8��p<�KܞE�z�ڊ[�*�����~��~ȾEE ���[!eD���В(���%&�Z"#��?�xjU&I����"
+���S�1T�d�L�	@�;���G�T_�s�d��q�l���p��jP���w3e�K��|)*Өa>!n_r�eʟv��vNd��ńu��3.RO~�݆��������3�,=��	1����z]�Y'�/ZLj�K���p7~g	��%��\SF	��a�Av�`��j�r�t@����q��pW�r��}m��ɿPr5^+��R������5� `������g����~���N�O�"_����TQm}�I�9��`�[d�T7�&���lԑ���A����~t;�am3R�1�&������Q�/[�,R�ܿ�r�3�'n���C+�q�����Nc�S��F=mȞ&)ղVs��/X��#����dG��J��IJ쒔GcP-��o �����yۆ�v]˴���7��(���O�����o7-?���L��dK�*k��o��@����1�`��-�S��
{��yN�pT��e��þ8�"ƽh��B�/n�0o���!RZ�5��]{f�D�PvzR-'L��F>������%-�e�"P��ߵ)�˖|y'PҦ)�מ�+���)�&� u��(Ӆ�T셊_Q��~E��! �g��A�@�y��g�;B���r��jxw����_ '&e�p2D��b�ͷ�����7�J�CR�L}���H�M�<0�ɺM�%�On]BY� ���69V�̽?�2R�w��p+�嫷}��)܇h�8�^-�W�����' �����c�v��g�����4`t��-?���:�H3[���U'yȠ�1�
݄�\�RH<��g����Lg�0������,��"7�==�;dc����({A,�����~۪m����-�Rf�>�H��_��/���[���\!s���)~����H2��wF�?��]y�0�-Z�\�^(��pc܍7� ]r�O~�S��\��EFc�tÞ�Rs�1��R�n� �\��T�N��W������>i`��,KwN٭�$b'�*m�8d����-h�����8��4鿕 VMa�2���^娌��Rk�F���7`'^7�0�-���q��qBR&��Kf�=��̊3�����8j~����^:uד-w�O �C�n���ϯ��xq����u���4�PP���L
��fm4���a��&��;RɈF��q8z���� z9�E�Ծ���?ÈUfo�iEY'H=�Q�ΔW2���h��@/<9�A�?��w���FR1��M3��
�^��������b}R7��������Xb~�h7ϲ���bw�?Y�W����{�0��t�������2��O���v��	�������lp�\�������#x7�(���֞�v��	�\^��KrWu��} �LI�����o�����G���m��d�R�l���B�'�ߩ�f���gQ�a\��yZ�qh���Y�-Z��&�8XB���,��|��B�,�?U�'ͨ�A�Y��Zj��>�ߕd�%ؤ��%=eaB�zqM������N�(��3�7�v���b)3W��Y�
�L���kX�H�Q�E*�._�q/uW@��"N����Q7��+ ~��$��0|�!��ߦ��Ws�Q��],�(?*X�#ͮ S��	!a8z@��8���]�/�򵖜�OaE��i��o���Q��B$��*C��1�����)��A�u�17�G��RJ}�1�!or�������Q�1����U��?H�Fo.)��\���2͑^ Nt?ç@���@���N-a�Dd'MSql���] w�-�;���`�Z���sBI���!�/�w�������������U*��p� Gj�h�y��q,5��"���)} X�2T!�_+/���Y2���1*D�
��`��9�	���r�Qs��fN��7��T�^��s�t �L2�%U��B�ubD������VB��|�����������G�%�(�/�`�]#TA�m8��a�Y��Q���/����Gކ�����VB���eiʆ3>�d�?�֭DcnF����n���<̰M�`><mw���G�rO�Q�]��Ɨ'��� Uԓ D�֭�[u��)˼�H���}V�0�΍!<�H�ށDK��,V"����w(����3dR�q��� +]��Ƅ>1�n��W�bnYC��O��4��Js4�f��o��J%E���H����J��SA���F�!ZU���4�p��:�@_�Heo[-G�q�F����+Ju��r.;.7��Үo�/�F.���7�~o���/q
�Zn]��C��
����ݼ��^����s�x���iy��|.�ڂm�N���B9��z"�,d��v�^����� 嗑���f���j
�_J�@I�띓�;�/�\͞t�&w<tf�D�
���qy=���̗���Z�*������8I��*OI"r��[d@u!1DͷGe�8@6�� 8ح�s da�Y�|�(�U�k�-\��ݲ������"�' -r 5 ��)����K�?�Kg�pr�����E�;���U��1�����ӳ�&��.އ�:H���Y�^U�o#�\����H�֥�V��Μ}�b,1�M�fԌ�'�O�q/��hz��Q�d�M^�g� ���3�#��Q�����Vaۃ��3$(G@�2��Ң����>����!܋�ϋ�͗�u�]��`�{y��H�d����|+��k�ҕU���++L�����ƛ�0�r�0=���M�A��}�*��8#ǔDVՍ�u��f=�M��d���l�̕�x�kCXm�$���rr
1�g���V��Y�fs�a��3wF�w.�@��Ə���kI ^��>RH@�5�p�C~f����:�Λ���k��bSi#�L��r�dj�&�o���S;���y^?7a��m��Ew�6�5p'm���a��ئn�^��
ߔ8V���g���D����T��;��L4�.�L�|Q�Ľ\�@��j������"�����L��ɛ� �
ʥ����w�n�p����6�Y;s{@��	�1օΑb�ܩB�k��⯫r���_��I�%��v������lp>9�%�Hd�C&@�<����>�6���8e<8 �ݣ��'���N���B��:�O���Dꯈك�g��~�N	��:%�9r��0�4���h���:��C+�?��ү������c��lS�of�GI)�9������X.Ky�sV^�гo�
Јn��N<Skᦪ\t�Al<�W-
��YjC �G��4��]Z�������6>M{Y�^]8��E�NVP��t%8� 52� J�RI��{�sv|d��e�v<�!�y�߈h����L�A�٤�x��Ԫ���U�����Ek�m^<i��*�����rzg�;�)e��j~���dL
�f���i��y;O/b�*DC��j��j�p��R�!��~��es@e���N;̮�f6���	-�o�ř���e�d堻���9֎���c�{-[V���j�IQ�7���ҿq+���`��]M��\԰w�Bn��D����^b�����q�?a˚���- �"�����&��oOb�#v؇�Szt�
蕨��W�[N��zTUOd ,/,'q���
v�d��cmo�f�3O����&T+�����BI�ԥZ�c��W����g��ص~���X>|E�3��4�'�"��23��5�j��O<�D!é�6<��&��6i���U���� ��<��.�.0�A�Þ��Ļ�O��R�p��@6�ޛ�Cpimo�m�&D@$v�-\j��%42��f�.?��t���E��[��{�w��LE�p�x6H:E�Ȱ�!>B�!
f�⣸������F��m����dX�"����"��$�P�C9�͹H$���@�M��d������uo"��o��	]��j"�D������J��E�H��OR4	TU�3'{P/���ĩ��g"�A<ECaK�J8���.��x>Έao͌P�YXJn���v!���f�'�S���5w.׳���@	Y�1Hڱ�v�!�`�{J���Q[|�O�p]{�'���MW�8[�a��!��>2��Rș�'�p(	�^ە�`C�k��������`����������s�j.��I�����qu�TA�(�&��men�C��X�i�	��6{f�=���:��)���.�{��吣R��/�9�=�[���J���V�@˸8�5��/W�U��T�I�V<������hz0a�opO#Xл�����|�X�f^��
ݐ�{�?f�IDo�TM�sjxX�ǃ��=YV�����8�)���I'�
3��������0H�?�4��Й:��j�����'�!:�ʔ���A:�?�P*ሡC���y�<��R�4�Ǥn�J<�!Iύx��
�n7L�rp�琫|@xwi%�f�S>2��kq�m#��c7��7TCNZ�A�+�y6	�u�Y��p����W�Y�~��^�ю]?!��L���&tL��ҕ�&�2�I�Ο�E�A��4�J�_op��4���My�m�H�H |�LΡ�t$�̣e�U�e*�n��)�� ��1���|�1Զ���]�L,.���bz�a���%��,�k����1���.F	?D� Ԅ�l�᪋(��c���ROi�TN�}�YC$��D��ι@�L�4y"����J�u��L�%z��AV��@I���)r	�?��d�ع>"�kg�$��o���>o���G.�&񑟕�v"I`�V�3�|�g�h�I��//��ZE|R���3bI�c��F���}�g�ؑ�dk.���Il���gW��9�l��Ր/��Aȑ��t�᜞M����:�	�U���6�rФ������e��f�W���aP��ı[���*�w�5"1���~Z�ud�V����9/-*�)z��)S��ێ���{���m`'Ԏ-/���30�^���9(�-�a����>[yd3r�~�0J�a9 "�7TH��X�1����
��m��̟	"u>�Cy�q�ߴC���۲�L�.�3o^N<�7���!�A�)���������O�	��P��s�����4�:%F�46���J)N�h�9�)�G\�\�^��0���X�H,RUyP������%�������h�����-�}����a��fИ{�(��u�SU�� ��YJo!�#��� _�,�A	20�ȣ��R�0��[7�5&s�� ��bY0�����P k<!��,8SM�����IrYO�a�����oU#;��1$��t�zZ~2}ƚ򖊈P}��R����c=C�&�"�E�(����\��!�[LT�R��q5�a�?���N�X~/�(F��v�H��3�h���c{����� R���E����񔮕�Z�<bk�_���=i�����������5�a�3F`Dќ�S3�̏$!9q�bj��/;��Գ��H�/6���ڔ!���V,lS@���!x1r��ĨH�n�j��]���8U�R/�3����2��a�!xvfΥ>���j�6=	!g��$�%�S��m��02%ʑ�s����Fٸ�Z����O��*<՘r�ތ���'�e^�LH&��_�?џd���T�?A�9sW���*,�^�>��]\����Ӗ����#���o#�E� ��y&V2e[�r_��Zb0`N����G5v�ƫ=6�G�H�,��Y�i'M��7D�'������a���	��D�E'XM�ml�G� ���6@�1'B{&��j쫫�R�A��M�#�ׁ�C��I�J'����V߇�����b�o���4�3��MVh�R�.S����z�aʂ٠��&^��(��BB�]��W�;'���͔�ޣ�ů����D��]	^��>�,����e��
UҤ�AX��Vk�A�S���d�'��U��\;)��k5�م����kn�t�P��ϡ^�)�v%�єӍ�SC@_��gpd*Ԫ�7T86��Oǂΰ���u6<Ud�̑�ӆ��)z����:Fq�.��z�>�1�{[Md6%���ԃ�VrS$̾9�Bq;28��^y����#��򞸩�j=�U�U�����YQ-%{*�8VӍ�����N|�s���ט3����s>�n��H^����Ѻ�;"�+ur��-Y�$m��0O��*��A���7�ROW-V`�����qy1�4eO*>%�<ؘ�/�^};�׵뎐��q�_�)�W�842��^�d��S��*|�N�θ�: ���9��qn{?aSsΦ���N�ڨ���>�F��� � ��\�Jt��P)�jG��8�Ë�L͘�Tq�����$�R��=�z��7^v%7�R�i��p��Q�Y�Fc�G�9%xp�&�%޴�a�Ar���2����]����@��c��?�X'n��}wCQB�> D5��K���������P_9�o����#?����l����6��%5z��o�T���s���t~f{�#�Hc��\�tb`���X2���g���F@�F$�l�����Έ.Z�_r=�e�M�!͈�)K�͉�ҳ�#uw���ER���M��Vi U��]��b1����w�A�g�I�����
��ҕ������t�OJy]���+Q#g�u��y-7�>��n�~T��- �>؜f�ޜ�!�8��kk��/V�.s-1�Z<b[��N���bѪ���MjIP�T����jE�e
uG��)�l�w��
fsN��L��B=EQ�-�<���EN��Q��)�DԚڰn�^x�����6�A�մyp��S9���{��G�b��c����~�׵ު?P����L��d#>|�)��$���~�����I�������'cCsx&���S��^�̩�:4Hn�fA�A�1�A�k�(��^�&k��0�|B]��͂Tt����Y'K4�PA}0��M\�& !S�?�`���61"K*�']��L<��HQ;�?9N��yl�׽v�x\L2[�=�I٫���5�}�}���`D���#�53)�� ��t�Dh	\�U��2���y�IҶ�W�P�H�� &[u���G��)4�"�A��6��������_�_%eڂz�U�#?B[(��k���7��z�h�������&w�sKMeiY=d�I�y3����|z��n�Z��*1@�	�2�b��_JS�x�`0i��Cq.���k��[*p$k��X�)"�k��Kh�-Z��R,.SR�z��0���M?t=�U(�V�i���~>�0��_�(���f�E2����*i��oAG䈒*#E��bɂ���V9�`��8��$O���!�	��Ί�-	O�WLF�Հ��<8�R�@;�Y2 ��|���M��_�u���^�f�B߄�ֽ�'F���$�?6�´���V�����N�f���>;��C6b��I�GH,�u5G��g����A�x+���1	�UqpR ��n��{r���Z�Q���[�/���O�Zw0���QRn+5��6"���=��2;�'u�\w�ޤ��t�52������R/�oں�h@f�3ٔ�KZ\9�3R~�O��B��G*�R���C6��^�<?�i��;��@$Xоis�pG�gz�����%m�J�J_l���b�)=s|!�'����>����%�k���"EM�=~7T:���I�^M�B��	H��C��y����P���.G���*8��᪠��+ڻ�.�� ��R\$������D��ָ-۬A��u ua���~�3�Ǩ�������b�r0΋����-�v���+���ڗW`m#8z�3+閕� �w���>,������<���� *y��;4p��c\C�0`{�@��Q����_+)���D4�;�>���
��i�1)��|g�G»���=�Ec����+N3{9��]gaK�EKj���xz�.n:��|;���W�K�w	G�5�%�'��kYha1±������*}�찞��Kq*,��u�8=�J29���ܰ���1C#T@'E���@I��'D#��4�.����&\F��A��ɂL��4\Z�o��ػ̍0�X��6Xk!#N¬����nB�U�+��y��'�ا�k(��*9�r�a��Kԕ�{|U/ߨJlBz�P����T>-J�K��r�s?�8�����cL�Q���K��)�����m6��N�mp
����[�4��c�!�O�.���Rր�����CM£j���)��	�n����ss��5�,�7` éX�َ֛냌�?֦���ɚ�g��/�{ xZ#i��%����S�M���у��x�0�d��ɓ`��u�g-?��C�e�pU���y���N��V �ˡ��<��B8�)ĩ�T�<B9�?R���$�����ܙOZ~iϯ���������_W��q=
�����pC�ǀU��=�>�M�r�Sg�sIL��΄�%��S��-v!1����-��.1Ϙ�р(Z�W�?a_MMDb�O丫^m��@��SعQ��V��m�L��Һ��O�)��9ϧ�O}X�e�d4԰���E��i1�Xe-nJ�r����xh'K.+���q'v��v#D��$�E���}m�����ʂn�T̖��i�!�ǲX�R�"C��8��Q���1ak�F�*B��E��x�����ӋFL���z�b:�tL�ч_E<�D���>R�U2�<�PF� ���)��e�n-����@�>���2���!0/WZ-,[(|�nO�)l�0��'�u��p�u��1�,!d��,+��x�#�-Gak�v@�=�`��z+5�	��K$��O(���;Ϸ���B�%!���V_?/�Q����Vô�g�P;R�*�����O\�"p'`J�t�Lָ�`�V���˝V�v]t�v*�L#)P{Ro�� i�#שz�C�s��4���Q�a�\�O��`�D�.�{�]f��z��P�DwR7IҾ�ڙ��B�!���̽9��N��L�}��v(�.k��O=� ZB��C1@�̙�N����U��y�5���ٟ�2��C=��f0`�1S#���?R�H�H�Fxr�r����g�q�bK ڞz6�	70e�<F�q��bƂ��3{v���Q��ac	{:H��Y�G�)	� �Be�K��>*��a6_8�Ø�=�C,���8˶�����$�������7�$=������'�~��1�}��e�6���#M�����F�[�G�y�H  ��zKk����fQF�J��#�W~�����%7� ȠA��TV<�}E�X��
3v��҂�v1;u�Vc�t������V��rN�-���n���Fӆk���w}-�����LL�Xh>;n��s�����l��+����h����#D���k���>!^5Y[Bu�$�w�Pi��%�, ��w�Z�WBw�Bj��^�lV�� ��23�	���m�@����?l�6,�D�E����8� ވI���t�nO���p�/���'�ޟk2(�P:�"�?K�r����;��O����]og�>�*���;��^#<����;�����uVa��B����7�w<�%0B����f�1� x�m4�g�����Ap�[���E&VR�^�!�bz����&ß��5F��ý�3%ԛ��J0���6R�����ۆ<���%�,�T���~��T�U���"����}�=S�uK��Z/jҾ��
;���_��0$
L����t�2�4gɥY��M��h<`�q�2��������-	}����wz�{�r��~Ĉh�47iV�ku�~���6�����?��Q;q��h̜��/Ij�Z��[� ��uy�;���q�����������[>��F�JK6�b��`��)����B�����&��U�p"�0���	8<�)�;�Z4Fl��ﾪQ�˔ǔk�"�j����A��� �,�#��M������B%>N`��˴x1G�W�6����F-r��^��.)���rIF;���❫V������N5��X���$�I;`R�.���(ט�\���1���@���qB���q"�
����P�+���]��*s�s-���@���ל )'�EH
*��v���d�� ��}��� o[m�s�z~���b��O�Pm'%�}Rs�Njh��Hfa�6�Y�}4���sTŰ��k(Z�`Y v�_���7IÜ�kv��cW�O6���5�a����Y�2��)RњC����F�9�"G���O���UM�֭�f�;�U��np,�3���.�nHs����Ln�7�A/G��;KGXx:W���M�j�C�.��܋�@�`��|~ ��fq�]���[l0D�j��	>�Xm�a;���-�f霣A
��_Lᢶ��b�8-ġT>���\F�9YS��}��ܩ����&��Z��icqIT���Ou���T���u��d6�6	��/�V|u����f�� �}ϩ�nIB���T�r�O��q�����[;<��NW�jÙt
d饁��<n^ª`�GS���Վ�mDiܘ̽�'|�^�H�O��م^,��q0D2ʼN���V����e�s&�M���0lmd�K� ���?-V�	�؆N��0��R�u�+�[§XjvǝL%cٸ�D��qm7楡��ϡS+��V��:����Ph����}�>��_q�.	�� �Z#�V�X��X-�fʑ�Q�5���3�T����`���昡r�N'�?p���g=BJ#�W%���:��~'��\�������zQ❆~����8��o�����u?��LK���;n�v�$@�L�t�B��~���S_�e���$g��h�4��@�zT���
�.����!^i�
"� 8؈ w�xH����:g�$-r�����=�[2j�0�}"���/�M�FE��w<��q@�g��Y|ESp�����UJ�Dn����UԌD��}��Ύ�"����ɒC7��>��nn��s����ݷ�/���g��e��-��݌�=��Ŏ�.{Bm�(�?���@%D�O��s��nd���(��l���4����#��ղč�S�^�����5�i�WQ��!����[a)�]��-~�3��pV8��c�('��^&[4�*U9��(����4*�n�&�+ ��n^���x���FZ����|�TLX��ݓb���q�H�����uGm�^��5p�Uk�~�!�϶z�AO���M��;�N�b%�� y���Zc�1s���~;�:i���� �F�����pWmUn�<��p����,���Og7m�yy��1�J�_������_�/-�7���J��R���#:��3�Ym̥9�����%���)�^����r-١��"i��\syMǔ�%��R|�+.&.z�����8L�y^C	��a"ʳx�J"�r�%�$�jQ�a||��?H�����Q��=w�h췹!�]��$}�?�ydlx�f��=�z#�#�`z�x'ؼ�l�!$�n�8h�Ǵ�߸ՆO�v�&"�K�R	`�!a�{v�NN����)�O�K	��F��c2[&Z�k����Y�$]�����j�^Z#�T��ݘv@���xr��	3��'��#o�+s�c$�O�<������ �bY+�'��v$p:�m��0I���v����?���x����.�k:B�D�<_�_��	��ꀧä���蝷^
��۹�U�k�8;�<b��,7��G9k�rNw�O���`���e�E�d��*R�ꬕ�i"��x8V�m�`'[v"=X���T�p�.��>�5���\�cL`<�Ż��w8�aw%�#��J�YM,��)A=���ё40�yg�I
fG&R��\]��2�TЭAF}6��,�b��{�k�a%��܎
'5����^�e��O��Q�)7�2`#�W�}-*�bh��!tĈ�o?�9_�DIr#)n2���r�����Q�߅�PF��Va��2��#PS5f#��=�ĥ�Vf��C���xԆ�' ��x҃�5�ѡRy�_�u?�=����~0���"��s����
R���G/R�C��<,�W�1b��s]��u-U5#/a~�f����_�ԭ]�#�$�l��E��;�mC
O�x)��@��e��k����)ز"�@�˲��Y*x��?�y���ByXlsَ�W3?��mڀQ?���J���%���@	��v?�cR	�ᢖ�ل���(�TW��y�R$+�2�/��1�34av��܋
Ц�n�����g㗙�4��:�>�����X��a��5��Q%ž�ݴ��8O�hccW��~:�ঊ{�m"���F���|m��#��3�~�w�L��.<� ]⠤��7�гhԲ���$�#��Bp{�cT�m����m����&��o���_�4QĚ;��̫��w�a��ҒJ���bJuAz��q��K�2�7.�D�G,�_��Vw�
�?�|�����Ԏ�w�?�`��9�dk3����#��w&
�p��ǏZĘ�:�gB���R��ߐ$י�]�B^�(�D0N��+H2�N�ozG�yF{A��r+��e�iA�]V��'��P?�#��#/�q_S�1�O� fA�<��?0�'8ᒚ[�p��D�h���$�.�{�����j��S.ͨ�����9�����߫�a�ۻG`����qe��w3�D8N�]wȃ�゙B�<v��El�o���L���<Y�2G�G�}J���?n�}0�� �c�C�>�đ�:$D�Ƈ����`
v8J�䲏?�pgb�0Dy�Ov��G�m"�cMm��w� S��O��Q4B^�]�+m�`5�oCA��O��.*�;B�f���:��|:�7��*_���_g����5���-O]�^��"�W�B�_��X�s@�q�^�@���p����XA��M�^y/��.�!n��_�o?,���y9�w��JO����\^n�|����v�&^:�_W��˴���A�١��p��[�Xo3��%t�I.�|`6�Fđ��J��KM�:�'�+@?�2�M�>�9��T�Bsq@U۰�� ����<�(�:/����E"s�G��X�XH�4�T%����tQ�O��	$�YQ��J�䱼\�H���1���q*Le9owY�mf�%���U�@�\Y�X%Q
Ę��߅q~۰
%V��d�-j�M����̌�y\�û�t��_��]3:'� Δ8��+�b~�7)FY�Y���rjs+n[M�&�rq�;��i���[]y����~7��ٞ�X���0$:�D";d/S#B�6S��|~���Ж��$��p��(y�/��������/�s�	&�u�1�;k��ڙɼ����B^���`;pM�'���3�F�m����ЎZ
����t[o{u"k\��� ڬ��W���Q�L� ?�_���5��
 逈�b�>����-zz�����m3<���}Xۥ�H��
�&A�8������5_�]"���4���q/���L��8�&�VR��aI(T�F}մ�b�j�~�X/�Aҕ�+Jm���}�����Qs/ew�x�f�SND�y��	��{m����P����$��{4�؊�*��W+ύ�!rR6N����!�\4Tj��nXՖ�KnZ�)E$ǈ���K`��D�"���)�(r#a=�$�J����.�^S���|18���+Q���YvG�[r�=êdI?����f����6��Jl	����)�T���f����ekx��Nl���|
"z���n*���f�;���7��-�����`�*���h�uU�>i���|߳�uI\Oѽ�'
�7������?�%K�:��N� Q �$(Zf�<�1�)5;n�N�f�.���:�C��?*o�F#rL��Zڭg���]���ĺ b����5jϹ��/r���d��O&��!�
���0�Z��	9��䵃У���z&/cH��M@)�I��:3�"����p^����t��.5���`v����3��`��b�s1����fFZ���"*?0l�d�TbI�JўOy�mA*���)}��Lx��V�^��Q�_�O	�*�,�6��=z��H�
�s2�5*�%��Y+��ac�-�)�&��<e�Eʹ�N�x)8M�v
$P�Wk��L�8'�l-��E� ��c���<�䙈0��;fo����Wc�P�A�nW�9��,������"6JJ��E .nA���q��`-��:;�'�����V�\���c/�bR�3FZscWyZ��4-	���l'#kk�u����0�S���k������햱qm���E0N�:D��$��pS}��V� �&d���Ʉ���A����;Ͱ�g{8��?Y��ꁗՆ�*V�?� }y��3AU��x�
��Dx�h�cy`���)l�СU/����έX-� �ø�\�O`�j[��n���)fI'�b�s�v���Y���xM�6��뤖�d.znA/V�8����D])��`UUt��)�{���I7�d���霈R�RS%��J�G�J�N���b�������2�$�� ����#�oq 7��Q$[���g�f�𺣚�bi<�h)�"�R�6��!z��M�ȡ�	�%�R�x�-Y�K��~AM��u������ᦿ�~��
��A?�{�����Xf "�<�)�.�3���ƈ��.ZG�6���	˪O��|��e��f�D�s��Pk-�K�Q�:��%��=��'�/X�� ��V-�]lt�@�~yw��%����ך�ی�����W�G<��*ch�0Y�"�0S,�WM��M�R^	�� �����v��8C\���e)?&:P���
�i�Бj�)�"B+����Ĥ��.t#9麕偝E@Ypc��B��a���u�K���.B����׏5tڈ��z�y%Z��4�z�r�Xz����|�F���6�yŪAj���9y}�A�{R�f�������C�]:s�f'�a��֕Ի:T����K����9��,c����X��J��|ޅ�y>��b���+Q��\��]N�.5MA�(�)�T�b	cU�:�E��d��RQ6���I�8 ��Ǥ�����m5Y[���w�窭/��ῷ:�k2Z��.���~����%��?-2X�5�)\3�a]@P�Tyv_�c�	`M���BhLV��S��Y�|m���L�n
f<
�Y��|�����+:s��ɾ�x�Ƴ�h6��v������%ଢv2s5������*��Ht�&�>�l@m��������k~�"���h��g��5�����Y }>K������؟e����?�4ԩ�Y�n�}i�}����|����dF3�����GLq���F�>Ub��3m��h�1~ئ�5+�@ ~��P���>��X@�^��1�m�$6G$wEHK"՚�+TЧ����:wtH����C�c��!r)С?P��09��6��w�rmO@����昊�z���f_�pq��Z�B��i�!��9&@W�}Xf���1���\)B�l�e?FKӽ=����!M/���g�3B-F|T�u�GъYh�n�,ͱs���Q�oK���҆<�F���-W�m����S�j|)��[��߆}~ ݪp�V:((=��h\���������a�q��%`4�>K��)墨Y�$�j2@�����I1.���V�(s�>��N��F��Y��J]]\��~%��c�>���U*�Jm1<���yW��`){g�U܉i�����sB|H7��\Y}��� *�V�����^�F�\Y���P�x��F]H�/3��d�42�d����c�
���;)��AH��ެ"��"��<��M���?���j�?޴4�,�I�%�V�1��3{�fNAs���k ��<��zw��8j��hG6c:!�AE�Ch�����|jFo"��x Pi��,J����{%���1�On�C�o.ڄ���h����T�X�~�4�/R;�2}��MOަ&v�.	g�E��k�;���[����?���_N� ���O�M.���-N��2E� ��7t_|�v����Q����F�C]�B�V��ȭ:���,e��J� ��W���^�5���	��#ʪr�W�#o�j�3�{�9=����fF/W]b�AP� ΃��T0 T,U�}��8�T�ޝ�:���?+=/�4Ë�#����	5
�7�@��-�m�A���c�ݯ��"H���R�A�[Σ� t��� 5��lc2{д���q��eԏ���h3��!��R+�W_$���.A7��	������۲���\��&n�����UDL	͕D�������
%9Ĳ_C�܀�[�������S��e�-~^-t��4�!����&�!�1�K�Z=���`z���#:�h���M�MK�(�ħ��|\�$s���q*x�>�����K]�6�B˚5 �4���!~�̴�u���t2�^9�Y!<-�

@$�uC9�H�kX r�~� SA˸\���U>�KV/�a^�Nz>c#W6�n+��N�G��ⲿq��8�=w����̍�.f�͚���$]	��v��KU#q�lo��*�@�h�t�S�;<��6>nz?6�k-b�ak��,ǁ=C甂R�kH�f=�IA�'�2�&�z���?�Pa��F�6��Py�
��i�&��T�3�<�Ѭ\�*2�[8����tO��ʟ�Űt��m��r����R�O���?�|0�� �����C�'�$?I���1���hm7m�Y�B�4F!�aa_��%Vj�84Yb"8�u2�J;�8Sa��}g�K��(�q�ݧ��������<E��瘫
S�Μ��-�~�h������=�h�����U�1p�����9l�����=���慺P�:���z�?��)�vw)R��l �C��6R|;��S
@�7��p�Q�dc=��|j�P�[���~{�����Rz2t�}��vk`����g�u�lm��bj�K5m�O�T�i���v�;�?��%*�-��bK���r���K�DI5���
t���� �#:�pҼ�F�J�U�	�맲��{��ӊ�.n���@N��\��@�v|�Ҹ��+C�ho��Fr=i��	����'0Z�V�R�
�sNy�E]%��D�Р�B��L��v-�J�K��T�	��� ��p��E`���m�b��� W����_+�`�7b�Y�Z��ٓ��g�.�yTdc��b�5O���j���tyF��]����8j5w�y+�����jP��.MMf��v�T��H��3��v�>gUK��ַif(�%�sH�G<�lk���R�U/Ռ�Od<l8��c���R����p&��V�>���c�.u�q�J�k��g�B/A�d��t���+��e�6_����.ώl��deD�ΛO�!Tl�ĉ7y�r\�ɕ�0nC�:�<�]��ūN�!�}*��������)%���H���mB�HU��>s���J��[�u�Q�snm���G<?Z(��[���I$��|hd)L�r����\���[�ɜ6_
Evi��Vi�������w����Dc�o����2�#��������tT&t^�� Q����a�i=�Ɣ��ABμ@��S`7�8 �8�x��)r�Q��{.z,�]C�J���j$��_�n�JԞ����p�m�R����yÄ��2a<	J��
��G�PE��OL�	��J	��hj�]"����ߺyھE��SF�uӂ��I�;`)���i�~ߑ�/�y��>RI�`�(P�!�	ut�m��xIP�.�&�� �ۍSG�&:gW�
�%;���"j(��	T�]q\:9l��0n�-25����
�M[l���0]x�g��r{36��G�N������w�<��޹U쵒wD=�4˶m�%mM*�ܓ,�k��ٶc�)e`�<��b���1=毎`��Mэ6�|Ns^ u��Q	H|Op�B�9�s=�&�����`8�zx[
��G%�H|D��'�S��8y��-V(�r�'��婅�YQ���Z�Lu��
!�	��4"*�jӞ��,���8Y���W�L0-2��]��Vw������qeX�S΁.y`y;i�P�������*��)� �` )�9go)�yH9*_7�8L J�Zi�Ph�]����r��T�EC8�I�t��\6w�Z���g��ױdY	vsԴ����i&%���s���y��\ss�iv���E�b�n�Ȧ�Ա��p��7������T�0�gM���z�{��>�ddajA��,_��� �G�U���hHB������z�c�o��Y�6��ZM�ф��7Cy8��҇����'���,�n�(�H�g8p��t4�g����~g�j*\.���.J��I6�o��%7�5��ť�8����[�=,O	
1�D�!W���;f��}�[�x�W	���3������/}�8�=�w��R�vY����خpkiWi�'i�A(���c��9"���r�i&e�U�Vw�����+�lpy�z�l�!ґ3N�_�X�$���a#�d �����G�b��2��H)6��k��z�=��[��%�q���J�I��p���ML���N0���&����
�SPo h\��1A�����1��f�M���r}Xͱ���ņq��{	U󞇝 {,��V�66����@KF�L�n��(%N�L��?�{��or�ݏD�}(�'GA٦���ZLN���àUy&MuEl���9qZD��
"�Hv���s:Ge��Hw�I��(s;��\�Rq��%8{gg�նՍ��F$�X'V�?�<��=9�]%T4	�E+��K��gw�%��PFDX�ϓ��=�-q����=���n�8�~�_�P^0/�wgя\��ںEX��>">ف��� �33q�w�.B"��\�|Ѫ �.����E>M�P�6X�ZFM�7Lj7��yI�cwd�{�n��꛰ Tl���b֡=��;��\��{��޺U��B�O\h����9��.�[{ �C��.�;��ӝ�h �ێq�	�83�W1�7|��րS�B@�F���}��_�]+��8xHJ<�C�8�]��3+T��&i�#�3  {�bӺ�ez0G0��ek۝*�P�k�����kTwߦ홺�;�G:%��}��"E��bkV�m�3�m�xk)	$�c���{��q9B��H��`h���ҽG�II󊴖��sP_�z͗���r�\ᥘ��{���g[�vN��PR�GK����H�������#�����6��Lg.��ݑ3���X/����<�e�&Q԰h��3\���_$�#��@E�)�h@�Qx�P�}k��!y±,�%6�2��y�M�g�-�Tj��*����A���h��Ng�ȃ�5����Q��ǎ����V-g��)  F��%��2�X�SĚd/�z��q���Y/�Ɲˏ�zI?�mQ�Ƈ�?(%�9tN�;�:m�p��QEoY�?/ny�cOe^��ɉ�1fZ6�^�l�
ܷ�ZC�xEB$i��\�"�K��(%��va���ucSm�O�3�26���@Q�mXl�@35evFs���]��?5S�Ot3���m����z�@{M��ʳ�� ��y�u�)	l�B!��qsQs_���4۫F���PI;��Z�Uw��m�d��R�R������)�[��	{���8��׶z�O����`�FVWeG�)��c��g"��t$|K���9y&���+ڻ�h0|���*đ,|�U�A�՘�.��"c�����ba����9������7_�m��r��`�\�����r~�-`��۸ִ�����.Y#%�'�0�p@e���p�w'���,��SlK���q���X���� ���F��= ��ɧ�����y�	�k��)GGܳ�\$����n�v�!�lFo���^ߩ@vm�%LB�+�i���ڵ�����'�i�L[�W{ؾ��/�A-$%2F��2[�����9�!����1��L�)�C����s}U���m~Re���V�[�<y3�?P�>s��:!�E*԰�:�a;��V���jF�Qq��8�^�$k��ʳr��&;���gɘ�!��ME
��^f�h�&6poE�f7�VA���B��؇y�n�J��srx�h�ݜ��
�p�1;_�����Ӈ'B�u�yq�M�p6��n��1o3�����$ أWV���s?��@�dU�^LD���8�͜��ۈ&�56��\CL}e��=��4P��9�F}�0�+3�C�+��#����w=	�Mk���6`��&f8^�6wY���j��!Y�1\���`���/Q�� �e�$�8A%Bj�}���}��f�)Qv��γ���c���B�g6�@��p"���S�f��r�%׃6�9���ת��d/Pbb�[G����e����*�� �;���3T�"��8 �ҋ���y���z~{2]M�	����L;��>?C=
��*�y)v��>w 
��e��I��������rw�?�{ �%�Q�x���1��h����Iؙ��fh�[�S�?�Ø��D�׿���h���0����p��٤�ϋ�z���P�0>�E���db�IfsѾ�&�S�Պ�8T&�]3�6N�6�A;	��%�=ܯ�k�y��O���ll8Y�K������% �8�خ��>��?�}J�n"�`+F�������3���0�x�(ʔc��$�G)�Ӈ����+� q0��K��~���=M�nn��0.6�Otх	�w�!^���V�E͝��Dv�T_�]K����Ӈ��Pv�.wk3��qJc=hn�y��#KK2�a/�� ����u�����?"����M����/f�HXMd!L%%[�Zf�ȯ���;��`����Y\�� $��F[E�����BP����[�c�S`A������;s�����OUEy��ri3��͸ M��u��e�܏�8ɔ\���,o(w�.ͫ-�2�D����ܘ�4\���.�6�4=ꍊ]�z��@����	��[(�Zp��� ���h����R�9�(����S�v����W3�T�{6�9 ��+%v�4f��|J�j5���I�ȅ�Ѯ��x��.b43�/��C����<�=㢒̯捵��MQ���g�0, \t�#����&}�#�����f�ee�,(tڵRWb"�6�mX1�qe��y�"�AR�-�­I���=�R��r`6�����}��
kl~����[�!�[iMD�Q�f*�)� ����@�����X�mc�p^������Ć��Zb|���8��& 0��@�Am�:���Ua1RZ��T��w�o�}Z�3ݾ�>
<)?|%�B�K5�i{�T6�r����+��"��
�V��Ș�͵�O��H�t��$� M��%$�~�I.�њ�P!>D_�:\~�Zq�@;`Җ��Ϲ��D	[V���
�&A��Q�bՖUr:u�ZioM=�Tߖ;�]&Q�l>,��1��>��sǑX2C�9ߧ���3�Slh�#�9��X9Ě�̨���^1/�D�~�����l�����~���#@�-�+�m)w�W��Hq�8?��9���+\s��U�UTctL[ԮQ�~Q0m�a�}R2�8P����޺
��G�;�I��m�a�ï�{��KZnZ`3_lbq�U�:*�2�Y��A��U�%��0��-|�r�
2�*B�`.a~7�$2�^ڲ��:�S���t��hO^������� G�<��d���_�B0|8���7�=$]�6%H��'B4V����ߥ��z���cfyF�"�ݵ�[�}[I��N���C3F���Tb���,�Ƀ��JUE-�A�H[�����X1��7��Pg�<y����Y�!���ŷ����CXZ1G
���f���R�T�Ua�c4H߾q@ z,g�T��v�>hrĵ!ɷ�]u: NZ�'�Bh��e�g�����_���>c��S=�M!>/h�Y�tnǕ���Es�a���+��Y����XT�L���Ƿ�b2]�Amki�@б�g�c� ��%	5Om%�����	)\?��Qj�p�XF2<�T�:����w����?�[,��� ��ON����˶����u8Q�U��������֚>�('Vo��V����!�1�t4Qdu����W�,�%n�����kL�eE�6H�G1�Ā���Eltj���P��v5>���9P��q�
��L��3�aL�}H��ܭL=�DIA)*u}6��K��3����Z�ҥ[���ޛ9W��o�Љ���i�uٖ�Ş�u{:�`QSE*�̥���S%A���|��M��L;�>%��������Y�G���i�����ʗ�:o�u� ��+?ke�nc��)W��rK�K��K'����?$&�Iہo8��})$�� #_���Au�s=t7��b?L��Q3�� ��f�	�T\��v���K���:������pT�(Z�bx��oa��h�����Y��t;��/ܼ�<�Pz�Ȝ���Of�w0&�������%z��5��\���e+����."����٤�(0��C�+��ٿ���T�	ޅ�N*��V��^xR�ۏc��jiOpD��	#r�6�e؎��JT_�4h�Ah�)��+���7�k']/�=�4w,�Sh�.�
ybl<_oʨ�����Zk};�G^ɿ*>���k����z�VL��JD��|M���9�O��c2J�۪DD�q�<>7�48�G���~��P;��|�.{jz�5� H�	�g��@�Ŵ���ηS�Y����W���\~�0uK�p!r��������F-�4|(��e \�|����*��k�tC`��\���L�z�ה��c��{v�T�V-���B �w�|�{"�Ia�W%�S������DY8�c�����:d���y"��:~��b�� S���9y����nOO�L��������ӱ��$c��L@�{��?3�3��{w�;jeZ�
�m�︙��Hk�D���Np���5|�K,�|2��n�T�uA+D.l��K�������V�ϠR�F�۝;�7�$�䡄�����'�2C��^�[6�xI��U��'n��N�{&9ni ���i�{i�09��Be�<I�X��=)�xL� ���k�~|��������,i�pB�+�����HEO�)���SVDB�I��Z_L+8̰ӂMc�������"��W@������!���� NK>���yv�N�?���vW!G@�К�xsh��q3���0X�5�����|�+뎳���[���]v�'��Xd	K=s�����}{c��\�n��t׍KӄiL�rC�P���-�:�6̵�Dǣ�EWWI����k�2v�O�S�`��ܮF�h���ΰGB�,�s�Lfk�\��9�Lǚ'\��v6�~���9W���U�ge��dm�6t%ȶ =�з�;��m�7�8��?�Gۤ��A���~�AO�*�}��D�>z��#6x�����v-xoV�ʒ��H8��o�0{mD�+RJ���/Q��I�:אc������;!P�� ��m�~숹��]V���WaF�&a�^�����!�����=ſ�<lC�����"S�CI����1;f�q�Sȸ�v�L-zi�<>�/����feV�K������}d.4�&Ale0�Ht˖���)�?��� 7���!��t�E�^�`�3�:��S�?� �I��#�✩|^O��8w9q�b���#%p��V���9���A�t�D~�aS�Q���[��*gz��˭�/zzfYn����!P�=�зA�5��?w�@y�~s2BU�%{q	�;B8{� Зx|��o�&���Q�"���r�a��zr;*c������@��ܯ#G�Sc�ɱ����A1�}`�4�����Ѫ��\����~y�m9٭q<D/F|�����Սy4̷����]�>~^$�m�� ��h�
+8���G�H�K��%B�%�z6�����)D�{�@���?1���M?:^�Έ���6I؟�B
V5Uι�*g����n���5���u�f	�֋����j�v�Q��p)��l<Gl!lq�xH�I����w.�G��r���f���f�t�55-����)
0N� �e��R���yB�������02�b���H'�W�����c%����\�jA&�8�GcH�"먕 �̺c�euwv��� y�QK�^4CI��iV�cE���歘M� Nկ�eY1�5-3'��u;�0��5�hή6"y�۰H�Ơx �M�(�d�K[-d���$Z99�̘�%YZlp!a)�����?���f�,^ �\��-�f��l�d�^�޳���x���l<�k�m|��s�F�..K�H�tD�¸$Q+����:{Ǘ��2�(B�/G�&�y�Z=s��OEtWKh���Q�E��-�y�~
j bٱ(��`a=�5i�=G�į�c1�Q���jH��]�A��q��v������G�b!���-���en��?'bԼsA
��3v����9���V��q�M�'����l�Y�!8.��sx/��4�n�a�_*ӯ�!�w��7�4�=&w�G�Q�'4����l��\`ؙ D����Ǩ�?���5bj��"�����O�u�K��3UL�Ԏ>���=j��X~8c��d;_�����W˕�:8�]c��%PH2#��Jiy�� -�>;�|V�pcHʣ"5@�!ǯp̦v�OX�H�`�_��U�:C.`>�Io|��$���;"�u�Z<rʞ����ѫ !�%|�r�O#?���e�����w����l�(�Y���V����N�}J��V�J��%Hg+�b��G��6�d��	��M)�Qy��B�j�\"ӿ��I"p��<�e�+�瘺P@&���^%�Cժ�ό�?55#�]4K!Ԟ�:�rA���ut�@�G���,9��=IχB�����ȷ�CX�k�4�_?6���4Q�N�G�N�/�Wt�n[��s���D�s�����2Gf��-�n����5	�y������#�v�{^��v�_��&-u�
t:YzE�ɔ;��|��gk�w�ݎ�l,0����Ͷ�Z�ȍ�OG"`�R5Ʈ�E�ou��s��?�"k�-1G�t:���dt�V�.��+�v,�d*RqˤY�hl�t]	�Z�OB��.��k/��g�+�0Ϣr�	�TFk�fBP������Ohs��H��Yf�4�G�
�9���񅣀��ܵ<H)u���̩�3S�;b`K�a�C�0�4��7,�����>R�{� 5�d��#(_��'�_�D�`����u]��>	��ڛCe�� 0�reK���bP?�ʑ�iӊ���M������,���J�G�n��������+�*`1����㥟�oWZu��,}��J1������S�D6�GN����
禟l�����������M���K�X����bF-�F���AMA�g���Q�N��5�c8>q$0@�:��`
���|~	פ����U���gʖb��b;m'���=$��H k���b�4��:`�[E�q�*w(��fY�[ڻd��������1V
�l��8�u�9)�V�q �o��,,<��.kb��ۅ`��Ӿ@bAR:?�R�(Ϧ��D=.=���6k m���P�tuNJx���V����s���!�Ś���t��4>��z�n���f�e�U��%v8l��4h����6KX�o}q���6�2�=lZ㗞%G(�~�Ǟ�=@�*��jWŎ���j��L%1�kzK���y7D"�|��2a�@iްP�jb��Qֻ����l�uS��m֯vS����>3ib�Ǫ!���l�E���Q�N����Ϭ}�5=�Nmco!��)������ea����J�v{�C�TL���Q�+e 9�m����N���s������j���FƌV�[����;�5<Gs�멳x-t�l�t����I�x���:=Z�F����VY �C0;s�y�o"�u� (�QF�޲78g�8���tV�]��} E
wr���`��Yss��a��e�k�~�a����`uw�T�k�8��6�'ܑ�doָ����і���2Չ��na $��ܭ(�U�C(mn�S����-Of�AM�Oҟ����\h%v�˙yў�����7�fwᭌY����..��wT�<9�C��M�]���X̚�r���4��c�ې��IU37L�x���X_FK�F����\������Lو�R_?:�2���Q,1�D���q� ��$��!@K[�P�4M8�W��6�7�&Dʪ��}�y�f\�<5l��(A�2�ܶ�8���ڷ\*)[N���̖̘11��c ̞��%+py�?���aū�)��E%���NgZ�?l�34�,cNb�1�2 ���b��Zɢuw�Ǧ8A�U�[�j�
��\�w`����f�\�&����,}>��ւ?E���QJ�C&��?�
���jN3X�͙Y[���BU�4��MN�����%*�_hq�"��U��*9�Q}�6 :K�-��>$n��H^8t��Q����[.��v�/���E�*�q�a�����X�`z�6ք��
6:�ס�~�]I΋�m�0�D�᥍&��I}?� s�y�wlp8MK�䲏���j�>h��u��R&���G����֐�~���i��]Oe�q}��2u�������%`�3tg�No�{E�&��&��V�3 ��Jh��o��"��2��N�8^>a��K�!��U�d�Za�^�Ԥ��s�O3;+�vQtLz"b�����SKD�ЁE�ISWTf0�/`���a1�I'beJ	Aj����p��bryi`�S�9�; dˇB+,�Z1�+w��O:��>�d�ʇ�x�x$1[��Nr	^�28ʚ��)V���J��w���K�0��@��{2[T� "�A�c(^�>�H�����<{?�z�!*�A�$q�Ӈ�I���1�g��!`%��1n�f��J6#~b��,�`��歲=�oY[��g���n��y,�#i��,�zު�����Z�vwd׾�"n��dlQ>*���HG$k�����T"��a�(����|�t�HiI�'X@��ə�(��$�bЉ|xUd��/7/�x�=F����H���P$��_�g�N�{�6#�FoF��p����B,X��"����ͅ�ӭ'�b$'�����3�*�Li��eq��r�,��A�z�o��^]�@Ej"O�1{�_P�~�ն���V�Rv?ܰx�"/<�U5���pE�O}�i�$cE���V��ꨉ�H���z�w􉄎�I^�X�!N'����4A���n+챦Nv���?J���<AF �6,�s*�g�y�5�wP��
��v�`A�K;RQ���)���?��2h�����טW�A���U��s���Mժ�YZ���ka�d�%-�)��[2�W�NL�j��?R4\|�>h��Y\�����4L���pZ�NO�_��O-/�K@����aƎ�q�tJ�?���8B��vy�����-����o'?"3�vt�<��N�e��?�ѣ�M��ڄ`b���K{ICTB׌�]��O���� �6���y����;��@�om��,}.<��c�i�~	�)�g�ǔ�̎�ǃ���4��%���I#D8�XÂjT�n>#�b��g<IVe�1�~��䚌VR0.�j[�L��4Z$ޜ�?�(�Ojg�p[�QAsw��+Q����s��ErIG�J08�j�E���r �ܻb���z𪟐w�}�j�d��6��1��3͚QXK|4�&"%��{���8��φV�g����T���	m̐S�C��x�
,2��)�%\#x����"k�
����ftAj��_��p�0@z=�V��_4l6��&��@&|F��\"�mh��[E)�d	�O�M@�9c��������`Ldɐ��d�Hd[�3)Z��Y�>�Ps�Eh`֥D�P��=�ŉ����o��F�Р��ǰ'�.:+��ரJ8pc�AE%��2��EQW��&��H��Xj�/i�ҷ�IJ�M��
BZl�55�M�������t2�J������z�^���	��I��HK%Ӹn-F���$-�ٹ���L*�5�<�"PE�(��:�9�}�"����:~����X˜BtJW ,�'�f�׎��	S�c�~���M�5�
*)orf+�%?o��N\b� >�w��NP�ꦥ�m�Թ�s*1��ЋA���gf[ w4��8/ap�S9�G���ڔ�@tA�	�atS驁��Q��}�M �F��`w�&�U{��� �����D�õ���1�*p�%i��^O+F#qj	��#j|�X�Ik(iM^?S�l���ެ�07��O�\9(����T+�Qx�D�.��8��y������D%)G���;Q�U��'e�1�_x���p�bq���p#h�"M4���W�ٵ����C��Rڸ����S�nx�wd	a)��Ό����K)�1�y�{snI��`�sʇI��}�vtm��ЫG^��3,�2=���S��xy�:{Χ��'�~��7⩵���߁��y���ᕜ�E��V�9�DM��+��LqW�ӳ���$٧���y\W�Ae�|�����{���B!�j��\b����u<;V�~�,~$K,�=&���F�>jF��fǲ�n��2����Sف��,�Q�����z����`�.k�U�^*���u �^ҝ��>������?$��=0��M���N�|pW����)��p��]��C����v�&���ʹj�
��G�x���1$��r���KKڔ_�Z|��)�xS�C��F�(\Ntu�XA�g#�I��#�
1�+��R-	���ru����<�Z.�q7f�6���b#)}�^���=�`J_v��k�}i�~�3����S9/�ŀ^ Vɍ|:.j Yp3�_�4�!���/W��OTe���݌� �u�#��y����3��T`@l�Y�s�>�Bw}H�߷h� c�6 �u�m"��t��#��Ń5��1 �k͵����^�3����ˊ�`�Dbc��J�>[&��Zq�0K��L���y�QC��=^�8�{��X���s��
��p�$XƷ�A�������e�!N����>�'�f���5�4�PY<����i��k&�V��HP)+�Ԕ~��P�9Ҟ@D�9̔���)@�ք�6 ���@)B�d�wS�q�c_��A1��È�k,��k�t7�	��!�������ڪ�?9�-�	���+�����C��"n� ��O���9��t� �`&�/���j�&��W��=�Cq@�n���/���8j�����-����
�\�М���
̸I�;�c�v�K��_�w8���o�1U�,�-�Q��U���#0k�|6"2܆�|}�k0w���*��c�̻��3�����ofߤZ8��4�<����� VK;��қ���/�X�|&�gq��|��=+&��T��w[�wҘ��b�n����^br4Ў�m,dQ^�������i.ο����	�<�K�E�*�� ����LH	��(G##�,�9%R^��!^T5}R�� �w����<���vI�wa~J��>��:��-�*nF����@���)�+�u��ut����q�_�����z�j�h�
�R�,�>פ�ҍŹ��V �D�������0�_k��fʜ7A�A$TDe��-�1&n;�c�/�aC>)��	���=�����.�t���x����\|��q�m�#0'8񔛷,J7 ��_�O��	b���y�#'+Sd���|L )��Ǥ�+�̗���	�D\�[z<s�pk�$p7��1Q�.L�䐊�+�Hn^�{�j-�j`�uK)î%W�WX봁���5�?�#��{����\R���^f?T��5�.�6��:��9�R��υ�e�u�z��o%ߪ`G#�.�!�����I��0anj(E)Z�����fb���=�P�����9޽���h�N��LM��vgV�J�+�`�����$B�C7r����Q׾�aT&��3���ef����/�D��Ge�U�B7������߇x�Ƭ���ܷI:���[���{�U
�h�?WP铨�1�5���{��Y��#��[��#o���OYg���W񋑄��FBa��w�m�@H^�C,:i��2%X:��l�����	���58������gv_��7��W�+��q�fi��+�@�����`5�UZ�,�����V��å�NF�dvMX[-�L+�u6kN@���>\;���Z�{��Ha�J���aǺ�E�3`�U,E�r��ux����Q���՘M�D�2T��&Xo o�ID�B@��6�nK�D5�s�(�QվT
�J��x(��XO񷺢��,��b^�Т�p(��S��;����^�e��3m�Ɩ�<� �U�d,�S9��LhaRA���2U�WVs{��*k��M۸������!�/L��L��e��[?E�ut��k�2��W��������<-��1q���f����?�=d����c�kу�=��
��Ka	������HkrQ]�<�nu�F]B|͔@uɬŉ��͓�KX�6�3o��ٗ��w�7���ڝ�X����gY�"]55�����n���E�c��n���K��#�����M��������k2�#3.59��b�H�-[����ݔ��]�Б6 ��6��h]0�Gm�j)CPXx�����񛊯�h<�x���M}_��)B)�F�`
q۰����֊Zg���1���ցl���#/Y���(6�L̯�;Y���>WwY�T��f�2�g�Aj�/4<zk���[��Ab�M�L���K��e��� ���rOP:�ꠔ3-���	�X�Mv�1C@�l&�k	�c޹����ý'���ڐV����m	sJ�Y+>��ȇUg�^��Z(_̅n��g�`nܭ�m���J�~1�ߖ��آ�T~N�P�X� S+��G9b�ޝ��LYV��9,�{��T�5lwJ�q=��6����J�),UA�����v���P������0�h����ׄ��fK��>n.׼7'�N�F��,��PKp�y����;��Ո� *n|k�X�YmV�ۗ�#�u.;&$u?�-�c�潚��~��O�.�8h���ly�M��ɒ�nj.��;5��Y}�1n*a�N8>̼0������r�iP2�62}:*���ʊkI���񽚷�����^E��q͆*EO�E�T{�=uQB�y9�6�6�,T���lE$���}G���^�% ���}�	���0�MD��wq0�t�mw�f[C�S0�U�I�M�v�\�D��8�@��v�>D���W�<(��W���Ba�%�� ��B+ٶ@9o���9,�}�{yK�k�g̙��@_㼠��Շ_��#�M�%8��kQ�m�N){\���R���R�@�UV7\��4	�2,ޒ�>[o]���1Ӟ�.9���&?FI�KU��Y_+;�Y���|i4��}P�Ȉ�.�fw��u���h�L�G<�����A�wP}�T�l!��6\�E����'�xԇ�������i���S�[�>곾�k�-�GZ!�D��u�����=�Wٺ @��2&��*gxh�s��Yk���� &��GS�&]K�B3��k~t����A�Ze�Q��,���o��C�f�����6r���~e�)������J�'�Wi�3Qm�����2ѐ�� ̌(.�^��*��#����0+����;�F����-K���i!�s	��{q

B*'(v?�_~���`�X�ԣ�9��&�Q���Cr	`��9R��Ք�J�R�Rf��di�����?	���~���3�	� ��ƛY��ڽ�v����n�20[FMi��D����6�}�eJRk z\��(+����7}�'W���]���q[�/�_{����+xT���_�0f��Z�^�/"2ج��M�ܜF7����d�> ��}~�\��:�p��:?���Bӂj��B�o��s��$�C��%���L�9�l�-	W4�����1t�!��p��U��v� :e@cD����+a��������R�4��^�L�������/�����*R�):���)Nj��z��8�/:�nO@�( 4|Ш~�!�6���ʺ;Y���%�����ut�X��}�:f#i �F�U�[},� ��9���֎ϯ�xEd9W����E��Pr��C��ˏ��5��|v��am�,5(c��*&w��,)"J�ۼŤCH�R��u��;��&���"���M ��+�*'��1�������k~+ w]�S\Q��0�2)����ǻ�p�w|,Ō��*�\U�q�m��	�����\��9�Z����Iu�n��`���u�ԭSXB>dv��ib��[��j&^�EӘ�,��2q�wk��p	�WxSL���,m��� >N9vk�H��m3���Y�(⇘��8_��	���#VO�{!�O{mW6�b��ž��p���q�X��e�x���N�<*��ݙ��z���K��揸u>ȴ��sXB��~vx�wb�ַd���PT~�\z�s4�Pnቇ��W��f���(Y)�J,b��L>���|l�d(!Ɨp��ѡM�@��F��2��c�O0a �4��5��O<�O�=c�B�"�t��O��9�H�~���#������q֨����3Kl5���|C���Q�v��j$�7�B�,զil�8�I|n�}m�\��I�B�����Oy��gɆ�8������c[���Ѵ��'�9&����-���/��.=��
O����8J̐$���)fD�y X��x4b��+@1�&���>��V-����>߶I�Gy.Ai�q_�����1��ݱSC ��~���Ƌ���
�ղ���'Xft�Q8��Oao��~/6-����5᤭Y2����[Qލ�P4/�@M�:��c?x#��!)2���W/,���&��A�ɰ��u��0����L��2�0���T,�h������q=S���)�"�~k�L3�?jѫk�=ǸX7%|{�?�п���"j��|�e��\�yH�����$7k�2� M�={xU$F�>�Hv�S�=��{MK�,q�b��m2���A>��%���׊v��v#�4�PS��q�΀$�w&�L��1�X�R�C��$FQ��E��s㗩��?K��A]_�4-�CѲm�A25F����-�DU�ݒPd�羂K�ɅgJ=�e��t _Q�+�^ �鴏��#yڑ��T���ځ���J��I�D�%q皠��_0��6�,-���;U����8�4��e�h>��ǯ:��L���/	��Ⱦ�ӠW����jy(�
S�K�{$/��G�5<���+�Ew�ļ\����2���]_�1w�C��C))mq�<l�{��^P�5y��r�1;���L7��;Z8={r׽�C~�M*9�'rt�p�߫AY�6�����)C���Rt ��ݱ�^��~Z++ 
�Q�j���;����IA�@h.�#R�4�������/Ckd�du����V����c��7�d��N�g�ó��kW���|�FQDҡ�6BC%�	5@)	?�B��a7�c�z��@�}u��5W����X>q~��r]r�T>��R45ϗ<�"t��`$?��1˥g>�N�.�&�q%e�?܊D@� �"��<�p7����2����j�����x�y�I��bf3f�7]u�va����t{r&4�=Y���C�6��a�AP�b�>X�V\�g7�����j[w)�=0u�*��-��ӌ�����+ GlP�Fg�{�0"\�=�b0��Z�u������=3}�YR�&�-�Y��dπ\�/��s<�H����a�����h�P@2��Bב>q�%K{�?�h�A?�6��p��/�
Ȇ�I�u?g��d,=��	#G#/A�ׅ��e�*�����#�9-�s&?�e���H<�b��3���E�=�Nv��+��%<�?d�l�}1�a�o� �q�(0K��X�qg�>�l�%q���jo�A:�/�`u���@
��v�Y�/��&Us�0_n�}��W��o-<S?�M���(��	���K[sj3{_ˣ���L\Z[3��W�?�σ�� ������e�G�c�	�3d�G�-��hn��9��G���jfQQ�K������e���ScY)��a�.�̔kG8�2�w`]����P�_	DО��l;{J��n>��]|��Q�[�3X�*X	~��+�3&��}b7c�ț߉�����*�ԕн8͝
|)Z����׭ΚZ`����߶�F�����i�Rl��fY�-[��n����æ��{\sN%理Ϲf�Y�xw7)�vXL-���\������4n�|Z���H�X�oM{j/.�Y��;+�Ig����]�y`��x--�[k	��Lf�4ú�M ?RU���4`�0��)���I����P2l���R���<����0���S�!��p�p�p"<@����IU�Z�+@oU�G&�${C��l��"n��Ze|O��)�u��`E���Wp*��?VFK��}�`x�.��?�!<������U�09����ͮ�&$V����&\���C���&\�T�>S۔��j-�;���\q�rF�gU��ͽ朣 ��6%��qm�C�.� [�	f�W�R l�3����\QG��
=7��$;���+���w>�=��^�&�A$�P�����k�_��qJrS7@<��5P��p�xfi�9A�t`C�����t���E���%���__"�Ie�E��Ž�T(i_]vdQ,��R��y�M4��GRv<S9��1�B��o�">�'K{]V�x�v0�k�v �H�>ThK��� �;K���^���M��!Mr�cơ	TQ��L���J%b��CB�o��q��?x��4a�Вm�4C�����;/��P��en������b��^!�e�fz�lˤlT������h��QMw�LȔ�zgX<"�G�Yj��hI��Jҡ;��r� ��.ޖ��"�~@\�'L����3�~�HG�J��	��.��%{���.TVG�]�Zi�di�[G�1q��T�Vq�?���
�|�[yn*�ʷ���!��n���݊�.2e�V(}R�c�ӓ�=O���B� ����V,*}�O8H�f�@v��Ӆm8��V��u�vt]ʀ��j���o���&��q"�wǻ���i½��	�֔X�ӟ��)X��٭n�[�
�2����px+T1+�"��q��D��]R�Zl��Go�ޓ+ktS�)voy<ڙ�i��)M߸�ռ���X�����j��}�������O�^	.��T*^ פ�@�a���0$�t��6&S�B��D���Nk^r��k$_$������&ݜq�����瀧�8P�e��geх���>��&�����-�3���d2��Y��`�[�	�>G�h�y�,-Sl�3���8�ǷR)_�?:I9,F�UIVJ�N��Xq5�b�Z�R���T?=	��=i�^�e�0?Ù�~�_��G�D��7|Z lw�_^�w����+���6{�#B�H:3@��|N�VM�`�(��d���T��P<��8�a�W���%����á~����!���Y��̸��	��� @Q��5�L�c!��[����Fؒ������ɽ���$h!��kL��h�y�	��M��c|r�9���H��C�c�4S�k�
Bް��(��|�*�j-�6K:�r��_ˑ�U
˘YuCS��|�������_xLI�+'�4S�˄�Pf�Z#yt��7@1�|�na�N�.��4^�'U�tV�a۪o���6�����O[�}Ć9���?6$K����SN�;<�(X|�(�N���z `�'6�
}#��Y&��	�Vn5�ѭ�'o���|Q�MM�n��2�/AY�ɒ�H��@r�
��RRE�}�&8A x%Zc[4���&��3�4,�l7�R�vP%����4)���s"6A�!���?��0}J�X3МMͼ����=�i�w\OG��ClCH���uF~��HilYL̢~������D�6��d�5-.��\�����C�j���F�P��"+4���PJ+'@ �/�~0u��ݜ,�щ̚�`kX�Ss�%*�[@e#��}"M��\�+��A�����F��3�h����}SLV�N�s5T�Q��i{J�^.N� |����co��P�C����5r�>$�����Q��:9�Kj�u�|zƽ�릣��2x�~z�nQ�B�,�W"��G��I��g,RΦ� �營t]�>G:<���M+)+�|:�sf`=Jc8��d#��'�U��U3���q�w����rA�������Nq��r=ҍ�&UL�;���q�=�&�e��g�:!ZS �`��t�K���d����o�5��7_W�75�������/�6E��Z4 ɬd�.�
����1�����Ht.B�%�%OV�I^F���"J�~ĉf�"�N*�mA6(��\�IHIe#?U<|�T��T�D�QKER*�������S(J�4Xp��8XJ|��Xj��~��g�T<�1Z�Tsl��=�c8�vu��r�U����B���@�q��Rǐ���vѮ����u1ف)5X�S��K�@/��Z�Ub�0L�}��s��D�~U/I:���=�p֪��leڊ�w��D��в^��X�9M��ɨF�xF���	~�o�T��y�"ԛ���D�p�ח9N��m�e~x�up	8l�4gۿ��	���,:HW����慫�GÐ�Ju����K�dF�N�T�,��B_�� A�A�4�ǚ×z�8H�-��j�>�}8��[j Lo&���s�B_����ؼ���}7cF�@��ё�|4Ċ8yq;���k ��?�nI�L�y#���}���o�E�|�M���p�c�lŻ�Y��B�H�YG�3�7�Ҋ���Y��������(��m7�v>1�U	w܀L�`������ 4�c�Ci}Y�Y���Ԁu��t�����##
q�-A�"N��"�b�@�8Qw��KM���4�u)G����*T�����0?����R�9b_�s�?NC:�a���:�r�I�T�ʩ�.�{'����:�w1��yĽ�D���o-�b1�D|����LA-\�9�A�C�9�/Eބ��W��W!�\iyA�/ϙk�$>�stQPPv������/�s $?z����T������@��v� n�Lw�7��
A�B��*3�9���я
�5�����@XMA'��Q]j���M 7�e=I��UY`��m>	}vv�����2�ia.��=��0�K$QZ"Jy���ُ�(;�K��h�2yߩ��N�1�{���.���6<@���U4��ֲ��\�K�২T�s"&l�;k��V��xDM���S��*)鉩 f^�J��_c�\����B�TT��/TL@:��S�����+��*�_�J�
�&U����&8��`�Y�mĳ��� sg��YY���3�����ё]� ~y�_.�RF{B�s�s�˃��@��.��;��Ӥ`�4=��p_��*�վ��=�G&�F�����Kk�������횴�=Z���	X9���^쀐�x���B�cߥ���o�`���r0#�/�2'��gle
*��Ee1h�����ɓ�v�*:�!�1��5~�EP�Q\�O�=��y�ެ�kW��բ_]A�A(E�����h62�%��c����ceˢ)F�(�D�`�Dg&��h��wb>��边d?��ig��'Z�V�FfK���vc0#s�������P�,/񹜨�^CQm*�k搒�ˉ�n��L}%�E�����`��ֳES���#E�F��BZTj����2�k��@���0N��t��Y�uJ{s�ߏl56��l+�Uh��O�"C�Ψ;��u�?������W�h��Jx ($K�\c�F��T
�Ľ��l������R�;��Oe��dY��C�9#�h����cNO��F�ʾm%Y4�Ww���v�;�L�S���Τ�Zn2���?"��y1^Ύ�BV�&��MB�=�5�R��[�Z�a�� c��,-�A��ڒ���N=C���&2�������1-�ֈ�w�{�vN�J	[|÷���5����UK^6.7�Nb�^�߁E��F��㔭�!����$G;�d��`�pٹ��#̃�-����w�*퐓��ky�9i�xֶ��Q꾵��;���x�YA����	��������*�ܢ��}���4��'@���Y��e;���F��7�A+.0r�]���zj/�R8�d�c���{�/0��+QUL�)�ǲ��^�sm(��Hq�6�ñ/m̰��JX]�ñ�L�>X�F��~?l�(s�|�vV��=�mV��w0��A��Ց33 q�'e��Zt�p�/T�@�����)��q�'��.�~�I1���a�#��;|����(�Z��kGG��YU�]V14&�s����A��L���L>W�\QfÀ�D����EXث����io��ae���v���Q/��ϑ�j�;z�J�u�U藟��f" Ӿ�h.2I��*"�XJ[�/U�Uf�>���្ǳ��4��<5�l�r6PH[�}���L�
S4�8��{�"5��d�-[��O>oc��J2>��ت	�J��qqQ��㔖r�Q1�N5��X�ʂS��6�P=�K-�x�]�53U�^z����PM��?��c�����WP,6�3\��Kx���k����r����yr���IǍ��Sak�������+�	�M�=��@�]#۩ ��ċ�ս���?�ӳ�S�����^޵�F�7�[���Ii�_�����Z�߯厉q�\MA֫��yw0��1i^��|c�`�J�(P�W;��G�/;����^M�_])�O��J��
^K�%%��TJ>�Y>�L��`��a8��_4|��߰����/��t�Q���������|�>��I�ot@੽�M2��> ۱ame<�����MÍ�/>�n�]$g4^e��a����%<���27u��N��>h�ܑR�uc�B��P2N���+�cc�&n�%�35���rn�䜞���j��+�-����L�yв��9uk3�Vf��t� JJ౟����*��KH=<	�Ʃ�7����L��8+�׃j��&�a��X74B2s�MD�	/W(����e��#Ҿ"I_��bgA˂��s��uX�X@:f�[@U�e�"9i�@k��>���S}����A��6����v��5҉ð�KƏ�뵏��|sUx�X��J�\�KN[�M�n�:��A`d���l2 T�<�V���-�c��ܧ�\�?P*��|�%`V��W��n����V�����W�hs�9�����xc�ܢ;܎�	�B����U����В:(�]֙�Y�����z�פG����<�*�UR���T�^��1��-b�.�h[�}$d�ݯia������h�1�(	�ҍ����u_S��g��n�BDOR
P��{��+�&f�9sڿE���y����܎�=Pf��@=�e^-���͑�
��6����ڃ�q��	2q"YL6��QT�\X�w,�v{���N���v|^ڲ>���?���b`�_��\P�r������)`0p��ݡ�@S��K���0�îo�pvR�"���0����ZI�WHo��{���;�ltE(Ic*2��۷�`���_:�R�~�������Y���/�gL�8��(x�	��k<zE�xK0p�E(SV�n[>�ܐπW�QN{�ք�~�:�-}��KW�y�!o���M�-�U�| ����Y�:�Si�c�Q������Z8�d���lBn������1<F��{򷖈v���A��t1�����֛Be����1�伴.ֽ`N�]��P���r�W��[@�r�5ܬ��%S�!W�-V���VB�:e��]"US��x�A%�j����UEPaG]u	�������mJ��C��D���:?��YW��B���r��n���Ի&���Ò�SQ��8@��$3���X������5�;����2=Be��p��w�� R��}�xn�j�4��Rm�Ba��5)Sw���C�9p˪>����+j�Ê�k�o��Z�Ac
�Do��-��
���3��f����c�k����n��^o�=�Nf6�J�$�RDo8]���0�J5	��c���q��W"<��_(*bD1d=�3�0п��]/��=en����@��}z�M�g�:��O@`N�s^�~ߑˉb�%z5��_��I��+򂬩���y����멆Z/��ٜF�eࡊw�C��4e�6]�����V���v�0����	c��2����C�V��є؆WL&̸U��5�iF�?�T�%/�[:�h�{����kW��|�#.5~>��Y���R)л6��ޥ�>x@�� �f�#�	xW��e­�=ׁ��M�7����X�6sr�G�&�Q׊8�ls�^��
>u�Hs�a�����@��n��)��t-��N��%����l�&�y:�.���4M�i��FJ2�1�i�\��8�W5���bq�D�Rg��[���u&�n�~�xK����>�����*'W��L�����cJ�^��h���K�Ū�<,�����sw[�f�j}�S�Hg��m�s����!m����������oyu^~`Z��{:㖤_^.�ɨO�"��p�<������ج}3cMC�5fk����s�yB�qD�%�ѿ�tpϖ���I�����+j�@��>�]��x�}#�b�~R#,�I���Ic��k��m�:e�s_�*����f����ԙ)o�
��&odUN{B\W�	�G �D	����bIT�r��jDj:�L}p}�Ȣ/Z�9	��;���	�J�:���pS)<>eƼ��O	�[�r���e��)S�λ��y�A��0�t[�3�D��¹^��r�?4�bU�x�{uȚ9;��P�R��n�'�c�����CQۃ���u�xz�p/�.ބC����@J�Z��� ��-³�T�� �E [屢3�gp$����<Һʌ�.Cƿ��Q�]��n�L���T4K}�}\_��E��|�j���놶����e^:��Aʶ�N��@R���o��P�%��O{�>�\jї�T��y���<�c'��?�[t,Bt�4���uL�O|��T�����B�k8��!}" GC⥱�̾᪼�fQJ�����F�ӂ��r/���9h+�!c2&.խ��J��Jf5m�6��v�� R�IW`^Aȴ�����Z�;����|�C���*z&|9U�;w���ЗA6�f�h�]Ԃ�W0`3@M̮�^NBޒ{�B�N�2��~6�_/��*u9�M^��jE���č���(rN�yIAe���:���d��.tg�{��K8_U�'�t:���f�8���)���=u�31���`AY��d!�<b����ć&�/�ԑ�l�d���tO�w�MR9ǧ�Fz�n&�fE"�/�Up�42�e�#TS"��{�5�J;>Ra�?�B��$Lo�;���h�w�b��2B`]�&Q�CX:�v��bO2lE��=�p%佈YPh�_�A 
�a����ڒLm�i��C��öMb�^�NP��bRN�Cv�����>���a�n��'��Ȏ�Y���qi7c���v(vN��Z@\V��6�����U��+���g����1!��U�oQ7���|�����e�y31��XG��{jt-8�AŅ�K`�G~Ϩcě[����$�QNa�GS�t���y{�K­Cmf���h !-���1ң� ?cL%���G�+����,sB���r��*OYWpZ��ܙ\8�>��w[���:1������`1�1-�K�h�ܽL�ԯW�~��y���^���{Zk��.�n�:��ir��"����:���q94�nb����P0WlH�n���a���x!�ajdC���[�9�QS[���� �-I0o�" �SU ���>J��w�����a�̥,�z"�zK<�x@��#���
�Y�A�:�n���20�!�؟�I�����-��vWړ,*q��3�+�/��&o��gR2�W��P�x3ڡ��F�2)�!��TcJ�)'��N��	�vad\�����;���'O���K�^0����-���(��m��.�H��_E��$���(�l�R�!c�R͡>ur�W��X3F)Ž�z���J"�?�a6}9�N���,~/�	�c#��gJu��I8�7���#�ID��v�����^v5�TU)U�j{|��7���������Zɾ�c����T%j"h���rK>��+ǎ%8�Gp�����_���wA��2э����Akg6}�=�K�f%�y~6�_o���>�D�z�r�	Z:�0i��!qv�F�<i��P}��|̀��ul��h�6Qk�a;@�BCњ�`��2fEv͔9�+�ʤm9�9k�-ns��K��kTx��+�]��H;��٪����N,�Yʨ^cqw��wѱ,��Dw���m��ۜ���ؙ+^�t��p�ȯ�'�t��7��O!�4�|��s{*�P�=���\z��I�ϊ�ʚ�Z���M�Y����4�ۇ�F��@s��"E�vY�UHQwp7NeoQpb�ʴ1��w�"����/�t4�д��QHT�{ ]y��n׮�l�r�E��!����j֣� ;8w��e�dᛝ�M}M�Q&�ҷ�-��?mز��������Gy����O:���.#�]ߔ�S/J�̷�����n�y���I�.��F�%�"�hRV]Ln�����e!�0���x�c�+�x*�	1�y��`���
Y�Q�{����U�'�}��G���#�(<�>�i;�iiZ|=-�������8,�E!���Ij�z��75�������Z,�?=�������]�RJ��wk�(JS{�o���v
߼rj�h?$JZ����gA�Z��tӮg�4�����X�ײ�N�a����@����/����������/J�������3�7^­Ը�		@@�.�2�W�;r]�|�1C�٢(!��a��X��"f+o?�z"��-*���_���F�w�97&WA=�1;���m�C�S�'C�?C�o�L��?�<͋م�<����G>������
5�\z8����P-�g��j���cM��F쎒s�/�(I�M6�x8=���M�AL���[��u�ײ���΋7�����A��М�n��YIa�o��\w���M���I1�h��c��|�q�ָ'�w�T7,���&ͮ�h��P�ɦ�
��'=�3�j,�E��L��C/�J��F���������ܭ�髌(s3�B�; �qH��H��&���B�YF�.�9��Kw��
6tx��Ë��bK���_5�-Y�Y:�`�[lY�����2��8_|����S\��;@���u�?ܘ%p����ExE�f��R/�g3���c]k�LJ�P �	M!��c�B�!� _8T:'�y��%�%��W:�T~B\��V"Uoq���r��S\�I�Dz3�j��#��u(Dj����= 1�-)���iL�>9حl
�w�h�����~qs����SD�,���54�,�}���{1C�1;��.�2��]4P���V'�T���xG:E�9b��
�m�k�R,�~� 3�*��J���i�j ����"z~Qp�L�D�u��6B����[je!�͘Se�Y�H"_`Vl���D�=��Jb��i;$AB�����������qʒ��4�����ߥc��s_�:�j�L�W({7��`��Lkv#b��M(�&�(3�|���q���WЏ�k�z�)�prvF�mQb��e�16��7���㷼T���m$�S~De�29��d�^�&�\��w�.b�h������:뻆�VEMg�F�י�w�m}�K�Qr�Q�����C��A�$遷�1�R�m
v��q{$;m�P@ݖ�X�Q���v�-!���{$!M�܈Opq��2X�Y|v��RW"�ζ� �z#~ȣ������hV���%���OМ��Ջ���<6�8�������%PC��b(��LIisy2<^N��/*62��L�ĝ)[t�@)B���}��LM�\	�¹�"�DA�|pxA��i�2Syٟ����¨�$�W�i�s>>�Z�M�AC��nW4�2@SL0��b% p1q���'�y�1]$�>��q�C�k�u��M��r���^HJ|�s���\U�Z<]�~P��R��C����
/;����B��: �_ ;s^��D���\������2暹�����A ,:vw$"�?#�-�y���8A4�M��Ka����׍ՠ�Zs�7�z 
�Y��� �Q�7E�)&0čg�<|��c�����;�d��ֺ��p�yf)D�w6 A�Ueno:���{¦=V@�p�����V��ō��{�Œg��,h�0V�<,��ڬ������u�o n�ؕmz���`Gf1�#t%����@eTi�}�'�[j�����bU���m�F��!��Gtι�s"��<��s�9..��8$}'p8�1��j"��7�9C´	p]�M���&��Za5��45(�j'�
�M�i�Htx���XIw��v��!�ݻa�*����I�elIg���r�}��
�Ċ{.��|�>�΀�����_��ðg<趧�t���4���@�v��Id(��{�dP���|c��]��y�kV�Տ��D(�8D��gB��W�D�9*"�2c�.�A�AC^�M�~r��jD�d�#�����XS�R��ӎ�w��	�'�6���q?k�J�F�VG�%HWd�fY �"�J�"�5�P�p�)�V�Z�0���ؚ��^+�hoo+���#X�,����L�j�&���_��0�ɫ렺��Ub��C�Q�m;���s�`+q,5<V5���e&���~�IRHƵ��\�/� �<��VZ��,=pXk=�%P�c��*U����c�e�"�R�0|Ls��ğx_�q�����YM��F"�4�1�P��5T�3���?
���b���O��A�E��O
ܶoX�3�e��굦2����Rm]'�Έ��91��}��dܥ��OɊ{pyF� �	�+�	�T�^]�岓t�*:�s���z.t�%���xRwD
���/����I�h���|[a(��|Ar���c�?��ZPj$��hdP|v_X��) ��o��Gj?8?#�=�C8��]���̢	�Ak��m�i���h�`��aR)�c��{f�K���˵����Y��l1�7�9�SO7��D��r*pȧ��~E8JA$�5Pz}g�V��c��jU�O*Q&0`O��ٷE��[�ġ��/aA�@������*�A����c��g�H�fWoNЮ%�AZ��<L�
B�'R�ƅ2(�F�9"�.�ժ>�9L���Y���3Ġ���g"=����ޟ��,���q�+�KTkmhKBN��şw�����%|(�4��<C4��J��>��	T\��*ή
�ϦE�e�7��a)�s�,m���X�f�^�M�J���݈�5�EOj��a��Yӻ�V/�,����������&��z�YG�$0�U�ܻG����872�R�{2�A�A�]]�1r˸���|�i�#���o��&�85�=��F�@�@ѭ�;3�P�s��Ƙ-Q?(�cK������"פ�����[�f���������h�δ�k��J&���g�9���v� d_
d�E�l�r�}�1Y��Bv�	��!&`�
>�yz�du7�����������d��wH�f����b� ����s�R��k H��Z����8�(%M�����t��;��v��I��5�bx�X�����*�
5*6!)᱔j�LC2���&=�$�M�،2��L�b]��<�0���,�c!�ڢ���#JW����|����xyt��}����ۨ��v)Z�$��=�J�x˾E��`�A���z�X˾�])7��l��YH��_��T�ycѴ
��O�����^)Zx�	�7����˔�	��,��b$g�L�*�^CJ��m��4C��dņ蓒��f���#��RA�b��;Q:U�x��T��S'�;�Y���i��*Xi7 R�TF�A-(�O>?��"��ik�&���L�X�<Ą;��}A��ſ��C�.N��f\�Π�o�*Ġ�PؐJC�q��Z�����%���n
��_(�`h�X���Ak��J3\��:'P�u����\��$��sK��1`zKAf�e���?��=imY2B%Jgj��3�"JѲ��M�r���g�HJ-��f�V�~ܵ�tI�HU�M�(3��Df{*�8��h�ඐ�H�`��%����k�."9����h���;y~6��zu5��d�^~���$�=ՙ����f.b�:��5[�T��J.o�8��El�E'�۝c����V�8�+&$��+��I~��@_��Ь�n�詗]��I`�h��?���,����b�H�"*c�K�q��2��4)c�w����{�o|82��Y�~��%Ƌu%�����UDd���*,ߕ�-�z���F�6?"t�D��$��섳R�f�|ՙM��'5}�Ή�N�V.�s�3c�d�0�Y����u��I����W���X�~ȝ��8\�[�t�٥Ʃ�2�&(����Ci���P�� D����M\6D���(����̖^�(��h����;g4c_Jhwe�bU����8
6�`��8	-�W��o3'��WU���<����#Eo�<�3�_.�3(X�6�O|��
�	���o�ת)����$��ag�6R>��0.b����<^NBD�d�k��K��wK]JgR`U�,�� 9�Og�^�G�
g1���~}a�^G�<@�Y��Jzhs��~���nk),u�%sgǩ+�A�ɢ�pg1�XS�%�<��}��e4�׫
�)��:i�[īF�^��P��ۗ�れ�71�y+2M�'��h�@#��#�6� �nXT�A���I$�G+�({Q�*����*�xe�p�ک���s׽3b��w~����i�[�U�-�j�j&���1����a:�8��(���f�)�N-[�9��Ľt�3Ů��R؎)���Q�4
��:ʤ��[*A�}��[T\bE�I�1�4�`��������[��~.��Z��N��F�R�L��t[�Ꮟ�4��{派��Q܋S��Ʌ���Lu���i��oR����QNdkx���{�'B�°��>��\bo�|��I��%�X��kR�$�C{!"����� �Q�˲6з\Ĝ���
��h�J�Q�h2_''7**��` |���+�q�n�u��<����������G��	�)�!JT�DȄ��М2�K��(ƀA���4���x�����+I�R�;�(Ә �T5���C�R����2�m�B\�/V{�	<�ˌN���Biq���9K��c$XES���̝ol����Q��tNiP����b'A])�I::VX}��dS�FA����#؝�jh�F��#݀�3p؂���z�s>�����}'���I�9e�K�_FӺ��Y\��F�bF��"=}�;~K�V��I�琽�G�O�L�E/�>X癢~dj��G^�����'Ry�S�I|{���I���ڳ��![
D�X*��9��y�A��}
�����%*�f����{{�͵'�8�2���]����dɑ V�Y���X��:G�͂�P�ժ����/�:���f�]K��%XS�"�M�9��3�6�%}���	h�O�#����ĉ�Y���ܼp�n�Sj�`�`X|�-�[�*9p�6,��u2�
 {:�����ĺُ~A1��@\��u}6*<m��\�O�@?f!�#u�k!5~ʶ޵E������"�0�Sz��ƺ��%mt���ҥm����o�^p�����Z~)�7Z#�t����.�7�s�0�!��|ĈG\wvftm ��5��
Z����i�mi�bڒ�MR�Z��7(�Sj���V�t�1�S;P$��e�V�k��,�D�2�c��$�ә��D>�j%�|�!WG���Iûe�,�e�{�=�6�����X��)��]T����O���@��ө��nbݽ��kL�)��}il^d�w����-��g�?1L�*ٯl��>�Z�^B�KV���#��za�,��;��l�+��8�)a��D��s���z� �iP� q�f[�uű-�D�DJ0��?g�����;i%`e)�V���FKc���C ��x0�19:��V�o�RW���u����o��яk�����6�����������&�Z5�?�x����R�)2�xg�B��Ak����\r�mJ��
蜙���W��و�5}ⳍ� L�U�˦rC�9WƳ��:����A1��i����v��a����մp��	��/۩7�9֬f]��qȂ�{�4vopn�Y�{���0�*ӷI�E�퉆��e��F!6C����2��Kr�ʧa4f69���կ�aU�7n*�e�b����	5Y�HG� B6y��ި�r|c���1�2�����V�gq�A����q	�s0��V�e�2��	�0k'���P��c�*'�xd�jB������������^5��C��Z*GG���nm���� 0~�	�
�3�+b���
���>d��'�n��JuE��5K~����[�l�yC�W����&���Fs���	"Z3�C�7�ɛ���8�+T��^�����U�GT��ֻ�^~u�ϧ�¸]eANWz�i�/���N���b�Ŗrx�[��Qt�I�oSR� �	N^���N���T�p��1�P�n�ڑ���`L>~W�1���ZN��`�XP�͍0�t����?_�9���p�emT���P4�/*}���@zyD�SˁK�)x�Q�V�4�$yv3*��e������y���93�6z-7�����p�o��J'���m6ɭ�5�x^�z��@y?��L2���zX��L_h1��c�I�Ih7��R��Ws�p�௕��z^��֋��oF�A�x*�eU+��O� ���}M5ce���_����L��Q�z�p�@�-m���+�Ϋ���`������l�;��.\tokWϛ�y����1�nS���Z�rP��8��%s0��i8�4����<�{6�%�?e-5���p��u"����fJ��a����B��n��쥧i,W�!W�kX��aL���P��	~��Ŭ�$*�lr��9�K�����;՞b����d��)�w�|�����ƥCz|�����<_�|���A�vX�y�j��v& C���1B�	��u�=�R L
n.�I�R�9��MG	�ݲ�L	A��u��9��\��2̱@S_��q���M���Y0c-�-|�½bx�x����B��I��{R�v� p�{+;����ҽ�V�[����I�b)ʩ�g�<"�;���ޜ��C��M]��F�Li���r��cf�tR�n�Z3��
��9F�`;3�u�̿�&j3�o��%D���=8��W�{9cm�߆��y����0L���f]���\U5�亜bjѿz��'�����C�Y�<m��u���N����C�ƛ��N^��bIS�y�>'zm������?@5�Œ��M(t�͆�σ1_�1��U�X�d|>�����$`�f֝2�l�л��=rd�@3�9[j,�o�b��X5�-'���Ġ���y"����Kz��h����r=a���p�S�᠕��u��zQ��� �"fNg���A�G�����"�f���$�ҠIs[;L�)^�W=�Z���hek��+�W8P(�ú����V�<-G���,W+�`+�ޤ3�,m���k}��2���E��E- y��U�rѱ����O��j;�J'�{,�X�b���?v�k����g�Hn�K�z�XPݓ(��X��R
ʥ.����k��á�����s˝�g�����dg�
z1	h��#inQ8V�����&���4ѐiީ#u>{$N�\��^v<UؑjO����7��-h�:7w['Ydvї}s�������Ĳ���~�'M	�^��kՈ��B�W9%M� 3���Ǖã��v�	� ��l`��1��@�!Zv�yR����ȊCIf��V�&��l`�SF�!*DC0-������fYO.���������
ƙ�������G tɣ���j�s�o%�򒺳���ܝ��ż�p�yOmDW,(5����~Ѧ�Mo�\���qyy�Vsw�슢}�>����A�7U8���;(@�.#��F�����t�K�i����F{��И�����%QơfXD�]��5�M�*(���"R����X�J���[>�](n�b�<�c,]~Lb#���0"_��$\��e�/{=r��SBv-}�p��u���G�W۳o1�:޼���٠������I�}~]f�ٛ��#�95��>#�eR�/�M?5uЪ�/���Dy�|��^�U�:�6��vÑ�!��z�+9�b��<�7���R���-wI:����|�A�B�?�}�ח���F���|���9���W+�_nVF���"?vku�t��t���/�b�p,��B^�Os���,��6ik��WU�n�i��=���pqq��y��7BωC������q	B-B��ƾrr����O�Xϵ�����qWS��|Ə3����r0j71��-��i�R�}�Br%:�"��ue�ğk����mq�lS�[*'���*x�F  Ͱ*h������h�Zo������1Y�|�X҉��٤���z%���;��q�5���u�����X�>��_Ƿp���W��:��S�E�Iӂ9xE��S�r�xשā�SՁ{�������]����i���Grν�>T��3�	� ^������$�{WA�.]�Hr�B�.2��7�HK�����!�J���,\�sR�^X�9�")4��~���\��v�="2e���3���pu�(���E�A���_�ܒ�4��s$��;�-���*���w����M�lq^+��>|2@Ɉ���"��Wi���E�'X�3�&�� �eC�,�I8�/�`D����|(kY�d��A���^pō�!*��F8%]P�A(��?��e�i��}��}:W���M�>�o�F犊�vc%�(K�J0��Ԃ��9*	��i2V��xNe�0Bʉ�� n�¡vSl��-�sV/}`��Mlss(=�(�飲5L�� le�T�0k(�;�w'Ͽ��U)��o�é;�\���P��(�Z�u�1f��c=U�����#�3�A� e�gضn�Ќ�:h���*B��-���	SM�p���q<D������ �Ëȕ/��(��;ߊ)� �c�HyI�."�K���6`�ӯ���b�q҈vqׁ%��G��^OZ���3LG�Z�Sv�G�K=�E��j�J�Ƈ���{k�9:��ƴXt0�׎�>�GQ|e��yЌa2��tv���Kr;�ؑf�~ �x={M� ���}XT�ٯb%��Y��0���
@����0��ےY�gz�+jM�C���:U
1`�D�1($���5��)~.k�^&�e��r�b���%�_+$|��h�Q���oaF��JZr��W�A� 	�%����)�70��F����N�m`	N&�[��������mT���$ ���&x�F/����:k"��
���Z��}�{`t��!����f�灍�,[�*��Y_�U��D�g���#���$�H<%�s���b�k�����O5ٰil9Aw1N��Yt�Ԅ`�Q�I$�;�!L�f�3���3�mxf*�asD�/[� ���o����3��K�v(M,Y���wګ>{�S��ߗ\6f`��C\��	4�e�j��$�� }��	Ņ.����M{� �z���5WL����f�H߆�m���<)f+�;���
�w�[9'�"E�J[p��
*x�*�4��wE����T~�
l}�_xl(�O��%BY����nO����v�3�v�p\�� )�͏�~l��g;h�_mO��j�
j��X	��BI-~#��4��-���cB�6��CL�jA�;�C0;�(��n��:Ĕy�}.���Kf|�Mepuw�ڹ���������T)��j����;�dZ�7,G�v�Ъ��
�:?�_��� �
ˮ�3�%˲N��2���h-W�h0�QC)XsR�G�QK����'@kK���T���������l�D�k�3�l�J`�ZdgU��O"����vަ2�';��%jR��R�8+�����tE4U�Ly��Ώu��p�O��X���wR~�i��vxcr�z�Id#� �g�߯�t��Q-r�N��]R5����6̙r2,Q�[e:�DC�И����"��7���"Y��h�&��i���!��\�`<�ضh�����u���풐&�)�=�u���M ���E*�z��1��W��7q�W����5>6ݖ��(����<e>q���or_H������Ȉ�X�*��才�WD�
%WUZ-eл��طpe��Q!]zR��23��w� ����'�/)J((�Z�" ́�^��mz{�&/0��J�ʀdM�M���k���8;��֙��%��>cGJ�Up�c����)�ԯYk�F��#�C�X�1\z9�*rwf��l�J&�H(t�/��J��cm7��(���=����G�?�O~�5��+����.൱��,��M";�������[ft�&�7U7քf��+\����"x�n����Tk1�!���=�� ����q8�;ߺ
�0���F�G�|�/�u� �B�z��.X>�����+��� �Κ�S��٢��nM���a�G�bSF����k[۞��@�������GM�35��1|�̞�t}�8��Eqz�S�T�� ���G�u�Rƣ:ҝt qT�ki��V���%���⢓\�dDFe���_A	J4�5�'��h�k�.��B�O�]��@��c�5Xk~�R[��=YM�skLq1���ְQk�^2��T�����#��Щu1�W�{���U�`�}�-��?N��]޲I+d�LǪ���~�^�!w��ׂ��"є 0go�<]�����E���=����g��Q���7�A��4%��3���`/����{�N9_��ͷ�X@]z��~��2�T�k?�C��CН~�u�AIh�4��^`^�\�h��u���!@
#*'��\I	�Z��{�D�[���3:��p������u�ّ���7��-��z!jN=���rTk&�r��o�]�}�<d�v���..��H=���%Rc���J��t����Ygj��Fv�[��+S}49�8w�d��c��)K��<��#١ڵO>Wj� �Q��N�x��ׯ�	���z�V<ǵ�V�-GʖĿ�`e(.K�i�������P����K�c�eV��T����כ�d�ԬG����Ѱ3�Y�f0�K��:�� !�_�X$�\3�2)�1A�dܚ��4��>�~O�
+���b�6�Cj���ӝ½��\b�	��a�ԃv YC�)���Se�Z�H�k'A��y@"���D"Ch�/G��:�w�P�<�ؘuF!�5s(�l�\�hya��[�Hޖm�^�"{Ӕv"�ڶa+�.̇�mi�\,��A��Eոa���|i�/�X�3��y����E�4�����#�i�:;fdD�N�"�Q{�B99�ro�bK3�Z���2E���� ���F�M���蚖��G�u�y�[0PY|��'�����b�Q� �;���[�s�K[_~����$�O6s�Ƭ�a>�>��vE��.����IP}|IRt[=7��f ��M���p�u�3�6|������k��0k�~Ӫ��?�De��\�
�|�Z64�oh��R��(�gc�@_�ǅ�	�RZ�P[W�MU��pr\�{�L����}��QV�0���j�
G�pJ���ՂK����K��q$�/5�wKC^'�u�u���z��-��
�ςW�����~3x�գ�>;��$ʹ&K��5Tg	�e!��:�.�g'�KY"�p"��N�ϙ����{�m������cVR�@�'�{U�E�P o�A"l������-l��6P\�9�	���)]�pm����LO>mS�sq%�4���F�f�]���Z���	���&���d�C��A�ֵ ����,�L��F*��� �v��mk�4�fER���*Z7��@�h%z����$G���F�V��v����A����n�o���V�����Rt���aj�T)R�����NkU�ϯ-ƣ0=,�n3�c);��z��%U.{�ؔt�k�{IۭU���27c��j���ˌ���V]f]*�i[]��eq�&~�c�}4Bw�vJ�L�Z�`�a�YQ@���0��H�y�hh�/ �yoT�r�swv�����6�[¤�Z��m�W�XJ�}r�umo$���A��'�|})L�ծ�lR������;� l��.�4\�`n ��ߑ[O�ƌ��%�81�&�3?Q^Fq�Q[H��lX���}�_U��?������H�}"�G��_�p;�KM/��h��Ar�۝%W��r� ���^�{�Zc*r�[jp�����wV��P0�&�he��&SY���O�'�֧T�1g���U����c�E�����u�L)�Q��ۢd�sC��T/K�U�ݚ`�@=�(���6��h�dz�a�~q�T�5�6�P��?��{
�*���+q`�9��b#F��f�Y�ph�N8��ݯONu�SbÇ�s�%ZE�<W�vX���K����ϲ��c�#�~T2�PTDMWn J�8h� �o��aӅ�u;���t�퍞����Mc�\g�Q:�xy���ei�fF"9B%��W]%3P)��S/L3��-i�w���D�6��Y�������}�k�V;G!X��?��ۡ�b ���g�24 ���a����`g�W�:��yT�N��u$8���bX���(~�+�|�~j"/V�*�N��$��[���50�����W*0e��bϴFJ����AQfR3��G!+cy+����獸��nV|�
��$%_[��ŉx�yvz�6�5Xw��^.(�����A���w2�}�/=���1F� 8@$M�����F��Jfw@��hᰪ���[�OpŠ���5_�IE��L?�����ýLU0��1YlԂ�\�tk��r�,:!8֔^v�t��Y'���1��kMvwv0�d�yS0U��,/'�W
?>�2Z�M>��Ru���R�f�!��|����&3�������ٗ�C��lR+�f�-,����䂗�{�R���iSʽ���5v����R�U:Է�Nv�1��o�T�+���K�0��܃�|�P�4��Vvy9�}资����M�8���uC̎��N ��.���i����?܄�J����K�B���d�v��JG�q��Aic�!�&d/cId=`Яٝ����Մ�m/϶s��,�&�r�dى��*�P ��	^2��RY���n7���=m �PP0��'�!x"Dg�CS������,̌Q�����Zt���:+BK�͍�H-�ʪps�/���1~KB�aЫ�s����!������E�����$��{�@Ebpo���R�d��J�h�R[Tu�
+m���8:��[���	�ʊ.7�6p����wǖ�:�n��f^��2x��`\V��9���K �։��|y��C�J�����>,�η��n`!�2����|��1������$�����@U���4_H�g�Xw#)��QgV�=���0R2�	S ��hy�;�x�i7��/0��arS�&vs�\L�k�+�".�IVAU���S��	�.�l׸��'��uZo��/��;��+���rb�E�'$�8�C�2�*����/z��;�o!V��tR�b����E[�e`��Ȳ����H���f]�%�Er*R���� �pXtL׬/�.{�b���1��6N��M�����Ni��O6����	�^��Ɖ��t�	��j �"L^A	�������]-r��nr:�H�v(©�:&��E��L9R�x�`(X�2��dA��vH �m�&��Kc������)�v�
�+~t?l�9=�"�cD���I�~I7���Ի��v惜ʹ/(�*8�\Z��6����H��#��A79v�xqV�

�8�\�:L�V(�󫶃x��e�3/]rԎ�k⯋u$���s1{ԭ�2f�t�tԣ��=�����p=;t�W�#�'��@?�MØ�&����T�V���e�w"��.#������
#��Ҷ;_�|�2��Lqq`�l3���Ɋ�R+�^��}�CJd��y���R����s^9�og��-3����c��C��*>�*��n�(>݃������=�[J��{G[��K�z-$r����ֺ�lP�Q����s�e:�Aa_u o�Oe� ;�i����n�|Sr�@I�2�L��dT����~���Cb5�қ�r@B��<BJ�K�cl�J̽KuW��aFM7[q͢:�Y���!�0��dU�����T�n�$8�z1|��o'�L ���f�͑e[nn�IbR-I� ��n� ���>	�
�U0��������@�a�a�7����xj�퓯X�Wq��ؒ�:�.��gL��W�YH΋c�� w�d'�z8�Ae���c���t���`r)/LW`�>��R��{r[���{�8��X��}C�7Tz����7���c�p9x#z�
1H��
�r$a}�c]i�; ��xbn�]�M��U�T�<O�J��Ahoބ�|�Z�j��j�z#W*�
��.
��U�3�{`����o�)YVr�Iy�R�e\J;u�25���,N���^��`7P�q�������l�Y��]�iL�E�s, 9�&_<Z{���̙��S3�P�B��B�#:x��/� c���z��sv��צ�!����޵U�<*�"�{�<���UN
`��6O�0I�>V�������hM�=��D�_���6ҹC���=�A�������gO���x��d!����L���%#����@�2�>ͅ��ҡښz�"��ӐG��]/o+�؋q�4RO�4��0ߢ��<�6��ì4�L�f��NU��?�AB��h8�KO'��,�׉�3�)ԇ2P��"Wď�ظ�GD5�m��iq\�G��� }G���`Sr_є���WK�̆L����lx�k���A�=�'�þ���y����QF\~��D`��V�=�����o�Y�\w�ܹ�Ș�K��A9<� �kg�������r�����q��~鯓��f%jF!��P~ald�WP���{	��Mv�O`����-:B2BM�RYW�g����ӚR�9�-[�/[�!��<Ȑ�B��۞>�D�Y)�ˣ����Oa�{G�L%�;�)R�&�mh~ٿ�t:�_� �������n��G�\e��g~�����
<�p
�D�U��X���:��NԕR����cK<^�}.�y��s�N����|� )p�$�E�0H.A�Kd�;�v{���Y'�c�	�hj�٩)c�@9[�r�<n� _ެ�7=3�-� �b��a�������2����q�o��a{y&��V�Lw�Ii������e�n1|%��OZ����[A2	^�:��4�$��y���쒍���}�
�w�D�f!���#��8���n(Mi��1M���1�_}�0�RD#��h��Ӫ�`��:އuRȤRσ'hP��{��������3�8[
��d�<"�*>d��yp�:�f��sI�@�+7\���+�
b���������p����"�[�o�'a%oIx������o�TQ�-�V,P�4��*����!���;B���J�H�7cX�Ի�7��%>W1 �U0n�ϰNTJ2}T�c�=U/���ç��c-�ͥ	���ӎ[��(�*̸O��%�f���
��S< ���3��������Q����9�5�$�G��h��z�#�8��g�l�-��r�
l	 ^DfZ=np�FCW�n���X���pF�?6P���1�^л�L��s���|���X5>�1�z7:AὊ�[X�ѐ�jZ%���y�	���:L�֮ѥޱ1WŹuI��~��1Vm�����*���y��X�����\�/Ԯ-�[�0%t
#Y�!������t��#��9>���>5	M��O�,1�/	�=���}I�9u�d�����g).�ļ/a�����0;�[���
[�D�����%��� ��8N�E�)�&�f�|�J�4K�m�q�\�qy�1V�t�r���7�].��R�}�PY�}H�7^�b\�h��sC�N5��:.60��R7a�'�=vl��Xp�#Y&�As�AB�c��~]��� ��[Sʣ�j	�E�$��� �3��ߺ�w�����%5��Rx��h-�e/߼��TaQ�V˔�`a�XL�� �c8�]�]cO�)f�(*�O���P,8�X���X��׼���Z?��*�SLҬ�|
�B��Ad{՟8ց?�}��t��`��9��=��u����$�.��:����1�5�G3���B���IѤ%f7�j�N���	#��U� �_�g���ڢ��{SD 9~�r�;��f�;��uP4=�1�?u�j�#�C���=�;qT�B��+�}�묆���K�����́�W�9nPC,��gEy$�}'�������M�R�g����c��'���
�4��o�&��V��Mi�H��3��Z�������}6GK*JXIgf�>�ʀJk+F�;�ÈE�l�M�^Tq3����|i+_p��@n�Y�yN �9����7�Y�w�a�S�#ͅp6��˶��y\�c��<����M�
N���m�r�����q����������<'Z���6�]�\���ν=���=HpX���U�D��k�]SZ����A������EԠY�<�/���A �&<��z���2NQ��>����CP�������VJ�vH�TW�M�r�0�ސ~\�-���.O�I���]�/숭��8&�3D����;e��kL��=�e�J��.G�/�K�M�Z�*��F�N�Vka�D1A�]؍Û۷�C��aVRl�\gX��:��??��5�S�u���P6��C�e�t�M����Kg�������R�v3~����b�e�'14�KLo>�,����0ɪ�s��.o.��~Q~b�g0A�ؼΠ1J�%]!�|f����ΰ�aO����	���0zo�4v�썼����Ў珵��h2���-�Y�vq�2��s���ۣ�,�I��Ky����4 j'�@J1a�~O�&�bG�/,�t�����.�nL2�����L�}���nQ���,+^�t�˟2�aw/Oۣ�f,Dԫ�dG�m܋k�a�-8����ix�y�ȳ�Ĝ�w0�_8A �E뎳�g�akA)��[�����&��j��R�]:pZ�2�?OD��}�W�,?��U�.ă���h�����ދ�)��-���9p�vw�#%�i&HXN)��n[V��TffXGxvL����Yx1�]a��#,m���$&~UG�ƪB,E�?'��OmCaJ{��7��iɝ<�m��A�[&��������[2�8ߊ-�J���H4���4�\҃J��Q��Z�[� K'��4�'Eo�������<�,�u&0����q���]�/��ƀ[b*�t �:��Y0���u8� �D��s26wό"������Uͬ
�(͵�B�R��]�9[�/���Ap�a�ٲEךb1�P4��:���H{��F*���Q�����~J���b�Q�K�}$7	����)�9;�:����)'��Wm�
[[4X�?�7��;��v�j����Uaڣ7���5ڛ�����4Sn��2��n�@�}�����a-I+N¹o�`�p�޹b�D��LC������lm��񷹉5�Y\�C2y�0�P2#g�D�U71ntu��aP$��nǵ��D��ݝ�n�>y��L�K���-Н z�^]G%��}����ex	E;�xg�-l���R�BAk_xhS�QFt����`�hʚP�ۃ1̌�WVi�E��jӿiy�����y� ���2�� >�*���b�ۇV�J��"�)�ˎ�KZ1��#������D����5̄pC�쌳T�##]x=�W1?ʄ\��]�$�������#���_;в����7�%#eSv&U�]c���t����h\wY��O�h�-�Ȗ篘2�ȸ	�~a[����]�����]�VmȌ��V�86E.�r	�7���kt�J)��I�ID�UrTMg�o�8��T��i��5���2�PB��ls��/%��xAe'7��Ds�
e��䏒�2�����:����};���ou)SV�q�>�X��dK�r�W�2r��ϡΟ��3|��Nߘ�욅N��J�K��W�D�m>�"�
�����D^��:
N�V\�`���*�i[�����]}�|�QZ���0��6�*]�68��GV��92d܊�x3���Dދ��&>-�Eٳg��m�mh�u��
��[@ӲQ��U��|9rw7��Դ�6jo}��X�E�y���^���:Y-���#��԰�c`���~��׈[�'��f)s_��n��� �3������*�3�(ACڲ���r�%�}�tA1L�zC�� Z���}R��Ȃr~�����O�Lt���f�!���0���NI�p�=o7sa�&�zX�E���&�7���ez�TB���6��>ܦ�t�RΝ��U�2C�P����\����-����6$���) �&�6 +3�$���7D0� �P\=�3�mMT{�C�y����n��z�e�~: ��G��+�k"dA���w��mU�T�njVrG��6e��}"���?'d3P�	Xrln,������x���3�YT�	y��@��T1����m2�)ʘ�p4���4��a�	>��;�yh����vK�����EЀ���V�K41�4�u�zbB|�C��--oWaq��M��Dn_���'�B{��a�ղ1ӵ��N�>f��\xÙR��g��tN�����-��j�x������׏0.ظ��ptؓ���2�#�����k��] l#f�?,;��|&T��x�;ZZL�]A�A�f6�m_8٭zѫ�� x-L����a�8,�S}b��!z��ۣ����4�ɷ&�/f��U�:7�?|���?F9�'� ��ryɫ�7Ja��N9Q��8�,k��8�dUh�"�}�2�����6i��9Y����㓰!�9���<��������\�.����Q�E�ұ����ǩ��P6$W�K�tuu�g[lŏ��#���}1R	K@���'UyE|��ˬ߅��]���QLM��(�L�!�dNnG�n� >����т�P�$$���]!*��q0�C��`��&�_Ţ]3�Tڸ��-<�-Ն��ݟ���^X�/�����E*�Լ��+͇���d�S�Q�?�=ҢÅF���`D��d%��H}���.�P��{]F���7�pǐ�*톶۬��� Vp�7;���p�?n򗁝,�s�R=mř�>�2�4y�ѣi��G�Z�ppSȺe	J5K�b��;gF��0�!7z�I6��1���7C� :yq�/��Bd��U�T���j*/QN_�T��U�V����r�<�[��y�ϊ��x�m�]x�]��^���D�5��;��"w�~�����MO�D(��^����?��"�Y!����"�+< ^����r뾫�1б����#[q�f�'w
etk�a@4U�@NM5��8\Ġ��;��/�G6�Th������!� *�z��Ԡa�I�Y*V�>�=�̼E�"���15��W6Rk�}���9<�����fK2�J��D]�&Z�68�.�4I�tp��d�"���=]���5���g�>� >�6&�$�+W��μ�Kߺ<�z�gu�jp �T������x��\B}&=��bbB��X�H�ffÞ�J���Dt���[��p�X���[�zQ��Z`��)�����?+J�K�bT5��;��Ov�~����j &Jͽ�k|u�"�/|#)a9��C�Q{�}[�t�#�d�6l��|4�I�R��@'���s]��t�f<LPA����e�A�L0��9����,�E�QZ�r>ޒ1�%ow2���"��\Y��(��,4�Հ3�����	�>>�N7��\IO�$[.�j��5�\����tUj{G���}�:	�3A�E/�Ţȿ34�AJ##$c��';fg���v#�:��%���
;٠z���jf'_�
AD�3M Ce�u�3��0�E���)��Qm�M8��J�Ё�Y�
�/&P����Т�5�(�n��@�A��df�?��O"�$�L�"�t��Ƃ��}$q����>����5N�Η�Xf9;/���	�"<��כ��Ž��K���_d�iՃRu{0 �@�{Ŷףb� �=v���w�>�.�>��r'.�1��D�w�����n�q���f]��ĺ���%����䕾Ʉ�h��+V�Y��g�^?�@���q�v�����{��)���hH��h���7��X ��|�8��\�Bp�ѝˡ��\�gZg��@��q�A�֭;�z���Tx�7�
���Sg&ei0��o��7�Ik�����'T֒���T���~�M¼�D_Ş��JEd�3>��l�֞/�KH0y��8��x�2��6-9�~"tp���$��mt��F�4�]�jӚ���n�����W�?Ї^w+�$�(�+<�,�%�v��@�!ɨ�'u�ֶ�ǣ6�U�c������2�-�^�$�F�ς�GJl�l3�%������pc�]^|.��`
>��F<�:���}z�<g�!W��_�*���y芫�QQ��l�O�|a-J�ؕQh ���)��5�Ml|f΍��W����#s�Y�ޮ �q�>�[�u�~���,���D�ٴ�G���H���p��(f=�:V�r���=k����d3}X�B�D^�6�Z�:����,���Ѝk�6����\1k��C�J_'v����� ��'s*�F������|��� �Iw޼�r j�\�'I���Ȁ*���?0rJj|�W0���.���W�m��X&?MZ�K�Nĩ�(�r�$wަ]�YL��[js�a4iZ�;wS����O=Q� �Ō����^�n5;|��q)���E��}��I�(�1�J�8��F�^mUl/}W�U�G渁��}�vō���SB��Dw����*�QF�:�5�B�+�\VTd�hiZ(rEζ��,�ϣl� �4���8u�x���1F)��Rn��!�4��g�.#c�
�,	�[x�r�zu���M1/XD�c�[�[�a�
k{Y��k�/�9>����%�M]��ޟo(d�� �uB�G�ё��s��X� ���y��ɥmlvRt|�#��ިv8Y��MjR�U��1�͵�^`E��@�󜋉O�ʞ�D���Çe�9�b5���|Y���hu(&|KJ�PK9�[���yjB�Z�țe�ZW�o$�ifp�P�w����2��f���eզ�I�V��?��79;��"n����p�r�}�^O��.|˾��'�� �9L��{gB�h\�֫��ɻ; et7c���`���@BQ�� +�[�x�H̐e�IB��O"�w'1i�>��x�O��3#�5��Q����FA�,���I&�Cƫ�OH��wO���T!A8�5T/L����'����)a��_�nL��#;��¸��哄?�F�{�J�+:VU�8���a�m+)��tr���h�d5S���sнs5f�����!)-�{S������qƳH�ua�H�6�*<*�v�"$��0�h�V�z�������}d&�܎#��@��,|$LzI
}OA��T�#e� 
N�2�>$�M|��}6��No?� ����uY
��8�[���
+����7�����l�_"Wl�~���Փ'�SjO�k��.��N����eNT��G3.�y�wܨ�
�&}�(�k�_`��8�'[���c?r� |��F(M�1�`�e!�t�'٘��y�����Y���K�s�0ܵK;�"��2e���݇w؉C�
͟ ))�D�ڱ����F/�M���t4 ���MZ��tg>��y~qN���z���C[^�01�R�΢��O���^������C���6iP�����J���&%M�}�)��h�H��� p,�?�۝i����)*�7��ۉ���1F��j��;�\����<(2����R<�X���Q��K��1���3I�+�lM�M�;Ed�ڇ)���n3�ݣ@k�\94CY�U�Q��T{ �6
���)-������M��q����H�(�WL�{_���{��s	��}��!��}�}�]��5��z`�FV�E�k@�"5 "�D�^ߚ3{g6}"g��Ju�_�����$�f�4�R"�Hd��w�̳�l`�B�%Lf�7yc\R�,#����)=O6j�>�ў�����p���KvX���V_��7;�WY&�b��®�����	�G�46]�Ư�,u}�����z/##��Wup*����Y���Ѕ'7}����<�"��q�2��1�h��5�2ɥ�If-�L�@㓰�F�}^@L�&���Y:�b�#��=���|��l�hP`�����B��)�H.�7IE�~p��r��dt�P�/�'^9r �����
Y���V��!T���Q��iw ˊ��d��Kϑ���卌G�/�s�����O�,�V6��٭&+g�Wz%%��63y
�Iq��E��g9�D�b��"B����
�#q�����=��`�]`?0�?ʬ��a�. �T�V�`0!��
�.kV���[�1�Kۤ��dަ���C��H��z{J{��D��:@B�b�Ȩ
�NOq�Ѐ0N��K�=�y�aq$D_k��>;�|l*@S�����kK��~���YMY�!ᜁB�ޯGW��MO���U
��Z�)m� �2&yC�rnHon��d�_�K!��1�<R�~�L���k����ֲ�J�T�!N�	��%Ss�z�� ����2�)OP��f��!CqÜ���;f�7�b'-������Z�����r��9�i���O������v��	���h�Ud(�3H���`�����Dym����:V���Y'�w
2h[������G����G[�W��]�oDFi�E$����޷�p�g�z���-�I���!�z�ӈ��ݑ���0[v.��S�󐔇��w�j��6��Mm��6�'$2'�s�tJKRp���
�-Hd�Y�˖��4xP��CAQs������[6Vv3�obah ��b�:���&�F��������f��FF<��<���~�H�N��,^��P sÝ|���U���4����T��a�H�a��/��Dɐf���^�~�]/_��� 	��r��B�_�(d��.uɹ�>���?>-��K$9�d=�L 9dŀpa��{�3}s%Y8
�ۗ����<}�W�?�T�\Z�Hs{'S�7v�
\�po�ƹ�A��-�1�{	>���"L������~�,�ۖ����i<�0kQ�dj��9٘]sB��`���W�ս��a�( �b���DnI�8@��D�Kj���d��j�u�:~2�ۑ�� �_ÿ}��Zy��PK] �4�X�U�䱡%b�jJXy�����L���-L�1 ��V,ͅ��vёQV���폟(�<N_�D.:��e't]�o�/�̗ɹ>�c��,|V��/b�1
�B�5&��Em8:l�n���愻�K�����?���i��J�齇�lX}�U{>�X��P�(̳X�l$7>��ՄO�`������Q���>�'j�)�Sq�2��q1��y5ɵ����/����O�0����2�/0��M�E�3Z��ո�(>1f�P/Gßd���T�0g8�v[�B�;��5Q������~���8O�Ϧq�3���8�#U�y��lP�z�\[XB*d�wA�=�"QS��:�w�s�k�P� `�J�Б��gw��v-���r�Ğׂ"��xLR�3��+y������j��)��&@Y�<`m��+N���٘: Ipז�}�s��h�Y'V��LOZ���2��Q��ϊ��䝎Q ����1-7�G��ȥ7�P��|�@�e9q���{�s�.^?��yЈ+ل�VJ���z��pc�fuw� ��#�,bDeￇ�+D"��H�<O�
ł��O��g�?֖����uVW�WO���zQ���B�=Y� Lj���e>����<��51��%Ej��
,S�I`[9Q*�&e+>�/�Z�Dyrl/���O�BI� ��݂�L�F�H���1�:�I�wO���_�go��`�î"��7~�MK�'̨{�mq�]�E�+;ql�����]Bb�o�Z����n]Q���������Dj���!��Eb�7+��h,�
tu�����ܣ�-�ĉ'�i�aj&3P��wi�8:�#(I-Ǽ�.B����b���^u�U�O�@�ր�#��A���Y��2L����z�]����q��`�oz�x�P���$H��8�Uk	������|G�_	��5����5�y�⥃�/)R�sO~!����P�F1��}��5��M͊��6�T��,��xi��j��J?�XZ=��9p$U�rj�Hu�ш�t���B_v�����*ˣ^_؁��hA�¸z�~����!X�[����m���/1�8S�Ő��5[(���t�ǜ�3|�K-��U���[�}��	K��A[�qFJ�n�q+\�C�B� ��ܞ�]V?�aKBdj9Jr�i���,L^4�G�e&v�M��d�%u�ݙ9�640�4�[�����y�l_��]pK"��@`�n
Z�������C4>ul~�U���ZK���NO\�d:L���6����<�Cq�Q���x_gge$	\;02�y���p�q���S8z�P6cG}tr7�7������V���� �Y���-�8�������&b�"�K�zyes�R��U��6��7:I�+��zT1.[m��48�UT��;�m��䇣�UJT��ce*�CD=�`k
OF<�)mM�Z�{����~�_�u�������.$��[y��>u�T�HI�z�d<7�'v@��T�.��s2��Oѓ�� B�)��~-O�\����3YN�w{��f,Y�o'�u��+�,�.{Y����>C�daoF7�_J�Rx�hm�i��j�֥A��i��*e����HB7s 2I�¸Wj��>Х*'u
����z$�K����rc�܈�r�,�I��g�z��'�y,0�#\v�]>���_.�����'`4����H�Ҳ��Y���T5����Vg�d$	���v��2�Ԯ^��=/P�=��,J$�*�մ?����uŅf|�d)iN$�����acbi}v�Ĕ�:�y4�5r�_�ѿ�;�W6o�r[X.��%\�̯V�<��2�mdNE��gp �S0v�s�l3���B��G��̸o\.la�oi�L�O!�\B�\�$�ay-�nDӠ�ը���x=�C$/^����`e	�/ʃ�?����Y0��Z��4¼gpzfъ�%c3ݍ���4 ���<PS&�b=���m#�����)U~ZZ�ᦕ+gK#�j��8�	�?5�PX^b�T½*��|6�ܒu��q=� z�� |d��G�f�ɐ������B�pQn8Rb�3�ތ�em}#�?�\���P�z��w�N�4en5[�RXt3cBqB��I�דJ"!];!%�q1��u�"ce��@�U�q����q����+Z�PRn�jc�4+nͳ�^rr���G�z'��e�$wF'��"�ntf�;�He�����p%R���m��i���KM�:�����)����9�H/j������b���;fQ����bc���s�!(G�
��D���J�����.��r�n�1������G%��9H���H#u��l�)�	�M�"ۛ����*�eY��	�h�p9���$W��_��;H��{�P7P���k�!��F�%~M�f�=�J����'�'hf����� F(��F�V���4��zi7Ka���j�^�$�FJ��ca�$v �ɼ:�K���.<�^���c6�L��A蒓�L�}�v�M�M�J@? r#)B��%��biXq`�[���У��Z�n��N��I�>��nC��퀔�$������M���0��6U���I�d^�zk�-ɏK�3@�5�^�V�)T✻���q�� O�T𹍋��hV����xkI��ז3��A���S9�P<*����_��p��B�J�ʕkg0ɭB����d8SCK�D�;}�F��m�e�&S�#�}n�B�3�Γ�C���O<����f� u��`��%���N �e��s����L1�.Y�oSsn�X�����d���[��røt��8H/Z�)��un�H��x�����ΦG�j�+�u���o �U�C-��H�X���Ԅ���i�^}(�
�a�T��`�Z������6�kB}��h�;�F���R�j��a F��8���>�H�]��W�]�5�գ��	�n[F;��i1�V���: ��'��w��zE�,*��M���w��@}��>�.��/0�	E�gh�1�[�ɤ<"�+����,'%9&U?հ�Y�G,	�W�s�ZE��,�fS���K4���X;.�� T�o�@K%X/Ǧ�-()\v�s���b���8���4���ᥑI�g�:O�6{mǅcX�Ҭ{� �1z�*���^ȸ4G�y1	?�n���tP��B�H�}ֺ��`(C��`���T%p|�"�B������=�di�ڹ;���O�=����[Ӫ�8/Y��(4ډT5!�W	q+�+��E��A��ECba��7�#�Żzˤ����� 7F�b�x#ݑI�~�=��9Onnɰ��)z�%���{s���ؿi��i���:�s������U�	�˱|�PK
�"�"��=�l�})H�/��$�e?x� ��}�*&��<�"H�9p{���dM"���l�X7�nh�#)�d�9ED�E����/gW�--����ŚR��� ��d�񺖮�i|�uN�)���ucX��R��C�����t�]|�l��_U��1��d-�Ə�=^S٪	6�"��=P0x��Y���Ƭ�ٛ�!��&w��墷�y!�^�H3C��p��)���u��oUQ�^�[��/��w�Z9a45(iK��{������1�z(e1j�c9�����9
��P-+�� ,ơ!�u�g�<�9x8˝�n�0��R)|���PEz���?�L��mʧ�z\:1}c�쮸 ƶ�N)�au=jC���vS��A�9ږ��%�,r�ځyy��i���--<�3�H�և(݁J� �w���(NԤ|?	�ĩ�p��Ajҟt�q�UW�D�fo�<��[i�v��x.�Q<�8�����)�'�+�)T@[� �?5�]�@���X�#�̳�xx[�F�u���֞�5(�l���������4�b�����Ѽ	�8���5�d��XY��P<����"XEYtƱ:��t볡�y�2���l�l������Lki��=�Qa4�s� ���H��C�����(�H���,������)sB�t>��
f#�K�l��h�n�gBʼ8��8��K^��h��c�i�4�%�v���. '���x�i,�n|_1�ErK��O.�_4�����$(詁tH#�Z��|�������s^��Z�\k�!y{�m��[�z�E�!w��S�����0�^G��E@]�~�̊�!�֪CY��^�>�!�$��K���Z��C�:��5��� l�u�h��(��^Lnd�U_=��OI���o�@}-ߚ��F��w�y�nU�ԖB�1��L0��W�1�"��)���E�M5�H�� 	H7�)�p/��߮��h�ĕW���w��	�+���~�������dP��?�d%}��^�j�,���ܲ0Z��;����]�Vt6@.XF*�����~��ʢTx�6Ǐ�%U6����ߎʃP=�wOb�$k��@���M�2��-��ɺ�6��"�n�n��ū9��ۣz�yTR܌`S�7�< �8W��n��;]{�vJd7@�B����Nn�����ż0�x�u����:?v��~��¸������^&9{�5�M��	��n�%a�
�ܣQ�b��o}��~��7���AK;�0 �R�=���}��n�B#1�o��\���C���iGt�
�'�!�VE�ԟ��g�S�y�u�P��-��,�������5ZP��5}�m�դ ���A�9IVd�a���(����7u9fU�.8�'��
�ˢ�g������A͙*��I:"��tf��������i�4�j�u^�AO�*+e�)����z���o�6uC\#.�B��S|�����-�����s��y�Z�wp^%�j/U�o������剮T�ױ� ܲ��hp��X�Ds"��J�Zt�݁J�潥�"��։��g���G?��{�Mĕ�;��Np~��ٓc���常.W�Ԉ1�U<���<#��ޕ��0��}U���n߈��E'BH[6�w�V���ԓW|t��T|/_\4�ޥ���Up�� .�oc=ݶua�����>g��c="X���J(�Y����-�6
J�����ߠk�ÿ��=%����
5ê~�ʂ��n"
;�RB�)f���FYZE�1Tx����YF�!�T�����$�p�13���A=�h﹉��/5ݗz{"��K��b��1-��cɝ�^�\�6�1
�ٹ	��N�W�8�܄?W!���u�S�3 � �"ozn��)�9�a�hp��a�S�C��=��#���ğ����e�u�)�F�e]:���Ohxf.luD��v����e�U��eUǵ����1j+2,�Qg��@M�Z�����_�Om�Ljz=4&Ħlɴ^%�{�=�B��w�,��4~�;3��v;!M(+�#��\
��DE���C��b�-���CnӲ(�����1=�~�X�K��R�B]a!�O^���b=.�b�ZW3����<*�>�����!������cLQS�קM��?jUI���@���o�C�O�SԻ:�:3lʕ跇lh?��HP-�t�!��@&����J� /s��J�AhI�t���f�{�lN7��[H��� 7�ecY����a�᱄���?�|���~aV3H�j�R)��f�@Ɨ�\xQ[y�=��L-W3'wܧ��`��{��A��<����^�)��k���S:�/���0�ܪ���������ؙ��s�i
/(O=G6^Y��H�Wq�)qɈ��JD͢�r��r}��.N,�W?�������Q���-k���]�L���gd�e]*0G�Zqb�\T��x�M��F�A��1�4x �98y��獫��kZBv��c�����f���J2A`6�;G�.��4���q�t��:������"�y7�ȇCe"�V���J
��6WC�cg���!k+�/����C�;�a�,��~�I]��{�|�`�g��'p3G�7Q���(iCQ��{Tj��!J�U1��Δc���Zӑ=Y���7
H�440�}��,���zM�霨�0$ϗ!݉`���4V���ܳ��oq���JV��,!�(ԛw8G�l���4���B�
<w#([LN���޼"��)� �P��|��a8�D1}&�fD�ܤ����3X��cK���}�6R���<9,a���Tu�S�&���*xu:\pd��ԙ.RUk����Eo8��$�j��x�p�eJ��YӤ�)[��6+���>Gh)���jJe@^�bb~�������j�s}l�|p)Nk�t�֚�}C����T�3R��
͜�lo4˂����+�*����C���l��.K�<�/0l�>?��>N��.4��5�6y��D�E}���wO���Ĝ->�uc��r��)IgG>������*�A�&�ЀU3�� ��T����zs1 �+q��x�[Hn-�ם���3�!����\�$V�9�5|%& N���DOrb7����1�݉/UZp�bhؤ����L9�&)� +{ �j�f�ɰ������=~�T���Q��f�D�T� �u̕�\_���\�s�Zl���!������E��t�&7>Vq����\��<d/����y[:�$�����#]�O<��[��/�d7��5��xs^��6���mԶ�O�ACD�>��q;8���%X�ƥ+�s����8��fO��^��H0+��9i	�x[�������mE�F���{�&�_�JM;�<Q��\�Kc�e�4w���
����Q&3�cl�$�D�Ae�}��H�q<G�]В�8ʩ8 �g+�����s�L��b���NT�kT[G^'`���xH,蟥�#�Q7iU��̴Cѧ]��A}�c[F��a�������cp�*N���z8熅es�X�I����l������׎�P%�ާ�{w�q��9�*�8���D[��|���̵������k�A�j����ug����Rș�[�ƫ�㦓2͇�L_lNGP%z�.9��ҽ��K�?�\��p�f�����:������FK�gwĽ���}<��K��?����B����>�ip9�����k�wm`�p���"�(f�%P�o�Rs�w��(���ƻ�`g�y�	�:.+��W�ـgM���]ۨ�$DV_���v�C�;��Xz��n>:1�ⲱd'��������4���M%E {�l[��:�P��R���&]@ɍ�`|�3Fg|`��~���8X!�d����J
�s[L@��g�3rr�h A�.w�/�72&E`&��9���/+ܖHЯ�?�d�����=�ۓ1D������_YR���}�k��XA�=�%ƚ�)�O���V�=�a��ӷ�U�3�<�������.�R�T��s���1}K[�3*3�9��b9�-�3t�:�R��޸(vss�
�P8�)<���G@�!���j����]����s����Dë�T;Y�F�[+ �S�oup���|����Ӯ�螡��Y�P�s�<~�x��z��ܗ�-�h���b.��鿱�At� ��DHk�#��/&G�������G5�fr�$�ja���@m9�?J��zxE
_k���V�3�-&v�1���t�k�uF�l�y�y�O�:�����`0I/�)�N�p�Y+�^� �_U(׀R�&�5!��*Dp���H�I�a8�U�3�;���#m#�Md�BT��f�!Q����d[Q̔�^��G��w��H^	z�gw��g�9�[{�g�*z#�_�|}����S��9��-�-�ޤYk���&��U{5��%dn%���5B�Z���j;`�HM�B��CMы���A����mp��9�(:,��1]%���䙪g����F*bճ�
�/�Q&�!���H>�W�5C�µ�|J��r�Lv �¨��\i.]�7K��=�r����+ �ɦ����}�|�lKk%�O��D���KI��wco��&����]�J|||��P�	ޮ�]���N~\t034�{1��/+�Gzd�g�e�"�1�c��"��I�����϶�P���]����"����X��}f�����y?hbi
����Q=��i}��u&�����84�v�Rv�2�O�E�<�tBa�l1�'��@���۱�z-$��f(���oݍ߫1Ͻ�@���Q_���Bm{�Cߝ��/�oR��ي
����^#���;~uƄ�����|�K`��a�iM���.
f5-E�[���ś#d �$��죰bWO��(���YG�1a"� �Vxr�o��ۗ���J�sR�ySP�H]�}��5�
�<�H�Q�ֶ�^�3c����"��.F\��hB�1�\Ϛ�bg{f���U+��bĭ���?��_�Wm��[�zT��d�
������Y�P�4DI%Dʽ�ǽ)^j�u1������L"�;X��d������V細W����H:�h���[l�՘�~{�n7��э���3�X�F{A�1�|���e����7�͒�N2�$���1��ZW:\ ��1:Μs����#��}��|�6��#PM���o2���1���B}��b6�Y�t����}I�KL٬ZVTĠ���ݽ�o�rA%�s�+il���P��lLboc2�neޛ�S���v�mi�~��P�Xw*O2Pu�Ԏ�ٱ�:K�G��І�}�5�D/5���������r���$n�3FB�V �7�:���r(�y��3>g`��-9j�JB`6n��� �?.�;����^�8��4p�8�{^��������vI�S����N�=hqP����������K�+:Ə;�䖤s�KJ���.���f��3�C��^|����D\؆W�9�T��>S-�˂��6(����["a9>����BDw  J�u����3�4��vR�� g�H��&dH��ı�<���7�0�6��Ts��,8_Vr���3, \�79���L�c��&����_[foTw�e�iI���x�Є����]�D�@D	V����96��l�Dw�/�[��fQ��(PFV9�U��k/�I�S��b[�o���h��j0k����Thi���������� �3��{0a`�@a��KU�\+��\OE�ycy��-R4t�kO3�h�~З�1�䊄�M���'��䊍����w�TR��{��Ƅ99����FJ��ƔY�GͶ�ip��Y;�����2
�x74���1�R��fv�_����7��CjF�#�b.� ��h�D�-��]�u|�G��By7(��cn��/P`�x����~���#����?u���9��wޖ�읫��]!�^����Kc�n���d)�"��R�b߿�p����_(�9�u��H9zF��Z�.2��`m�ݧI��mဿ��$꼰L��S�Q|;��͗�ƪL��~���r�� �[ Do�geoI��I*b��������d��aGx7MV��~G�A��_�xe]+�R�.�^h��	)n����#�Wq�D~�3
���:V��|��
�
����T@t�+�Y��� 5����1$�'p.�f��Īd4,����lq�7��e1��niD��mk~���#�KT�纶�@���aU�w����."�q5�O}���u�P�)}6eW�]�\�	]7!��f^�|~��8u�B�	/��GM�d���u�w�4|
�?%�Ɨ�ԢLȒh�I�&�]3n�"[_���ɬ�mD;��R�o��O�;���1��4Ϳ�Ǣ�(�Iis������qϪj�GG'��*�e��Pym�V�ʹ�����X�c1U����0�##�XnF�mO N��Y�k5x�M\����W�X+�W,��1eZ�v6��HF�_z�r(s5+���hQ���*�N��1_'I�a[\1#8cM�ZXiU�"c�p���iY e!7�؛ լG��V���Ht��̬5�8'��gbCڙ&�^�p��H�l��u��>���>= )ۘi�k�,�	�e*�6����!DI�ߵ��c��ʛ����_)��lҭ�$o|x��	�;���netD�n������F��`�F�C�����9Im��2+*�E���j������;��!���a|�J^�fs�I���C���	�HM	Sˠ�(܌�i�x���E�����������s�u
��Va>5��$}w� ��F�MI\F�x�bӐ�\6W���t(EQ��Q���X����c��G�K�	�u�Cz���r��b(|ڍ��y���=;��3���-s)0�J�1���e����17*����0���Fy<hh���o���N�ϨI�㮌����|E�p^�^(�'���r�t�4�U�$vK�ukE�ذ���I��ٹ!Úl;�|Ś>�P;D���JSH�. ����j1K�,~{23�L't;1g{��©����G�Ml�T��'� �yG����i5n�	�}��t��G�K$�|�J���o���������B�Cfܑ���`�E���Cd.f����ծ݌��Z�K�+^����{ាƐ����?��k"b|@ك��:4�(�鲣�����?��~]�{�{r'gN���H�B��I�MD�(ySs�xEq�6ǆ�V�i�L��箪S��'1�����]���[���!�o�Jh0��DH���C٧����x^��B0�������q+�թU�O���G��&�t
��"��zp߃/�7\n��_�8K�Z1�}���n5_EՒ'S�i�C��n�u�'�g�->~)�1
0�D��,�� 2w|�8��>�����6�����mD�����=S�d�Z�s�Eg�.~�1�}2�{�ΓHz+"F���5vr�xb�#8�*/Խ��OjTa6p%_��z�x�k��u�n�io�L��ǈX\�+_/����oě��G��uΏ5qˏhq8�H~�ZB^I���>(k1%i�
 ZQ��D�ˤ�ߴ\pR���^$$����>0�tJx:���مI��*�#y!J��L���{30]�6GO��b[�[�`��+}���P*YR����B��C�):�p7��e<N��*���2L��_1���<��'�}n��M#���@�y7��R�ރ��ja��N@�1�I{�������*��EϹq��H�4;�o��^B��W�AM�x�k���L�0Jܬ����'��|<�j��}L0�Dŏ厙7�c/��6ɰ�[��ф]ٽn
T��"d���R�d^��G����.��u��N�\v��T�oMX_.�j�(�iJ�)�&t�+oZ���\!�k�K{~� ����mZk��L:*F_��[G�WJ����e�8`\AQ}n'��O�n`n9����[�D�{R�f�BC�]�:8��<����L��4��� �<}��y�<Sxմx�P*j�@��n���$�V$��lQ,.QWIbV���{A�k �Uº��I"�q&WZ�b��GR�-��3�-���F9l�E���-���6�?�z���:���;}�E]U�q���P!:n�U�=㳇�,�K��+�[�_���.W/MG�<�o�s�(�	_9��M��vB�dc7WnM#�6.}��d��P��Gܶ�B/�{}i$Ӣ-���|�V7SF�ZAH73T�ɫ����r����ܴ����(��n�@���gñ'	�ů�wK��D%���f�+��5��K[��|������}{S|�$�^��6�I<�3SNW�L�_9��G�w��MP��ł�/)]��[+2}��^]�o:�w6tT7���׮D���sp�h	4��ţKn������妒
q����LYk�+��0n��hR1Ϣ�����g��S6����n�k�&��&9��e��[�$8��)�'l(�����>�v�kq7��T���e��4��4;�/v4�vp�[>wq�ΓA�ζ��V񬏂�\�]��h�܏_R������^�����t.U%�@GBg0F�`٬*�2͸W8��m�?�߁<Z���3�+�T��8����R����ՂƩU08["��Va< �4R7tcUUWȁ���R�RV�	R��vV+0\jL؍�9�K���]P�� �����J���cS�G�OG2,�gרg�Sh?;^ϒK]R�g�̫�q�Iןx��V�%iHe	p��}�����v��tFE�}r�r��*�8����+�vFr:��w�%�:n}�/R^�����G�V���:�+�����f_��w�6�D�)�������G���3�rWă�N.�G:s<��V�X�/@��et�{����F�aR����(��G��SZ�ix�&j�	v�Yl�"�iw��7N�scֳ`�2�����_]�E4�iP�����񚣆?R��o��W��A�.��v�+�ڏȎS�W�.v$���B�id^�V�Q�wEdӸ�:�z�n��De��z�����F���j_HG���y�|�0�~�3(��M_}��.�W������2���M��(�Dd���+݆�4�ڥ��v�#�~y��G�����������������y�]�Qz��uMo�g]6����+��U��۬=��l���P�U��`���F8542<ׁ(U�!�^�1d���>߈g�co���n:w�����5H`b��0	�1%�N�$v���.[Gm�(�VLh"d.����<�9�#����Ρ��O/w�Brݗl�<Nc�&GL$m�(e� X���\-ݟ���T�WȺO#��N[��ϫ�2���F���)��cF^���؟���d"D�b�&��#���jj1Igq�,��6a��%�����H�;�KV�r��:��1�� 3�;�s���N!����I�����v�s%�PA��o:]Ά�h�7V^wh�L%qv�#�Ep㍃����	���,�Ջ׋�����6�R#\o�9I��K�=�Eඣ�e�_�Ij
"��5i� �����54?��� M �M���ѩ�x�^,�>����wϙ�2�af�B��~���V��D�g���刓���̜Aۙ\�n����DH�M&!��Nk��3�������E��X�>~p�y��d��Gz�\��m�&�X;�y
N�F�����ߚ�6mn}�˖F�)�Yx��ɴ��ɥ_�@*_��S<�u�`��4A���������x�W ����垶�tτ��؎(��z+8�E�efp>��{���+;���q�g��e��$z�
��fVk��}[P��1b�a9~���. 9=>oo" *����yf%�h�m���ilY��b���:~��'�}�j�S���6��ɺP��!�Ch��^��A�X#�-�Z,jO�9��MY�R/�ee���oi����8l��ޣ/41��m}�5z����g��� �:Y�pt�W�/��Dv�,	��̧	8
��-'��W�Wbh��o���ڄ�s<�A%��]��q���%E��1#	RΘrŁ|�����\.LRp -4�J�?�2"��F���g��k�b:����]���P������|0,5Gq�ߒ�}�t6�'��7\�vfC �ޝ�5�c,Mn㼜�q�փ����~_�D�"+N�z��ZUnT�%uv���9���վ�M��:��l���e��p����bT�mߚ?������}읫0VԮ5P=~tK, ��-n9�ѯBՐT���E(5}+��b�����V��>��̥��a�,���� �9�<E��?؊V��[�y��}�����e���� ^���f��������x�j�d�G�+e�'cɊ`�)�g���\wMҾ@wP$�Cj\\�̏}|�g��B|�;L�y�ӳfD���r�SVT�F!}��
h8S��=#'0@��B5�{ƴ�L��#O)p� �0f��$S��/R�Y�
ƞ�uj�_ڣ�L��ڧ�a�Eb�F�ļ6�Xa�Rbu�j<�_����wlwk�:�h1�t���P�K�g*,�F�l[�ݝ&�'&�\(o|O��o�${z2hjn�a2R�Q��WOC��/�wkl�s�$��1���#�����P_�"9�/������'��wK�-<�.M$����m��:'��0��4���:C�?�f��m���}m5�8������ ��|��-V�ukJ�y��?�K���Y�F����F�q�?�ڙ��wip��&S4 ��
+��j���H�j�"R"��Pa��������s_\����P��^�x�Oʫi��/��'�!]h(�+�/<H�5�� �~��c3�uO�7r�i�Z��FY�<����E��q:S� ���Ӹs�g�y����R���Da}M�_K��Hͦ)$P@f���+���x��>̄�z��B"�����B`�x9(�S���v������Q���ܾ( �d%�(R��?+��g��.�}}ϑL��ݥ��;lM_�E5O@a�Ae�V��ʫ�X/��n�O���Q�;�z_�^���uP-���e:z������_��)ڻ���8P�s�J��z��R���дq�A� 1�q�' %�K�u{j	��=d�}�P?�?��h,��}�0 P�|KՀArj����f����N�0�����|���qqj�6�S����\Wl�w��ӿy=c��˚��Y��15���.ˢƸ�N�݀���>*^�;�����ީ�;*W$�:C�0��^�\��V.���]UJa�f���]�e�u�_~���Z0�Ap)Bcd�Y�?GFRf��Ƽ�I�n��������e�2�kE�q�m*0��cT����O�ak�(�+k?u�8�K�2�h�6!�(�Iz�����f����7�E6��s�w�� ��?Ct�C�7������xr�z��
��lUU1�唖O���{�uK���M8"����'�9s.S�-���	(t�(Z��7���ΐjZ�y\��r;�	�U���C@V᚞��}��5�?�m�
R���]�f��2`���T4[<���NN'����ɓ�[�vד��g�y)Α�Đ#�����Ty?GF���,vܸs���t��I�<��� ��6�j��+�3�AAI�54�NJ,����s�[��͛��eޜ$��6��0�3؜�`\�\a����M'33��xO蹳[	����vbX!i�h�������'D@f�(Q�YJ�M��Ϊ����}z!I�Ą�H�G؅C�Ö�Q����i�vyf����b2��C&2��@��1��J����N�6wT��N��+���Uo7�;�`�R���ǀ��%��G�IC�#6�h����A(��}��=��M~<j��T>g��N�V�E�F�dxw�H�I�_�9��zp�7�v����j[1®M���������Okl�zgU�V���ViX�.��	�����_?rY���GE���\���R1��O�l+�@��*��o18��RG8�p�&���������e��>�S~�+�v���>�.'��	���/'+��$1�Of�i��Z�ͯ�a�L7]�M>���P�-+��m9SN�!�W�]k��Ftz(����c���T��^�
��=s���^^����� ����G}�]8=8�������샧��<�(S��窶�����87�U� u(�c�����s���_�G�#:#�b�&�I��a�f;`6�NZ���������
��%c^Yj��r��g]���;>|�(�4e�n,�p�J�,C�B�$�|{��V��A�����*7\)�����,O�놢Z��'h#k\�-f�0�P����wrӯl�s��k�j� Ɋ5�����<����΃�J~�����	
�&��k���h���s����Ojk7;�2x�p@�>(aHF�G"���f�J=8�E>eX�A��ȴ�;o�v�0XLf&?R����>���k��Tr�4T7`�ۮ�U�wD�[���	������ ��/X�����.j?L��chR��%���'�E���	��e�6�� # n~�G�����2��N��t�3bT������w��]a1�Z�n�����.U��W��٭ǥq��H�ڢ�ս�>��k1NR��C 9��AL3�#���A�j��!�!,���O�
��e�$��� vA5�9���������1C�˗ȕ[" �*�H��)���j���U���n�I���Ee�Fx?o�y�gz�
�xD�B��<p� ���<l�l~DpEf7���ü�@��3��f����t�u���z�`;�p�8}u�&>5�iJ�ݳ�˘m�O�a��^1ؙ���[�FH���oM�"������%ϕi�8�y���{	k��'���!�S���}��l�$�s������^�Qgqz	�>̗h���[�g�s�4�UӍ����#�E�!���dy��J/��?��RH_1��s������EI���C�,tKMH` ���E�r��x�A�����.�CV����k��m`�pʯ����+ ��_Ň�I(�p�V���)c�i�0hd��
�_����-N�N�ב�o6�lD��ʷ�2s����y{��Żb�-T�AdE�3�8s�Ҏ�M�~�E�>J��C��i�9���W������ �`�G@��4�-�:�
|�~=5t���F�_��W_Lڀ/1;4іb��$FP2泒0�n��i��me�$i��������5�?E�=O����B�[M����fV�q�j('���}
��>�����X��&6v�R�*�����R��Ʒ�~ZB��\���|�-�jIҚ� Cl�.�jK�HOᴺ�I|����>���49"r����y���o�x_�t�5?���7/Wc��(��{��!��D���}�T������L�8OX��oB��0K����J?X{N�),Ŗ��2�4x�O&f&��$]����F�`��-�q�qxB��<n�1��(��*�B"��L���~�2�ƭ��P�I ����αGc��i�[�5K���Q��̕�@�/U�6g� cUQY�74O�]�k �B��9B��|Q���-PYp����F�@��#���rd�mM�g�;�=�Y#k9��������-n��m}���l�o[	�5����e�O?#�V���j+��p�py��ؤ޳Q��P�,g����2K��SA�̫����Z�������M�`p�ֳ��2�Jo(R�o	�1mM�`M�mPE'����t���a	�+�C�&\��c�)}K+��[W��{�hXy��.�'�eIA|�{�ZYޑ�\]
����}N�tMԥ�g�?�N��q��($+�M��)�$��ma</��m,�ds�4B�L+qkO ��]�67�����(d
�u��8���eZ����,���$����v_�"~
�B�J��s�\&t���[4�t5"�j�]7��n�zw�	�ؘ�苏��?S%��J6�v��oK)�m/�4f��Q��SMh�\8C\P�$�K`᭍��K�gY�k���&
%H�YK�gJD�b2��T#}-�2*m�5MKW�*�A5�++��Y�P�H*#�T�z��<̚��A0�q�@�d��ߛ��Gt}v��g6R`	�@�Yo�<�p�+J�ᰒ�<+@�[�8q+�E0����:�D�ḧ,h���9���?=��� ��C'9ƦF�n��j�z8��^������L�-�H��1�d
�B QI[���M�<o7���}�W"Psz<~�rfu�fڻ8�ʻ�$v���4��׫pMb���=[�S>-|���0�P� �����u"O�ލ�A���+k?��e�V2��������8ǻ��L�-�:IіN�M��A�@�$��wY)C����j���LP9]?e�B0O?����%x�{f�QE�{2{�nDis�m�6�����Ȃ���J0���O��D2��/yP�w���ƐU��`� �,}�&;r[s��K��k�0P��P�`�tS6�[��l������9�G�߉(�2�3��羇Fi���:�Գ��ɑX��I��Ky�gSO%���)[�2�޳���X�Kw���#>��;���h|pyD�6H����<Ez����g��}�WҊT�ص
_�o�|���R�4Q��u�\Di�_�2�s��ڄ�+���"ۥ8�o$4[����{��@)�^��`�L��FrY��˭Fvu����	��V\�����)aR8�_@�>�K���R���9, X2'��>���|����~�g��\��?�q&�*��<��c؏�~ԋ�q����.����3l4�i^�q���*6�]�3aa�qԸS��&GvVh�B��^�ɻW�H?�ʞ�X���Q�6g��C��M|}Rܡ��o竄��S�߀�=�ʆD:�Bc"�-�	� �E%��5�R����Q����G�ü$�j�L��QK��vnZ�ٚ|�Cz��R�\wn[�n�_�A��ǖ�-A����@�z�?��L�Qs&�G��ߵO��+aͨ�z�U���]p_Qxպ�`���K�/�|)v��Ϝ�W�9��zov63�+m"�]��?��.�
ԵR�g�7���c���Y��w෡���\���
ޏY#5i)�9�5M�����0�5�Z[T�F"��C ����v�l�CNw��<%3xp�J΢b�u�Ӣ�w��H43[.�2L�j|��0��d4f�vl�]�T�M9�w�o>�p�ߨoԱ���GwW~d���H�mdd^�z������'�3�����fd��͠Ӭ1T��P]{Z��}t���QxC" ��>=V�]�&��-��x� ��xUdE�`������mU��
���5P�&9�Z��3�22c����.���%#�xl�-�i~������Q���>|K*�>�����+��4�/�힬GJц�n�#T˳�ʵ��::�˧Ä>��x�3��A�cNL���6�L�%kfg��>��3d�WWm?����_���_qֽ���z�D�'h�v{��?ob{f9�X�&�\��RG��%�<+	�ӘRd��)������W���F�@��aO��Vw�7#M�N{�!&:�4 �;|�=��G�BU`�Eo��|�peNXr��`3�%4�J��¨lct�v�/�QC}ֿ�U�1*�bB���g��3�HP� X�M�Y�2�E��Xx!��Դ8��M}���`��n{�'��p�z�C	��Jb��w�wX�^sc��R�`�����RŧMP��q	1ƙ(:\��Cq����{�?������|�Y$Nc�U���� ���QZ��)4~��J�J	��p�{�Bx�l�@�VV�7[�KL�?��㥃�LD����t܋�,Krű+
@j�8W�m���x��q "�]��\$�ۂz��j�7���U~��(*��6o�CX>ΉE!��H�)1��>O�gl�%�����R�В
 ے��I�t�K��h=#&�S5� �Tb"��{��'�4u�)G[��M?oh��}���Q$��Brcj���E[�s/�t)t��4ڦ��
I+����R��ŝ0���W[b;�[~�P����1�\}�;�U�6��쌷�[�&Aq�ـ|s�V�:����1�J�?_}f�Ö wb�ɂ7�� b�iy�����s	��|���-�h��L�Y{N��G���T�D�,j�CƗ�E��N
�\���8���1u4[�𫿆y99� %�2�
��6�ǃ�p�B�;2����
���(�;�|h[h�7�҂׶��n7���U���h!a*$�q��<U>�I�D�r=���F���x{
2�^�p���"ĕ}u-D��U��n2�A�MxN���d9+�ڰ���Ǫ�b�x_t��.�R�?4�������J�*��#��8 �1讉Ƨ�(�'B͞��A2�]9 ��1�؆�I�gS���9���_�%ܮ�1=�ZB��18Z�����z�B�^�!g�=T���rrSv��ə;ð��_<.�����h�|�5X&���fbQ�h��9Pvɔ�C��_4�$j/	H��6���N�IT~��wѮ��h���i�r��;*��9����q9�l���oDe�;3$��=b�O!��9��m�+9~�-�L-I�V��ȏ��˭ԥ/!O�:�zP4@��=�p��;�Hq'�Y��d{�F:���o��U9�n�V��8)���&�Q��[)��ّ���dy�!��-�\ Ad�*0T:�!��4��Dޓ_SбX���=Վ`@Z�W�A{�z�>�O ���c$8J�iu�t)˥[��<���Ma�n��9�h�QjYX�J��~i�v��C����;��=� 2���s�սC2,�Ҡ����,�����l�Moz�����M����(  ��`���ے��� �"��Udu��<�:5�e�sJ�#픹ڐ?���믙�(m[���aNo����} �`5W�"��P�g���x�*��r�`8:&��:����q�Y�UF�,�A|Y��=G����ϫK��raA+�֟��Ң��4w�����:�%czSCd����Ў�_4�\6�pΆ֬���ז���8�8�'.T6`�l�QR�\�c���i��ňS�^���=�����j�U���ɰeo`�($l'�i��3(�g����6��V��T�E��VW���2BI��]���^�m�#�ݠ{Z�����;):�qzƋ�h��!�}�!J5~�s\�-��wG��T��8�vR��T�'Ɵ���v���`��g?K�R7˾i���nA��z��Hv����3&���eX�H�7��@��c�6�J��=]i�WءBp#/�rNM?�k���@<(�ݜ8\��&a��,(���r���5�YO���:�C�	cה�[-_a���ϔc����n��V�� �d��B�������*�H��׀US����Q1b`�[X
�c j̛�6���͓&G����گ�}%x�Q�ܤ�Ap��v�M}�&8�n}Oe�)�Jk��]��aFߒM��15���K"��4�FQ�KߗLD�?�������`��F�@v���	W����U�ɿ�u����;h�A�1p���d5S��������:�Ի�w[��_uX���HB��ivH7�V�-�	�A��Ҫ��3�rg�K��(s�A���e�G(VX��W����Df�f�4�9yI�����ioǤ�P3�ԒV\�{�[V�q��	��{z�{�V�Q����)��?�YBؽ	�/�|�w>-͜�r�T/.�6?�\�.To88 O@)��� ��'1��
����V�?�ԝ@ V/[�m����nmG�4�B��K����܈�7����@�C��F��8�`�ɇ��@�5U��c���ͥ�|Q�?�����ɧ�8٭��Y���Y��\�����.��棵�Ԓ����õA�Sk��/��+��vb] 0����Q��?�0�q���!���6��%(m�$@�G	[G�h��m{�y���<���2��R��:�ᄾ�e0��=� cP@���^6��Q�K<��`5�J����c�b�~�a[��v�7���=lz򝪆�X-�/�o��Љ6�n��~�D�{w�R=cٰQ/k�ZדN`G)�՛Ry��
��>�4?���O*�'Iw�@ ��E��=P�+��z�h 08P�V'=����u�H�r��ݛ�Wn�r����!�IT'8�d��+ћ>�u^
"U���	�E5���Q���/98����2=����eo��k�(F��dwH"z��~ۗR;'���b{�0��Y�e�uz(u�����MN�$C�����]�7H�8�]h���4t���X���P��%
������=���c�P��ݦ���g4�F"n�)A�i4���S-v���/!#�[6�Tk'8T"��w�Y:�!��ᅋ�Pݕԏ�����\2��}*O����d���V-3ɡ��y>����!�zu�v���;Չx{�:%��^�Z��<F�	�J����� �J�)�Z,���f���U�e��Mu��g%�'��6[���j�-_����A�\�n�(��Hi\�]�LٷI筷�����LY�7�oD��ӿ���Ql�� �-�ۛh ����t�(��q�0�����L�ADh$f��LG��H���,���	����F���#)��x���:*��LKZIOױ��&"�>Q]�������R�gtwU��."i�u���|��d�Su�5n���3�5��}`
�L�!P=��������ϭ]. �X�Wc�W�����N[�����ƵF�� ����Yp ݹ��`��5r,S8����K}o�8%��:�c���h�CA��K;��Qwz��."�{<rBb�`7�2�8h��[��x��n�g���L���0�z�����HzQB��Z�A8�/�\kA�_�4}����M�c3:�|�-{�^�]�G���B�����HL���8���+c��9F�?qڒa?=�v%��3!"64�]C��
�ΫZ����H��FB%,�9�e�k@��ʪx�s �h���I�ӯ������<9X�c-Y�M�
�G�r�>��s�0�lhڭ'%��-Ѵ:�4�H���wM]�UT/́+zd�kD�Ʊ�K]��8:,�yz�d�X�Ҁ \��3g\p7�A�|���	X�k����<46�{D���;N̈́G>O=����&�� ��F��O@k�^���z!�e������.h��.��_�nZ��5yw�4�Pԙ#�r�mkĹ��^�To��d!����,A�1�0�{�?�Ĕ�u��rԔ�`]�A؁���l��+��B�&T��A��^Gv��&,>3�H~f���i�L���)�s�醝J�r�!CJJ�K����L�歵k�k�9��]�H�9�P��\>�,H�n�]�!��D�O��[����������;���V�:&f����gLr�am������&�~o��=��A'_����:)I�L��'e�!��w���o����LVF"|�0��=ѱؕԑ	@���s̃�/���h�h:/V��B$�g�����w��c��w
5�;v4yu��`wܢcX����[�6^yZ~\\"�x�z)��d̨��~s!qd@>��hs
�I�.Q�D�j��P�7�0m�;�'U���rn�N������#�./8�~�d���Y�"^��P&+95�^�Nh@* ���(��y)�t�����|&�4O��2�|�
���))�Z&��N�E��A�
w)�1�1X��@�n�e�[���y���(ßh��Q��։�����opa���*�븄Dd���]a��i�,K��Lv���ܲe~�yvi��{�`���B���K-N��Bm� {�j�/>"�]���&[ZRh��}��?/�b6��w�����+��!ӗ*% �����z�ϵ�'�h9]a9"�� i��[�O���1�^"�W��φ$����z�?�+]��RO���Цf->@II��k�l!�?Y�ҍP�lJ������7 �+׹e&��K|z�������!yE��c���p�Aa�ma�	A˳��l�Fk��1O.<⢳�)��o��x�l`���eo�1�KB�B��|�$�`�T�g�>s�s�[[�0�a��7 �����
ɢFw�S��FX�]�䦌��FW�k@�e#n�!L�	�@Agȇ�3c2�\�� �SM����גuiB"VA�����08J�l"����Pt�̫�#<BR_(���f���꧞xU�83k��4͆ŦR-������e ��j���A����g��>(���{j*[A\�I�{os	�$C����B�2m�[X��Hl��f��w5�<L�u�25�.(��(��\N�o�v`�sc��BVoE�f��e�8	��^ZSocw7���e��>lW�'q2�^���F2M�N�Kq����;�^������[�h�*l���O�#���AE�nh{5��)t;�<|b�^d�Yt�T3�Z¯͙c#gw��Z�rY�"{��-��YC�p}:�\�ta{��y���9Ƨ݈9	�9dA��Q��\e8o��]�y��Dh�4�{Y`�NO^~���J`���l�
�0tD�sڒsua�B�"���X��膀��X�b�E5s?���q��	gM0o�r� D�\�{] r�>lM��l?;}и��{��Ţ��$�s<T��ޡ#:�kX��㌂��QB�)�����<��q�����`��I��қo(�4�����e��ߒϬ��v ��O�2u-ܩ�|�z��0&���C��5R��\�'9�����{B�o�I-���\�N��2��_v���i��Dբ�*���D��bGE:�>�D��K�:��[O�B�9�(�K�s�Zi	"����hi z�[�z���˯�ߙ���C�����9A(�T�s6��/���j�y���!�DS�����PZu��#���7iw8���t\��иO��e�X֣Bi�'�j���QC�<�OXs��j�U���1�X�QN��wJ���L�U�HQ&'1Nӻ+\���S�w��I':D�����	� EɄ�zi'�'㲆�c�HIn��lgͮ�����~��*�`X [)�T�qm�h
�wa$�K��.��3��v���V
x������=�@�Ym˲Z��0ޛ�`�	���\��{����벴�|MǢ�0?�k
����dа�#Ð*U�M���>��'f���k3���$z��RAߴ�,^
�2]ĞY�f��b�_@���Pc1u��Nΰ�1���3���t�,����݆��R�؎p�wR*_L,k'1?���^�q���H�9�����3���3I�*��M�^#K��9ZSd�ͧqu�S����2����&�B�О
2��U�M�^�e\�@߀�Q��=hH+������҅|Ue^�5���N��%�<N��C��FN�[��R�I�UR�	xr��9�3g &�!�G� G��.R�q'@i��zA-����CNWE�g��� ���)�F��X�mP�Z�qX ��GIbtӲ�I`G��&��4��|���
�aٵ٢����/%��7#�F�c���e�M�"`[���MM��}L�1�˻�t*d�ʹq&ܖ�a��:A4'�����&� ��V�������]�%\sNw�]��Q;�)v���YԂ]��`��sC2�>��e�X���|����Π+����k}�o�3���fα�\�~��.��w(�;��YheT}:à��_����F�#�/T�Nݳ\�ʣ �;�T�����+�L��f�,�C�ܽ濈��>=�W�WF�w1MFyCSCǓ\jr'W
v{��e@��ػZ��@X0<�^��[�Ճ�M۫_Q[�2${���26׀u$�x�V�͏��پwRN�O�n�Π+���bS�Jz�+���kM�Ls,����V�� ���h�i>%�o��I���fܘ�!pJ�=e�a	G��N%��TqQ/���[�l��~���2D����'�X�ӀR6��4b�n���l~���@7�{�
��;&2^|��U4'��t�7(+4x:|�n�;%M�	�L
���`e6�\�.)�Y0MY�&<RIe��œ��ȶv^�B	�k�S��/'�G���B�L��^Owh�W3��x�˖($�ag�Hڬ����X�E0����YQ��)�o���{`�¤��:4|�e���(b�b�i�@����@��<��O���	�����,����}3�3�o��}0`+V"����5��bg�eo;��͉��0n���й5���~5�d�|����6}4���Dۚ�.�&�N^O�:�����K@�1#J�K�lo�����>���ӹ��m��e���.�C����ф��B�j�z��Sc��aTn�E���&���,�H���OIy�h�.69� Z~0Jɽ_G����	x_��~�_2�����[�1$�AV)�#�ݔ5�Sg�:������QY��8�~�#'� ���r�T�����l�[�^��|�-��z�n�����2�H���6�i��G[߲E
�\��|i�ː�g��J�Mx��:���a�"Pm�>k��4�-A_Y�ZB�0�$(.v���
»C�D��8~%@��@<����;�SȻ�[�R\�צ�_IZ$zV�'���Җ���"��@�%�r��	z��:�%3�g��`=T� ��{��<FY�m�.�����ỽ+$�L}{pc$�6EIբ������QR[Mx��~��i��Dg`^"d�jآp���p��|E`��</�d�Vk��{T[�{زj�3�,�3х!�Mн�d�Ӈg�]��K���t��\7��o f�U�vg*vw�8�PV&�П���O�O����g�"�!9:�DH�����\�4Bk��n�UE�D��Tm��*�2�eY�Z��qV�������z0��#k�K������B��"�������-�}�6��,��Iq���,��ML�v!�cF�b���x��lȠL#R��P=��@o��F�I��>g��h0�X���ɜ7 �e�֪LY�,���=���/�i�L/���i���˃����^2ZERz�£���7�2`ȪRb]��J-J`��a�0I �l��-bz�G\.ϐC����0"/0v�R���+�경o��b�EuVTyD�-��m�L_�{�[!t9�Z��Ή��Be�3L�3��0�0����"-c�`9����`���i1a?�TO����̫�;�5�1-c���;�/Cl�NW����� ���V-�C�M�S�i�\�i}��u6�˞eR�)��qs��݋i������W��g!�����ǝQ��%�*�x�W�"��$ʎ�ѢM ����!ʕ!�N�Bn9m���?�V���X�E�tFx���f�{�?՘�̶��{�ښ/��#bi*؞q;������ML����^�a���tGE�	��]�ɃA��M
Z���礔��)��C4�I,`�*��a�:x3Q��E_;�c�|�EJ:�kT����5o�l/P���&��v���	�w�Iu�[-�xSu���B2T
hd�6mۀ3D]�r���!����R�:��Y&e���,Q ��Lى3%�#`>���j��,���#ob$�� )���ﮆ.�Ї�z���#�oBP~s�#V�/�9�K�O�%j��;�1w�Y��ki#R-?�4�p�\�X,\%@QNhz��1��D�i7�H���� f"؄�s0(� ���|�l~E�N�,��]�ug�f/wjL<B��s/Pt��	�ա�덯�N�pHD����\*�I�	���V�m�XK�"���w>m��eN-�>b���dS��&NТ%��5�R�9a�Y�j4�x	�(H��7�i�u�W�S'�%K�O,P�ĵ(?%����ۺ�������w=����'�X*;4�\��
����o��-k}4�y ����]����&�Ny_�D�]C�W�p�?o�j]�}��b%�Q�F�D[��T��r�g}�P.��j�:+�@2�&	?L8X*�t�?f�'�Yw5��\?ho�8rp�D� ��s1�lf 3$%Z(������u���h;MJ��J��ߜ�\56%��*ټd����ߍ[�t����=��O�� ݺ2�-� ���F�roM�Qό8��\Gc�2���ͳ��Hvz��H��Z ��k��̶�Q�(�W�y�4Yu�˃
'@vۓ�!2ǻ�Kt�ͨ.���H�I�tos���gv�\�F�g�r�Y��WWǏ,���\YM�B$�m��ݻ_�M.J,.�t�Z��Q�V]4��=�3{�I�  �����&�W������R�1�-)�7RȑK!V�TG|�H�m9���ዶ�"�fd.:�8]d����?��H!��S�dx��kǬD�g�Ε��%5}h�/N��g#���\%Gɢ�	"�^�:,��x�5c;�fR�{�)2QZ0��B��,U#�ttg�	�@��zEq�_�o�	ÅC8qk������w��1'An�_x�ڲ�-\�+	��^,����:����X��.������{7a]g�f�5���c>4:A��d�Cs"S�?Mb��W���h�I���%��J`���HfފJ�ߒ�D��� $h�;<�t˕�;
��>~�ܛFU���j�؛��N�C*��p��/�3���b��[�ԕ"��y�Ď��|�S�)�;���%�d6��wO���(���ڬ��fI���أ�]!����n΄)�Yr�\h>j�<�By�,i��D��XLy�C8�� ٰ��˛����;���+�oaܮӒ����4��yiZ ��e�3����++����fs�Նs�2};�S=+��aK���hVo��s��..9�^����炴E��lJ#� 6���x�5\e���G̋|�Ep��:E��9����X8��Ȧqߌ3�Ր����P�7��R��fPXT�fQ#H���m��Un��D���x�r*��D��D᭵D*.��lm$#�W���ܷh2�)C�Z6�2��e�Q������(On�lAä�\�?!�mO�Q�d ���0dv�g2#=�nH��T^�gG��rԫ���0�}b0m�n��w�Q ;�h�����')�%���0&��w�xR�~e���g]3���his�R�� ��)p�3s������B��	��e�+�rx�H��j�`u�L
�7ص��7����C�R<�7d���1oC��������۲�x��L����ܛ�`��$�-��%���d�#�*П`	7z`�	�a�q|6vJ�e,4���!J�	
ҡ��]�a����e�)Y�z�s�	'�E8@7�7�V��o�`�>��-�׊ �?D��6�3p�"��i���u�o�G3R�R_�}>�E$���Q�فA	w��\��=�~uw�Un>�nN[��P]Ա��6k�������mz�@�����=a Y���H���)C�r���M�?�I�*Su�zF#�]�ێ��k<>�9��{l{<(#�9��@�4] �"�y|�3���Bc�ޥm�(yb�i��:�R�wh^'V���S����"�@;�d%9p�%8^R�%Z�-��	P�~���(���["H5�4Ϩzօq�Go8I #ҍP�ɇ��(�ll��#�����J�>&=;N�6����̘w|>K�E��nDo��H@����S�e[���ʾ���!����~�?ѷ�nU����c&�W����r�bab�_q�|�߂���'���Y�V�bg�_u�H��Ms�ZC�+���eZR��SK�F�Ǐ��B�d���Az����p�DIݢ?�͒�i+1}}�^4�Á�������p6A�V�Z{�%7��.M_�#j��6���ש���\4�Z!K���S�Ew��2C6��֥[�����r����Y��1H���*t�|��]p
'Mn4)6	����B>�c���m���'���tl���ųL���A�
��8�r�m��$�
=wtO��g9@n��6�����&5,7�� �_$�LՅ�X|��� �2N�/��yMG��<��:o5��ȭ�{��\�ka%��ѽlԫ����<	%��$�\sI	�>'��景ͅk?}�%a���7��Wq��j��9�^�;ZL%��)�ET��/#��9��+��8�F_1yY޳�˜x7~�.���(����q`���	)��ZXk_��+-E���㊽7�
�����ݺ(2G�D�i:	�x�s�Le��qy��0Ƽ���C4�������X4(��9�,T4�@�DRzc��n�/N������4 �v(#�{^@��Vթ��ى��rs��@� ;����f�;�&-7������ʹ�8-ݤ�,�'�c)N�h>��Ϡ��Ә��B�%Sj1 ��0Ш�خ�����Ov}��>�z��vnן�G�;Xw�$��k���r�u�v���#��)��o���u%�7�	��˩��O��@5h>P5�����l���1c��jSPICA�ˌ�[\i�V��O�hϵ� )[��s����\Zr(T2-Ԉ�
�	 |�g<�-�݃��0�W��N� ר�eK9�����s^��m�)�{@�v�B�����`q�)�����;< {,,���q����מ�O��j��V��">2Aާ,w��S��xC5(Q'��[�gJ�xRu��4��7����f�%c�&�ᨠ�i�h:b�~8镩a��@�JcG���9G���Z��qvMv�p� Q�b� m^b��f�[�Δ͡"�\�V�Cc(%�1��w�1�\�K�:����=˼���f�3�< &]��YB�;nѾɍjs�ۿ�u�#h��G,r�h_@d��q�b�{!A:�d��:�ѽ���l�^�p����qD�!0��T�N���B�YN���$�_�;�{��+�V1V�1��_}�������X�3�N%�����ʖ�0ҷ>i�8$��]���L���J���@f��&m"L�X ��S�#�{:�Í�@������������HùHʴ|aѧY�M�kx����׈��W���s�%&�s]·Q_�n|��~S�^���sHh6H�Aeȏ�Wd��������Ĵ������Q� �N!Y�[�����HO0��{誑��0$���.O���,�؎Rue��0�AQ�@~��>n��݀��l�
wP[eO��1,�@�M�]t_F���5=�-1����$�ut�\B�b�M�>kb7*,���d���¯]8;m��]��MZkf ���Y��7x��U�l	�>Ђ�8Y�쨫����h%Cxk����b�2',�1�ӳp)iߝ���J�K1���em 8�E:Ns*���z*�f*(�b��fM������jJ���#= K��5�v�5�"�_,����@^��#2��\�����ɫ�=hxީ�L��'sƆ�CS7`l�4�au�3�5�݅F����&: �\�W2M��'�xl�-EH�ꨦƵaN1=^)��C^��t��I����Õ�ҿ)��l��1���p���Yd�/�X-42]UT'=��J��	���;4Wv=�w%��&\��Nd�J�!@Ӟ�7K3T��	�$�c�G��Yp�a�D�q�LoF�:���6��%��"�.d��ٍ#^i�t�������~R'?�ף��w5�Þ�"馒�ߞz�~?B��`	����kw��/���a
�}�trvE�Z�������O�����g�
��i����xU���(�f�1Hu�jI��\˧i��'�W��Q��uLR���#�� �ٹ}�n����Ys��[鷗��yqK}t3����p(ȶ������^{��MSg��>��~//�-�Q�n������
��$609ne���I�)����I��f�:kJ:�����]��xU��UDu[�����b�l��GI"@7Nk1ǽ�["�/��î�%P��T�w���8c�]GK���J�*��	aF,=��cC�T�JQVV_k�(
<9. ��!!:�IQ8gFW-�xg_d4D�ܬ#w��)Ө^	XcfT��9(l�řq"j]���9?N5���D�mӘ�8�U���NX��y15^�i���w��쾭N�����NfP譤��'(I2�g=R�RB��T.k�W�A�� �-^�1�Dˀ%������7�,c}�_�1��5��p\mJwɌ��x���I�e��Y/�Z[
D7߷qZ6(�F��-Հ�����u������Q^����u�饤��2�{&��x��ˮ	e��S�FC=3uC��'�G���gd�W���+t1���7�/P�'�����ͥ��t\�c���jcd7�;�/�jkg���c<R?��K���{���fM�ZO��ӗ�檞t�1L���21l����7���k�e��͍n��ϓ�0��v"T��	�ک� T�?�,�0�ۡ�#K-�c�4�cM(4m��y��5vgL�d~�*�N�nf�m|:h��<ô5�߿��TĂ蔖5�M�(<�J���Z�D�ymh�q�V����>�<F�7DtO����C�[�o�
y��͏�P�xMN� ����Ԑi$9�t�3}���m�X&�8%���&&*�_ǹ��tg$��t�,����x����^���
��(S�U}�m��	]����N��e�����O�_��I,	g��MT�
�#�4�z̈́P!�o�a�5����׃�y[K6�Ы����ѥaJ ����,0d`��@�jmnqE������{�=��@�����={���i�-��9�jt�0��+�T�/��5Ig�-|�a�n5�<[�h��������<ݤ�>� @�<G�k�Vq����4yч��Yr�L�)��i��ZG�HC���Bҩ�an���|�Y��׃K�x��ކ�A*�(��'S;ˆ/��SG�ӭN���u'�����^G$F^X�E�IY�e�R�m���y����[JN�TO�1��9���Hd�h�Nߑ�ԯA(�a�dQ)�ףL���D��ںY��6zy�Z@�N�k��6�T����/�O\���)ť͛����NÃ����*�R|�3՜oUVr4\��T�4������e޳�o�*��'��Y�9����i��>ѥ�<AF�0�Vd�X�m]�H�Ze;M�G���R��W}. `�9����m@Bf���g8�y�ޅ%�l�����������c>��ѻA	�g���n�u���/�s_�s�m� i�OR��`E�r�A��X4��_��,$��¥1pfV���B
 IJ�a;<�U�[3A��5��c�/ya�k�����Hm(d�:w�n��v��˯�o��|9��N�O��=)��Wu��"�j��uyu�z�}�ߊq4ŕ��@�*[8��s4V��Q�a߇"i�xi�˄�YxF���хX����f���n�|�o��J#1�h�~O"��h��]\�|��foZI�����{�5�� &���]���0��k|��������x'�-;����/��h��Y�!�m=}�n 54dx��R�ZN���\F�U|Cu�SӜ��?_�A;�}�Iϊ��׵c['�a�ѭb��6�?ٛY�"	E�	�3�\�>���yFkMI|�B0��\��~���)LF�GIoi�`���)��[�� I3�s(l+P���١�tŕ��X����.s�A�{�zeh%]:���}��}�MR�r���l���i�+=k#��c{@���vٵlB�"�C�D���C,Mפp6�����z�� �0���Å�]��m�-<Ya��Q&�l�?�[[Y\�4���jb����ݭ)!�/'݁�3X��(�	êC����8TUI���!x�`����"\kW���$k;k׳�G�8�>�Xۮo������=Q�D����5��x�f� }���?<��U/��-���|}C�u4�"cY�WzA�ю������`h^_�kk=�Dzs�$eT��Dx��1�	�1��i��9>I�ܦ"�}�l��<���p�pq珯�Y�3ks���:�*�Y6k��n`��Sq|���ߦ���ԗx�:TWH��ī���6IN��W�8�atPyP]�.��b?����h���|V�QP�-c�Z����y�,z�	`��k�7�2?S�	r���f����{�iB�ׂ�7�`qe�z�_o�zt+��="Յ�ktD�2�57H��u�QN��es���%���.����Ӏ��Q��?6��E:keP���j ���/n�.�}��R�u�Z6��V!�<�
�C�u5h����娻kya� ߬�CI�T$<[�}��M�p�ι^P�c���B��`�V|`�a?#@7�X.���m�ٲ��ŧ����P~k=��ǌ�����}9�SQ? ��8�ܓ잦�w�̀�~� ����!|�����,!k�Q��,��G������&߲Χ-.�b�h�{s��s�Tʵy;r�6�k�1*��k}?a��(L1s�Mlάc���B��B��Yr870�O�\xҨGX��z.P�;k����!��t:��C�hvX�|O�N��|�v�w%�Ok��>R�Eض��q��ɀ��]��/IT���*��S�*f�t`Z^��g������{�����+ū1��Wa��}O0FU*h��;�BT������>�޳0��Q�ʚ�x�7�<�+�g��V�G!�Z�4����[e�����������`���(��2���i�9�u�ӇWǸ�ŏ��Z��@�^|�:B<\b�������9�LW�zn��^x���Вl>�0�d�h��r��:�WВ �����U������ >3��
T:{>P�Wu�*���9�`[��g�3��]@ŗ��	���P�UGk���{|��F���;D�v��;j��Ob|���R�C�	���%zbt"�0(����i���.!l�i�e� �x�D�S׫�t:/���FWn� 9�'f\1O^�ɥ���{3�\q8��Ǎ���L�վ�l�굹���p���V�)��4�\��g��q����` Y��s���=��Y�{�u�L11d���){��x��sz���K�A���(�'u���%0��Y�<�m&��;�=���~0��D��nl�ۗ�aBҞ�6��6)VD^�|\ѻ�ŝV�4��3I�,"�\����m��ͤ(J.�,�\=��z]��yo�Փ��|� <Wz�C�_��!��O�c��8��Jo�߳�<Sz�|S���
r�>$8�GA�i��jC��^V�w2�ٮL��V����K`�>�,�����$�n��O�i��
���@�����7�wY�ֻ5���3���_���}p�'����
����w.̜͚U6N,���5��VK6P�H��;yA�q�^��ԅ�b�ɛ�??��.���$��┅�l1�T =�q%����B/��A�>9���
᳅Y�	�#w��.�-�L�����@��7O�����e�0/��C�`���;�P��G����A°,��Ȭ?o;�e��lc?t�"�Q���H0�gQ��
���7ʅ��%V�k[*.�U�� Ǭ�Zf�k۟����	V��f�0��v���^��[W��
���I��-���<p@Ć_�����)�۞�jT��v���\�¨.
��#�,n'���� h�y引�ڊ
�Ű�r���L+->�z�������V��?�HtR����GrkG�@�<�r��o���	\t���	��(�Gz�?�]� D��^l�Y 9����:�I�<bQ"r�~�#��U�L�K��&� <�<��H���c{&<�]�<��|C:�Kl���&��r��d�&���	���{>Б�U�i��m"?����j`�"n}�W��~!*`�h�m��<�ee����J������HH<s#9�w��W@˸�5V�e[������'?�f	&�s����'�W3ti0m��#qض��`�w�`�z���O2{�T�5�.ֳ�:���yFF�҃�6;��V����G*�aG};�~)���͡�M�]\? �����$"*�ZKO
�"��[��N|�'s_�w��X�~��>&�<��Fϕ�O�`��O���\O��g�S��4�6,��󯓍�1;�Ձ���1�j_�&����Y���U38`�%T޶�����FΖi{'	~ �� 寧�ϹW�P�C�i�l��q� ���E5�N����W�TR�F@�[�9�/���[���G����`���}*�3�K��`��7X��A[�_"���I�2��y�G����BҺ���y���N`�Ө�Ĳti����߾�(�'���y�3�a��{�$��@�OU��[�/��]m�ap�2�lm�4��3Z���/�q�&Xvl)��Kkw������;�r�}˵���r� �]U���R�=4F�����L�!�D5�L�b���"��A�M-� ��P%���k]i�gJ���;,GT';I{L
[�F��oM�]I.t��7�
�7 OU܃���c���{�gҾ���!�PVOl+���ES9����`�0��/�\���eYB_�0�?����]��?�MV��_����7���VI���&@���oz�M��D�Ү�R?� ��Vb~�M��7�!��i#�cq>hmS��!����.&&�$P"�<n@�;V�x;�}7�aP��5���}�M�?5Kf���sLV��C�)q�y	@�#Trp	�b�mO�/Az�Y1����O
�Qn��x*�M���\�t�Z��'eX�۽`�vT�>�w5g"=�������>�NS���NI�P�!X&,�����E�P�y��[��~�K��>���V�6֐>������T7������}��s3�"A
��	|���qAɘ܏���(���6�]�2�l#����"�����p���� O��t�������������RW�k��5h�x#ÞU�z<�r|�ͱ���*��ࠔ�6y��2�sÿ�нG:7���iר�##U�:���\l�8��3n��l�R�oɢ]y�cyq2G�W�n�K�L�G!y�`���:�e)*}4������Cg �ҏ^1�����4��z��[����AsQj�ߌd�hY�)VZ#W�>��}GT��:��Ҫ���t�Ө��bb���[���?D����S%�T�i�/�H�	L�NN����_�V3����.o��s��j����7�TW��vM��-2|y:�Q9Ъ1��n��0�!!�f��+�7�W��g6Wy�����pg�1[iH�u��='	YRv�N�8�,��쏞�YbryH,Q T�ZV����0�	�`!=x	�͕��+Q'�_���Q*n!;Y�+�#�����h��`�/��^ћ�Ww<��nB�4�Q��<�z�ch|�O��É�nS�$.K�Vs(! s���|�w�{(��u�ydU�5�;M��|�
�`�c[�B��:���Hh��Pt؞�}��F�����`���ĺ&�1�D��,�.��/��b�{� 3&X�'�>82���Lgc!����+u(U}���v�責h31���]n� T��-�S8fuE�;3V�����jkE�ʡ_�L�e[�\��"N����u���"G�]�������:��YP�~�+b!�NDs�28q�һ�j��T\~g\���&�m����,S��@�5�A������F�Y�ʙ�h"dύ1�����*����R�m��L��{g�w�e	s~�n���=um\~no��^cv�X�V�R^�!�5��dA7@ڋ�R~�Oڥ���Û�/�'�f�u���G��w$� �[��q����ۭ�V��C�,��У���U1,�)�C$op)>�?ᰕ(�o�p���Ibo�o�n&>!J�!�	������2�������#+�=�ǂ�Ơ��������?�:��b�Ī��R��U�d�ѱJ��fr����6�RDL��1طs��[5���Y|�sF�y���� _�_��
��O\��8���@��|D6�}E~j�%f��LߔJrƚa4ܘ�aޗ?F5,��=�����%_�m��c�t(!C<�|��R����1d�����/�c{���77XM�tb�a��/V���Ɣp=e���Tn�L�%�D�t��,⹵����Q����q;��}W�NCGC1|�1[&t�?��l�x���Fsg�4=_�Ӥ\Ef�p���T�-ۊ��r���yZP��DP������vĻ�a��O�`�i�ሾ+�z����Ln"��,�m8�&�A�=Z�A�����c���(|ai�Q�ʴ��4��qg�p}��+��{����NYKz�|Uô�q���<MwuL�R���Ej�ķ:�E,���ŶSs/l������&��+�����f�[GA"��$R�U_F'hƞ����T�Mi�r/V��{��ldd�xC��&�ǟ�I����^t� {B`��ba�D3�D�f����	�쓫�-7�V )O{.yNyyn��-�:�"!���j��_S_�Wui�@Ǘ��J���#��1d`�dy�i*]�}+�D�^�P�n���?��S�s3Ys |�����H/S��8r�z2�#:.�8���82�gW�ٿ�/c\�xF��2�O��m]��� �lO��z�'.f<H-\7��y��4/߃w��F���;TK6�U���+���%V�?
���:�3" "xOum���a�O�{D��,F�Z�v���.�p��"�Ba��[�8.�G�!����:��l�����D�"t�Tǅ��P�a���1+p��jYA�e�l�]�p=ǯm�b�����r2���;e��Zl�s`�ÎCCy��> {`�V����ƂC���w+QVp�w1	�����w��t�0I����\��d�o,tP@E���q��
��
�73q-x6ZB}�F��0��"�=Il���Cv�'�h��T������F�'u�:�%��(�n��B("!%��U�` Q�x�$��iw�ȌwT�aG͓w4JQw��w�	����Qn� ����\<����_���L����u�U��]p��;6�k㢋*������0��S��>;D��ya��lP�}Dc���aB�v�|�q�tH�s�����2� s��p��5�ե?A1���i<(ZGU�0"R��FY_�� ���@���\�qiz�}0�E	]��kx���qԻԙ/�2�����VB��2����`��>H2Ih��L\}P�}���#50غ�����U�H|Iȣ�ޛ��yGN@手K6�����EW1��0��K�i\<�!_k�M��^S�&\I'W�1�������ۅ$ʎW�xT�:���x��P����줿��nrj-��p!����ےeI%/�CU���o�"Ȝ�-Q��Y���Ǘ)l'�
!�X1�q�Z��=�o�<׆*���h4WV�m�o�[�
#��=�ҹ%~̿��P!SaY%!ŠjOO)����|����80���Ԓv�(A���t���U�ӄ�Jp�of��ْ�3���J���d���3'��5�ު 6�׉s��0���<BF��Uc�����׬!�٢�+��
ѳ���ș�v�./N��8̱�J�Y� =�Y�/���K���Y�h}\l����М��s.y������炜b7n��)��am��"1g�0�gi��4��De0)�/|�in앇���E �x!�e~�#��UV�n���Ox�ޮ8�Z���%1(��u`�G��:,nF�������2�6屲;�x��w��AY���Ma2�y6�jJ��F��q(`�n�V���(����=�i����6���q*�)?�X�~�����Ap�n��a���$É�%4T��[�&X2g�W��:{@�����f�'�T��#0�M�q!g�9��7|>�����������������aj�xLn��n�)q
�1LHҼ�b'�N)|��;.��|�x�s^��؀�y0;8�n���*��=p4��?�|y��,pH{O�󃠌�һ��351�C�� 5԰�9U��,\���b�g�����X���������Ճ+7��gm����E����P�,a@�L�C�˔�$`AL�xU����|����n�Z���5R���F&NIa��]C���r�^��X���tb��s�QX�J���H2�wY�P���O��6��iɶ����d�mSb���XYqA��:������}�E�ӸQS9֊�uY?�wn,r]R�۳��F��s ����L���I�8:	�`��]�gZ珉!l����"���"yr}�f�^�y:��ҀQh����kt�����7�삄������h��e�I�w9oK_e.�i�e�����*�H�M�V�n�\`���SiF:Ww�.�[c�B�JS̗+&e��qB��6TC9t�k2f�e�>����t�2�T�t��2��7"�K4��Q�V� �����XA1�.�J�#�S6��6�����J ���򸂊�"*���31dB{p���Ț�}�(9n��R�M��jܽH���k����TB}�X`�ܨ���۳~�`�2����lV�F��?�Ѳ$)�o/���y�QM�L��d����LzȏX:U:��bwF�fK�����������r�C�����0�+C���|R��j��m+%\?"��N ƕ�-{T�� n�p��Mӧ�9z� s[�El2=��u������\_�Y+�_*>fB��~��5��_CR�=O�Ә�p�3�pC�Z2��/o�"����{�<�tAE���Se�w�����c��k�+m��1  =ۘ8UEi�f�6�@��8�W݊�7v���,ɣ�+��N=�/c軾���!?�+���������ke�]1�}z�W27q
��Νʙ��������,Gx�q"��\6)2$���э�@!cr�h���'�\SЇ"���'��;b�م�D�d��8aj���-3(��̐�Q�y����L��3��V%i#D�H�4�����e�ܻ�����J��Jf2�~����?�$(�+5J�
��p��.���Ҡfɓ1�����6k|��_B�*����� �hs{�U�t��i��7��y�CZ�A�_'l
�XiY�.w_��Zk���;�~{�ȷK4�_0`O�ǬV!n�A����٦��_��	~�g�;溺c�u-a-��)��e��3~</n�[�Cg,��1	�r�Lv�t(�����ϭ��x�j�~d�7�����4����66��_/��X�3F���y��b�&�2�+�~�
c�6QF���`'�d�N�����Ɯ+�C n����,6���1�hΐ�e�@�	�`��h�JK��_e�]C��S�M!s���2t���@VPH�jH#��A���do����*��:XR��&	��}��[2���(}�ў{z>����g��_�$�A]0��%mj~w�	]� ���� ��n�E^`������n���_����-���zvTBt Q�R�R�:��'���2]���>�v� g�(&¯�{085v��Q3vк��׌�������˗��;Ķ��4_n�R&�:��I���px��35.�Iu*x�!)��j.KS�-F� �"��p�Oh�z�,��jZ�&P��Se���a	��/q��F�L��!nU��t��aD�ǻI�T�xz`2�M��ƭ6�����Ѯ��c�����	b�$z�Nk�Fŭ����О���<�Q1q�ֵ�6n�fS%5ʥqjo�
q�[[�eN��Ju6�K�Q��)ְd����S�)����i3�"=�l����'3oհ��>~�[k�Շ��%^Ar9�1�(/rt�]31��tI��Bm�g�Arnn���]f�,����f���q�l��	SK�i����̖�՝3P�*|@�g�c��~+��ҭ�
83�]3[��aZ�0�~qb��<ؿ�d��a�H̥y��������"��8���AG��80b�����o� �]`��;�@s.	zJ�"�[;v7����/O� ��'q�~`�!x5�Ge
�ík�Sz�&ojF�^Q#$�t��31�X|�ᩡ��潙���b�������!%$��X4BU�*�TlFgsK�X|Hj�;�/���x�b���`r������SD!�fc}[s�YYA�I���2Z�J�e���7�8>l��+D,��(��Ծ��C�꒖���.�b�������P9XZcŜ�X.:��n�H��0� U�`��QX�@���ڡ��]�������9F��f�Q$��09�s���HP�����liԄ�)��@z�����O�	�u��^z8�O߃�ٷ��+���ϒ���z\H�2<͡0��x��&�\�#�����m����_캑��T��R�c�4V#���%}�ޥ�V~XX�(�I~Ѵ�8��*^:L�8:'i�>��J ��n.�ϟ~���u:Y�I������_���)� l�m]�;uVh�'����>0ܥ,�Ѯ��{�l��<�$��iv��ԀdP�7��l�G�-_���-)���Ah�#��>_c)�tV���潾�@EF���G(#"���G��2����Ҍq��n��t6�;��7���7x�˚�e�<xǐ��ն�r�����ѮrG^q��wn����K��91��^��!J1��=����ӭ�0�3ߘb\g�����Uk����f��h=��#5�WFLX�w����#[:Zf��帾��S� �y�c���uH;4�H�b�gr�$�@3�)V�� �@x��<�E�zP��Y @�[ܕ���yZ'���)�NJ��:~4����N�L����<�j�lK�XP���.no�r����N O���'9�����)?as��?d��[4h����u�ے�ygR��h=������] +�
�T��Kab%Þ�ի�m�1N�����Y;G�d�Ol�f$�>�Ad���&�R\+���4�n��Pb���%m�u&Kl{?P�+I��jh�Y�l�/>o�>�8��/	�16�N���i�6��xk17��/�K\��3#|J}Yz(���c����t�A�f�Q9���!d�T��jJt1�}�
�@ڜ�'�0�j��0�a��L�c?�g��"o��Vv?sy����!_C�A|�NJ>�����,��������5��������hN��BPY�uT�ф��gt�c
����Ӈ]����P��'H�
|����ۤL���#	 fS��v��k�`�	�0D�[�2�W����b��`"'|@q�f�3Z���@
�Χ)I��AV$�s��og�j��؀��I�~�c\�K�CV�J"8�}Y��HU�ݜ%35��g�3B���w��h�=�n*l�Sj���q���[���,�32���âĖ�Z�Sd�*Z�0�<h��9Z�նV��s���-�E�jj�[��c=�z����%7��N��Mz��=��;�a�fu�"+��s���.����	l;+n�,#^Z�Z#�:��R��P��s.�5�՛�S��T��K�C�~��ڞ��#��	 �F��Y��\��mC����A��u��
����ż�W`�?�"W�L�ri�BTv�ߜ/�7*�n�1�ʍa!p���9�>䘯�7Cf�}�%��y�ZKw�B���a�Ԍ�W��Li�Kq�d����l��=Z�3�B���"���jdc5�!^_����O�P1��BDy�<N��G͐\��,��şoj��;�80���1}og�RG�.[,��b��S�;��6C������9
87)���W����*;��s#k�!���x��)5c��F���Sf�6�~������{�fN{>���c{�H)ww\\4������<KVΣg���j����K�>]}�����5���-!�4g� �"�W�����s��sN�S2�-#\T7�wC���lI�;\��"K�#ۼ��q�"�gQ���o 7X��`��!�ڭ��/C�ZweN+x1<��:Q�%xI#�R`@�3�q�9Rm��ܴQ���{�Y�w��o��n��f������Ms�j�k�-�MXҼ�[�����X��0�ٚ�T��O�?��J�1���0`�M���m������Kcx�Pe�k�'	[���7���ް��8��ZP������pvM���J0�3����`�ȿ����}O�&_������-�J:�~t������K�7&��\������,t�����m�8X?�7�`��A�.��X���eK�^ݯ)�:_g�ܠ<P���5�� ���x���[�%#���#';R�+y����5x���M��Z����-� {�&LB,X��Fdq8�U��Fד�<\�)>]�% �k�� ������w����$밸28��5L7���W�]��y�/&u���ë]��7_Y�6q��mޭ�F "�,��n���^rr���ұ`�Ń4��j]�MàJ$�(�x�5h���:k{��/gAt�F'�p��NH�4Pl삃4S2s9��9[��y�\��x����.�L��^Pݯ\e��-�����]���ϛE?Ͱ���n�'���T��	 �ff_���l�o�r�ٮ���B�ֱ/g8g-����F����4��A;��k�\��ш����+��6��K��伿�o{}.V�"�+�G��p�?�wm�N�	�i��D����C��{yW'il2q��v�I�`�c.t���Ӗo.�*�c�#�0��)�N�Aʈ)�
�a��-+���,:�4�OP�?�������~�_�1�B)�3�������ږ3�� �us���[�r���J��T`�RE��V���-�@0M��(`u�x��PAײST�a��z6�+4!�/f�.�`�N�=;ɳ��t�������;��kn���]��p~-ŠM�gަ¡��ݬB/y�@�JC0m ^	2h�[�r]�ŀ�U����2Y�s '��h��߱�pM���:g6�^�6?��9+n��S�_����ŗ����0sH<<f}�	�R�I�A��e)���Pvjh�;�j�Plj�!%업A;�0d��lE؛ɟ�UI�B�=��Ob9e��]� r��Oy���Xb%c̩!�΀�����Ƿ�1kµ���7�;K�x{�x3j/7�M� J���B�o	z�'�Q�&�mr�2��*�	|����gclP"����*��@��_�	�(p-Sɴk�X$�@��֮�[�9h�^*W��{컈��� t*v���c����̳)�>�$�ɥue�$>�8Z�[<_�gvZ��W�a �=��#_d�D׊Fz|\P�Adk��I�,�~�	�`ܭ����e�͒>����H�!	Ž�
�w�<���s,�i����K���T�D[�N3��s�@���`�>Ȋ�7� �nB�ߋ��Y�Y�|�>~P�!��ú�?�.��()�Tݘ�F�
��1�u��V�4v6��j.�.��|����<S�q�ۮи�Z��3�\�1k�9�@����fSA):J|*F��qO���H�j�,��Qd��cl�0��F$�ט1�M7#X �-��.9$�Y'����3 �Z�p�iz������/��� n��,`>�PVË��'��x�����#Ѫm���)� ��,	����O�Lĺh���k�4F�w�|e+u�f�b�.�b��o6ƥ�N�8����E� �5ÁմP�g��	k����;��O'��lQ��=�;�U�>���LsP���1�5f�;�~;��=zΆ_��A�&$�~Q�3��<k���i/�e�����t�\�p�#��uWs���:���+m�#���ޜY��~/��2E�����e�D3!1��~;���z��\C���p���iU��M��|b'[��|r3=	JV	6�:}�D�mE�U��(H�{����Dpm0�Y|ZO�B�ӛ�ha3��ji�I�è�����{X0�ǭ�:,�Mu
x����k>�fi�O��uv��6�s�/'R�y~�����Kl��:7�W8�e�M�+��Op��������	3??�V4sAMܳVW�1�Iޏ��SמyO�ϝp��t�&�]��Kߍ�"��*�9G��Ű��h�\���������p���'
�-���qg��N��Q8�nx�p���!DE$�T��#���A���~���I�z�`����?��5��7�c�f]mޘFP�»y�Y4�-�m�!��v}���np4](BmW.@���F�P\�j�TK,��,W�>�����b܍��������	]GB�eTn*�v~�x�?nw?���T67�0���OKg1�-
�v��,cn)�ܡ���*����r����&H�������$�Y ꣦��L��U|UMͧ��1��A[9$�3�b����oc{���4[`O�2C�@�.k�2I�;9�?#���o /_��W��iI�ϲIM��1w�����s�ͧv�MT݌�z�$�"H�cҹ�F<��ޡQMz3[̝M�������C����6����q��:��"5�y���H�(���w�4l���,�-�٨z�}\v�j��x����Z\� �ަ�:����%�Gw�l��`�#�V���Mx�������:	��Ii�߿=n�]��%�?ޤ��s��)y���B$������e����@OFXHH�#�p�����Sim�-����S�#N���b�Н���
�o9T�_Ǹ�=л��Ұ�w,��!��Ơ��i\�!�.e���C�����4�v�9="�qwɵ~*=}����Q�<�XD#��p�cڿ0��W�'F���}2Q�Oi����ăpf�4�..U�D�y�ӓ
B��r�����>���/��Rc��7T��ObL�j[DA�Į�����}�W���99��ha+<�'���:K{�զ�C;���c8}��8,�W�Q8an��A�z�U�����o��G��z,���Wk��hNTf�`Oms�2b�ئ�t��ň;XiL��������7��'1�C ���~hNp��d�e��_55����M5Nu��r�7:yDPK�0o�� :�46Q�0�c��}���F���$��LF|O���7gC2:6
�%&���}k��Fz����zF||K�3g�<�O�m�Ο� W�́:�Ye:�tL%Z 5�(�d4����
W뎒{"61�h���4���!�������T��wO׉������'�Fw3hi��-�_a�b��N(�x�]e�"�ഭ$+�O�+9��{�w�d) ��\�d��y�f��y*����@Ͻ�b~�<��(2i��p�y������� ���`��5嬪Q�Ǥiǹ᧐��92�/���IMr�����^��~���<^��'�Ts��N�*�Y2�'����b`��������b��3K@~���T �U#��G�H:A�z�5��t,��\��
쩞�	Eg�.L�'���mjr���n��fW���56�e�ʴd�?�A5�yv�`D9��E�Ś.l��|��.;�[��n�R]-�J;ų#�}Q�	����*�m�3R��g#_��a��Z�sF���t��Ҥ<U��S�m����h�����h˞�c����7����A��G��gA�n�P�����)zǵ'eL��y�ކ������y �^�߃�`(�<rx���"ZM��<�ϮGؼ[�x6��yێg����T������[�7e�	��QZ�eu� �XI�Sb�9@o���E'7�����|�^r�"_?*���ї֎Q9�t='�����gHK�r�SK1"@HP��~�*d"��6	l�m�x�f��;y����`�5w�������Մ�tQ��P_�3d���tn�>���29X'x?i�np�.� $��sE8�q��Fa�PZ��#h�Z�/�X���������E*� H�9� �����&^^�N��Ky{��XQ*�����Ve� I�ϔ��x�SJVd�7��A�c,ȃ�p�i����A�U08r�,A�T�B�� #�aO>�Ϊs΍}t|���Q������SF#?H%������%��s���P��4�z���2b��/����0�j?^�/^Y��7b�3r$�4h��FhNgl���Y_+ݕ6�?��lM*;��<�!>5O��Eo��<h�bL�l�2P�(��#���A�.�x|�P�H��!-�vc�SO:>"soM�?�$	�@L����H6�g�k�e��zz�%P�������&�?� �&��v`2>�����+x2��l@j�t�ȾI��s=�s��x��� 'h�6�l��B�0����A�{C�6�=�!��-�ȡ.��2m\��꺒����v-D6^�\.[P/Ԑ	T���|~WgLu�`�'�R4�)J`�i"A iO�Ke��_�,e@̜ңD��#���zv�����ּ~�֑�#���衤Ohq�=go1�xK�����HM�c�Rd�E<��F�3�31�O�=��ETřI�7
W��	M&[Ӕҁ�ܘJ���9��=���n�u�^�M���C^��*у��h�2t��f��:�O��rcf���0���9��֕a������8R�GUM�B�9B1τM,�����܉�T�D�?��m�װ-��,?EU���	���Lg4��!��W��;�x��E$CqX�N�#,�}��s�P�W�7���	F�Z��.�*^mZ�`�$Ӷ�L�U��*x>?J���)�ē���Џm��f*q|e�&�v*sx5�栰1G������7���hQ�1��~8�8���U���u�a�g�p�����2f���\t���������Z��CYՋ���v!0�7V�(�y���;�������y��I�n��I��
i�xYK���x���ж�B}���xp !"��B������B3�����A���f ��"�}G�nU9@0t�Ot[R��u�d���&*V���瀎�!^������
� �9�fW����!�D�nc91�u^k3?. ��o��Q�[�����f]�Y�.�ZH��7�'�5��X������T�.ធ�TbyٟM�)�8�A�8Rwa/[t�9B�ۊ��� `������������X��ݲ�H��|�
HM�Ȏo��o��k(��H(�Ɠ*��h��2
ћWrF$��/����t�@CJ-�y�š���_!iP<Z�1I��V�;W�����>~�Ǥ��BoN4��
|�W�/HT`��_Q<���5!_q�:#�0o������^g,��B5�Z���4/�c;B�ӟ1�e_�)� �0R1�P����m>�����,�=��m�vLF�wص[�6�*�u���.g�Ǣ���)}q���:��OI�H�&�u���@�-��"\@˾�lM�gF�4�_��z�g��ZE��5}1�r�9��3��U������Zx����9�`7s��^dJ,�4f]%����\�*t��>j��p1�A���t��f���t���Z��a 5
�dd����]����P��z�C�éK|�3���.=�K�AN%�����k�#KI��O[E���� 0����>�"��feΠ�O�@"\���88M���Q����a��zI�e�u41��{���S���1%��
ɻu���c�'h�<+�_��E���߷�ѓ�pJ��7@q"#�|�_#����w[� p�vZ�^�v�Cn:hKzԞ��ߎ�XV���D>�Rl��q�`W�^<��"/6��3�(��oNm��B�9�aL�f�5���
Z��:S��~.en�VX$����k�],�,A2�	sm�*E�8�\���{��x�L³����&���s�{��lꟵ����NXL0P�{� V�e�wȾz�e�{�l��u�I{���5���ѩ�� ��ů��c�C�r�d��iJ�>���o�-�˱�ߦF�v����un�����v��KHd�F�ʱxvC��(a�f��O��ZJ��'�ʞ(�n)-��&�T���k]�l�a�4W���B�s�PC���up��3�U
m�=�1��p��> Aҋ!e���C��G��lT D����J~O�M���5��}N��"@|󋵎���5�P���� ��|�X>���!� 9 �\8�VN��{��N.�� t�9b��>|�z����oH��F���ۂ
�:���-�{B�+|6�'kaxOg���Q��
ޥo�r8���p��1�Ix�8�&�[&��If� ������c8"|18��ߔ����;�uܝV�`�;ii㈩hep~�Ȋ���<q���$�����On��p����������Zyrd/�e�A��'�,R|�D�'J����VZ���Qw;�rН F�( ���Q�5��}p�vվ�����l�n �.&7�UL�"�V=�@��J�ӚjJ��&�j3�1T��F����#�@V�-+N5v��1���%)Yf��O�8[ST�I���3
�1�q�e��='��t��cOԥ�¹a��-FQ*��i�:�𱖴� �-���u\`+-��۲�Wϰ:+��U�������3���uX&=�l�����{&���I������|�a��-;X�� "�����u 7�d,:c�a;�� D�@�	���y��L�с����
���|�V�6��%n�p4�~C�F5�����S[ ^�'�~+��3��EcL:7R{O����)��Q�0\>��K�q)��:������Ĉ���ꂆ��Gl�[I+��^#v� �Ɋoi/u�kd�ЄȶB�q�L>�mnx0��!=.T^�T<��-�8�̷�W<�ը�v�s�NzU���)rp���w��\E��3?���n�l�2־�rW���]Lj�P���qt;�MΆ�55�x���c��"X/��R+t۵���nOt$p��XD�y^�6���S�<ʜ�'�j�x�Hu!�BG-
�#�(}:�/V��6=qT�f~�kK�|���Z*��F�!�{*!|?�<9]�PC��:)P	|��p N'�t,��e?�����6��D��{A��K7�_)�50�k�U<���BfGd�K`ԡ�����a �,�}�Mq%_D����y�wG����ɽg<=(yJ8��*�q{�x�O$ؕ��p,:��1E�,����4����xFQ�����)���R�BJ�'Dݱ8Ʀ�1���_�n��;)l�j+��Q��UPk�����A��qW^���V&�P!�ef1(�C�4��pdWʀ<��6��xyU|��ا�~78ceLme?��A2��	�L�Dk�q*����vUBe0T�{Z�V�#�b���Y�� @RA��d�˂�L���X<II;Tg��B=��%(l��yc�z-߁�
�UFU4�<(�e�,p=*�8�����2]7����sH�=���I�j63TJ��O�t���4@��,��2����2�Y�ǰoI6^�4-��k'"��$9 8����W�P��O�y�e�?��	��K��Kɇ:f�@��ɝ���R<�����o���j��"ή,Y�F��/��+嚓^�ina㟮D��1*��,B�Q;�`�o� 2�KH>��.��ĸ�A֣u�"�TY��{ھ���a���{����X*�=�5��&*�ۗ|\����c�4P0s����O��t]F�U�H)�?���ԝ�v6g��C�&,3�e���s�MU�����E�����Si�R���O�>���'z��4�U˘��A�	5�6�wjV_o�H�g��g#��&���ͣ�[��s��~���}�������f$H�r@�|�ϛ�*�|٨o�i�<.���A!^c4z{X��>�B�\*��&����	�����F���O7�����~c�u��;��Vw�E� �a�P�w%j���\�}��SdPMKʚ�y8o~��:�׍��X����� ��.�í�vr�����d8�'u:7�>����u����偙�K(��0ⱌ�Y��Y��NW9S��W�[�BR�B�VU�lSF�Xe� {~�ɮ�`r�:}�9�X��[ ���P���@������úE�I��H���t�Lռ�ށ)����`�yY�K �AZ�犻�?�F�_x�)^[��a��){}�N��Y��ޥ͋�LVF�(^Rj��Z�x���/� �XG*hN���������UÔC�
���}n���J�o4k5ۢ��~�nN|R>B.k�|>k���g�^85����ǵ,j�p8��:������eFh�Ҫ�{�u�r
�2u�dL�X���s+d��m�˲7O�:�w���w�r?�=�Fdqrd����vuj�B�V��r��3yT��I��Q�j
���nGP
9:��F�� ��f}}p]��Uݹ�.?�^���[���zBS�P���vP��e�9>��gwU.XCI�|�Cxǚ�P �%�W�C�����I��{�C�=8��K3����Ǚ�!&㎯/���֯�~,,��|j�ٍ��������3�����`�̳L`�xa"����=P-M�j�x��*6��c1ɖ��x���8�EٛQۑn��6)l��I�_�Z���W������]7��Փ?�����YB�k%�<��l�f��-���#�E��T�|o�~�ǉ`�ΆH{�,l.,��F���ŕ?Q{��].x���dfJ��l�m�ќ!T�//�ʻ�3̐B�)3zC5���}{��d����LP������θ�v-mVnjL�բ���|I|Q�ː�y.:�4��M���8]�[u�D����I2�~��?�uI��qŖ�� �ꎈ�³��Z�"�[�����b�w{+��b��A�&��6_��(���O;��[:���'�� ]�+�hq�rG�Y�7V���l�� fw�6����,�uΔ�$�N.�uGC�U�ui���|�x�.�,*N��k�(�ҕ%�w�l����)�Q�8�����t�?\���`!SP[����N��=p��\����d���-�m�7��Omډm���)�K2pB$�:�|��"�m��/Wb�N����&�!L���o����v:�3��?0zk��;f���0��.�1����QIU"�j�3S�܊BS�7�cu� /�= *ߙsէ��L��9F�dU�N0��4,�?�b���>������䔏{F5�9̭��G{���#a��&��A�
��S����!�,a7>tg]��0��&h��'7Ͽx�v��U?��S���% $(N}S)�k7q^�����Q���2���/)�y���#=9�g1����j�o�0��C0Ri#h<��S�>$��YP��3�J�%,tY��%�O:��у4�9�������bL���Lv��k��ig����eO�g^v*qa�	3f^t\t�Tr�c|��Toa6M��S�d��@�)x\�� O����X4$u��*�gٙ�ty�C^W�5PC�R� �k|�?#����ed�py�	N���"��jA������T\p��9�Zu�D��h���r�!�d�+$��V�R�ӝM"SM�@��Q3+�G�f=M�.��,�c�s�2�(�W�ڰ��ݎf_+����SJ��<)a�_��m�r�!�6iX����N�G��<�wy�)���q���$�t}׳n=~�)��LX�kj��a�B�~x�h$p��}�"��?��Wd�f9B-�j��?���mw�������gȷ#�j�'dՌ��3,�Q���Y��Ў��f�����f�2%�&� �``i�����������{� i��çL��H`5=���В7��Vf�F�j	q}~o���1oGo�4��-�
��	d$��١G���o4o8�3f���!5&��Ƀ�r5�e�(#>��S��M̽뚯/�ð,��c�a˳2_ '&�J�a{�K�u��Cif�['�s4]��ql~noK����H�
�|o;���WlL�;��ܔ�M�m<�u����M}���:4c�R�ͮ���U��E�������GY<�Y@�����b<�ߠGb�Y$�n�-�0��H�xD�s�4A JM���,�r�o�#�r�`0��S���ɏ��Q��"W����l`v�QN��߇��iU�!1�S���$�p9�����n�VY<+���C�\�!��&5+�P�/ʥ�r�4�g~e�6Zn��'RС"��)��>	����.|����#k�i���."'��Z���p�G�u������o�+��pr9wM���0H���Ƚ�y��נ}�im����/�_�:�TߪKT���e���?:1��|�&� ��c��{~hݰ>�	�L7)m�a�FP�������mP@����{Ga>�M��6�����J~嫀��J��f�q�]�:��F�6���K�[� ��Rгʶյ�O?u��Qf�_�H!��޸��1�Bmk���ʜ6�����B����"�)\ YŻ�y_q%��@�#�]Z0��:^�>@�k�:W2��>4��ĞmG8�ق*�T�����a�UkW}�����3�UY�f�l\��ݓ�v�����*6��.z�oF�$z�7�?8��x7���;�!3�����9eA�u����<�e�I���b�8���-���lf��A����L�8������t��M�jq)e�Ҝ��M ��1XeruT+'9�/����:��)&�ظp��g_4�d����ݒr��JB�T&H��OD�\�X��B��v�韙���D�v�ibg<`�߿�����F����$�עu�"�Cr�7���ʚ��}�`��%;ΊL��_Æ&L�V��NR?���W�l[£�
-3T؁��Z��]�J�ُ���٢)�,�$7��d����7�=�2�@%6�Htڎ�i�f���(^<RX���O*&N��wK�u�W����m����[�n`刼 Lz�gm�c� ��X��.}�,���"�+Fh©xJ#�	ln${s�'�u�)�`-�E�7�N����k?!;��������8�n�9���~��@�9�9G�\�8�i�fEd�c������>��Ӊ���֧'ּ,�;fl�� xc|~ǐ-�/�5cȟV����j3�~��̮K����.�Qo7fS�XA�t�8������o�p��g��*\�6md�o �eӡ��GF�~�r{6���0�� ����<&���M��r<"a8�\���pv1�^���3ы����i&P�Y(�D�V!,?AOC�I:Æu��̵���;^Ǥ��E����Z.������ZC�RNG(D��5L���-��27v����=hË�?(�:���Wzs���Y�r('����`�ul'o[y#�OLw=�0�Y�uE�"��n�"ϲ׌���]�� ��X�Ni��,����j�?Pe�����b�8ƍ�:u���DШ�i
@P�{��9������72Ʃ�4>6�N;��Xpr-yB�%��M�9�����������C�{�^L[X?vP�*�{�n����ם���c<��e����#ڇf���% HN��VS��:N���&|ùjl��;�����頒hb;�tҨ��*�ۘ+����~���Ӂ/+N~C�2����ܸ����\}F�ѸpY��>�mM5z�O�
`�+�zk(����2t�w��ܟ�4�bڡ/B9�c�]�+ɨ{�/���q�/��|�Ȭ龰�--�;�9q�⩨�Lr�2��_����B�E��D�pێ�D٩Ԍ�v��IXͽ��.�
n�޻3�&)$eP���嵗lV�_`3��P�ȹ�{��fQ�,�"N"���� ��v��x7.}i��p��׊�����L��j�6F~��G�Թ���pT���j^���Rc0uً�H��|�>�)�tq�E��Mxҙ�i�n����*Q�Y_�F��D\7�_(#�.�#t��	G�o��;�*�!֔,s|1"J �@F�"�B
���(��K]��w�pC�*���wݑy���Dg*}50����w5�!V)L�-?D��~�&M������w�P��e М��؞��.����ݑ#S��t�n�nɪ��E�ρUi����}|k���q��"ʿD�1�����x֪�^i���D����@�n�	��g�����B�������Q�{ϧ�Y^q�/g��n{@�]��	��NwB��a#xM���_f]��V�Z�CE��M�d˸'KJ�12y*3?kTuR��I3�	����9.�f����(�:�ʮEp��X�jG�b���#�O_���S����%
s̤�D�� �"^�pc|ގR���{r,��
�K��Df&>x��Y@vs)t ��r�m<NpYZS��5�t}���Fo [��_>dȚ��L�V��7�L����]�n�!T=OSM� <\f�V�FQ�<0XX�1�=g�O��Ҡ�N�F^�v�e��[u�N {��,�+�,�zf���g(�Q#�h��C�!A<���uY�썋V��]������--D?���V��r�?=�CKL�GcO@?`�?��!I�%���_+��4a3
���Y�f%�T�g!��(s[����-~V���:j_�O�bM\��Q�s�B�>w+Q��S�/��G#�V��kR���nT��ȝw�&� ^��v��Z�����5襁��R�0MA�� ���PA��eg퐴�-ָ�Ö�ލ��W�����d]�(�!1��(
^<җ�����I�3��uA�!z�T��D��	J�,䍦9�����_��8�V��I�D<0��+�����H[!y�W4�(���sBC��O
>��M�В">5C�IO��[h~g�B9��R�0D$���f�zI�80ۿ��O���-]�6�tn��ƨ����F,,<~4��\���Ԓ�z�תK��ea�A�*�=�N\Ǥb��-��I�C&�K]+��n��B�A��* ��Ⱥ���g�E��S^Ա�aos�B���ʨIi7�.������K�Yd�'!�sbɟw �ݕF��3!D�%j���lC}��	Q�4���ߠ|"
�X�Mpu���]��(����
>0�������Q���/��W�S1�䣅5_�&'7�[O��V |�ҟ:$�:�t����`f��7;V��ڤ0 f(V
O��9�\����Af���٦����
��M.����p�G��.%�g
��O�O:���#��3ܗR��?� �_	$��O뫤��h�D����06d0y=~<�uJ�MzP�fR�,�~��:�L]\�NޣUK�5��C,ߌ�����; 9�?ĦDY�}������m�w��~��0�9��d�Z�ޜŃQ&��Ke�����Q̀U��MXR�#.d>R�Qӧ59�u`��\L�4�;7փ�;=\2��U�$��Qg%���[���XVts�/�B�q�ΨY���Hj��l�6^ľ�'��2���N��E���媉�������+�0qsk���,�����3���3���n�1e�6?++��I�N��(�ցՌ�C֯/�Dn����R���Ӫ�J�$3��:�8w0�&Q=S$��\QW�;�4�AF�e��J��Y�n�mj���m)���X5.�Ϲ���Q�� t�nt�O	�_b�6����K�K1.{Z{�*1��L:�8R��"p�[��Q͈���֜Q=�TS����E��3\W��ά7�8&��S�V7v��K��y��a���������H��SJ���s3�wI�|i�X��`��8Ɏ�I8���
��8�K`���A�)������\�@��x���C!&��p�>1��Y���,����h��ߩ���İ���B$:G���"��pK�Z���=�PZ9h���k1���l�)� �'��W1?;ϊ��:��=WY~��m)AԆ�e�hҪ ���)�$�z�iv\S ����0����/db:��h0�Ai�pјH��Q�#mLTBg�2��m��n����_���hi�j-m6&���+�jxQ⅄đ�ݫ� �r��t�A�z��KJ�����\-�0�p��j��(����&�R�M����*���D�y{�W_���z�Hq䞳&�-o��F������
ʻ�If��+3�+��D���m.y�-���.��X��\�9��)/n��}G$J�1��5��.ÉO�	�j��%�1av��\^�h�On��1�2^C[���0<z������o#��/�ym�(\uOK�Y�'沵�آ
�p��6�NYNl�5,U�4%��{F��s$p5����)s���q�ӧ
��R(�É�/o���8��T*���\~�b^3��*T���|��� ='��w���:s��.R�@��BMuV?�ꣴo]5I��05̈ �<�M2n�ᢨ��� 7L�gl�_1���"���n�[C���8-]q��>�Qk���Ma�x�^AR�����w���I�jC8՝���3e�u�p�����[&C6SL�31p�C;]4�8p���8;I�����X����i���M%�7闬�cR�t�Dtfiؔ3��k1фRN��D�k �ߵ�A��;����O�'k��[�Ϻ6�zg�W��i���_)U�;/����Q��*�QK�%�ˡ6��j�~A�����
V���Z��:��b+�WvȰ��w.�#�g0���g���]�þ ��8�jȦA��{�,N�-{�[�O�f�D������T�{��R+��/mr�\}OG�%����}��`F��
�'��?�_hC�F߻�B����������K
?��\�"ۡ⧵r��@T�v?����&�B>>���_Pp	jCө�_�����I�MrrE�~��ſC;��岜4��k;�p|�{O�����[�UZ���l�.c���E������a��w	6�zQ)�9�rT!��v�"m,8%�|��3EQ痎�^U)�]�x���n&����U�'��.ϕwYm�i« ~ܛ8�k�fsV�D�czӷW���g���"���}���ނ���w��_�g�5 ����k�h��� (�ʵ�sk��/�QF���/�aH��Zmf?�@�p��UP g�;����>���3���z]>򈒠�1`n�$5F.;ڷ�ܸS4[K�"��!$[k-���l�f�IYI�@�`�d$�֤d������5�v��9w�^ �o���xe��u��.�ʤ���"�
䣄7��r�N�Y)��wf,P\t���BUg��V��w��9PrZ]�za~/���f���d��X��l  ��RC�
�Vd�~�DA�9J�Y������{&P�E����,�\����J��;t84��)�7v&�/ho8�U���wxZ��EiyjK��׮�F�
�%)�"���eR��sl	 ��a�#I;��@7qZ�h���#��ti;aY��A(�Ya��l�u(�x�����W�|e�>$�'e��ӎ�x���._a�N���*S��%�/6fœ�� .#02!�a@���gE�$[��&����2�98��X��NfX���p��:סs�%[wK2`O��$�k���C�Z��e�5��BVȣ#�� ZI�j���px	�	yC�Ύv;��G��J���&�|
$P]��߭��YA�:t|ʆZσ��U�1+�İ�D��	���*�p�N̇�s~�3 ��\,.p�(fg/)}�%�h%Mȶ�u	�ŠJ~��@%�h���Պmx�� �)����C��=�aFcO��HLvR�oԸ�{-��h;D�����$$���0�+�ŕ�j�n=�����J��� �{�gߐ@����g�S`	������ĕl
�9F�asy���.�<����ȶ�S�K?OB�K��l�^�R�Zf���ie�EZ�>$z��z&տ�9�<t�8Ǭ��Ь�	�|{�ȕ�����g́� ���\Hϝ/j���G���3��h�x[l����e\�t�ړ�[| v(L�ڙ�)�%<4|��r᧶���tE��V�cΈD�2�j8���{N8%FnѯK�k'��-�@�V����
�Š����ꃱI����5� ��K�Qm�uY�8l36�x���{��kٱ��Q����w�|@��O��7��]g��8�_�[��/���g�Ӓ.ER�5����j4�M��O����Q}K���D�1��9%;~v4�F����(�g����[�]�ޡˆ;��utI���87�<YEbuaf8�n�Cb!�{A��<�����WB$M� L��f%��c,�I"�r-E�)�[�َ�@���[�~f�K�T��i����xKV.Xm��fp!e_G��s���H��JA�oSN���>߻$����j$eN���_�į.�Lz�<d,Rcm]r�o��o�����\�7N���M��sdџ�"@�й^��1L?U��۪�_�����}6��n�)A��� Un��R���������#ʄ'���"��>�60D�$B8[�>l�ΖQ6�~��kH-���a�ݏ�޵�P"��.�UϢQ�V0ų�%��1.��?3�l���Q�!��Ǻ��=��&č#4�p�\��'qo�C�4��c�8�%��wɧ�2y'��1`��_cK��t�01�P���G4���;ѯ���1�U����c�b�u�
C��N��6�nЂ���H2�	�WQq��]�;�6u�|�DCf���-x�R<��ޫa�C<~���6+��E���/����tW�;���Qf Bx~>RrJ4hX+p ͓���Ev,��+�]����$�[�|�z����c�).�E����x3�"��ݱ����
�M��CC�.�R�ȍ�d��Iճ3�����{�8�t�1H`Un���|�q3�0I��9Y��݃��Q�7���;�u����O�"�S�t��U�Fg|���P�P�Y�G7�F�M�~�2q3�=��{g�����R�����!Ai�
ɗO�6�u��?���=!�!�`��֬��w�C�F������"�RsG���>V
3�_1�̒Զ,�P�iiZp����",��֚�1�
�f�+���`{2'����Z�&8xL)C���o'�j�����JG׺ߣɫHn�5"1��f�ļ s��X��<�e�r�I�ݑ41����@��NF4u��]2ɸ��m��O�f��^����P2�p]��3V�w���� �,?�ht&*���h�H�c��M��,{�=��*B��Ʒ��mf�\9�kf��8�n��|*��2����ڸ���j^)E�1O%�+��t)�i��e��܅����7g��w���+p�"��J�{|�y|�g�]��j�zL!Xj<����Q��IgIO����&$���G�`/6�� p#���jи�g�V3��ꔋT��q��F�����C�}�w��\p=�b�P�`\ ��L��):���v��Ů�w�H�[��v�Vo/�9�����DE�m�)��2@-�����t��A���^/�<~L,)P)&�'�	�/��Il�%V����?JS�'5�4���ٶ}���nF$MP��C��W�������2�Y���B�R=���߯b����$�_tɷ�T�tȄE���8�^]�Ռ�-!x<i��j��*��Lr�_{�d[�<@�LL(Ωg5� �2wJ6�E0[�'"}���wAW�dm��g�%���QV�@��%-�һy?s躲�����J.� hC���p?�И���K���XSq���B1����3�+�I\;�U�}
�� �r�	��vj&fj��ȵ7�3��{\�w�]�#�؄�d>jC�=�^�FIеA�����h	�����%�!#�i!���#'w9 1�� ��H�F| �񛻃T/Vs�p���=5W��U=(4����c��D\ڲ���=,U�_5y�6�V�1=G^{a��uMW������1�K�GXFTo���4&���_��Ū�σ�H)m��0�'ث�a(JM��5��-2�L.a�Ru�gxL���� �>��� �o�"��=��.��p=��LX ~�QV�^]2r�Kn�ֈ�|u�!+_\l�zY���y���bs�{Q�~�ܗ�p�)N�%f]}r,{	��7�`�����Vb�Ml�(����D�]����h��֍,i�}s�~���M��!2{4��߃� �|��j�8�Pp\�ϳ���ۍ��,[�=�>�}�8���
ɘ�>e�,��S�i��/3��f_G�?s}oy�P�Y�I�1G籕���S��1-pɠ�V7�����A.p�s��)���6�N6�h)�L��l1`C%~щ�6Z��M�~£�(��J��n�>Q�m1��;Z�O92�zS����8$u,:�Ɠ �`�Yީ�v���~����;���� w��}%	�J�:kv�����W��	J'k��p)�D3��𜎑M�ѣ�.טqV��Ⱦ���$vǔ��'���8I�:Qtj=�cu��P����u��w�D�?����d�@�6�{��u-��Xp1�wsD��.�#8(�f�@��in�([���2�� -I�Z6&��ÿ��n���[塚�_+%�_���L��3/ɡ�l��� �Y�4k�!���z�D����*&
�o��3o'n��w8_�4�P��q|�:�4�=;3��x6�S�-{d��e%*�Э�z}Z�3i∖� ����6��~��h�py�����H�N�r蝺j����q$�<]�\y^�^�p����o�t(�)iݹ��'�q��N����Jz�J�/�B�U�����,+�fgaE;���͚㼾s0��/�"H����,=�޴a�uy9���еW`�;�!�4�s���O��Pa�<%��fH��D�
U^���|1~o1�؋G�B�� *t���OH���Oupԟ�`Rڗ�,-�.�% �;i+�[��9�@�Oy(&g���B{�$���*�����^6������/b���A]��p*����X�^�J+�\Q�`o�����[a�&��������=�\�[gH��لb��$\4��	ݲ��!��G:�tƠ�;DX���EɌ��/&J�Ԧ�nE��pR�g�Գ�2�b�A�s"��K�G�����߳pQ��1�4�5�0v�"U\T�jN�#5<!��T�YE�'ޓ��jd����*{���I�b��Ч[���B�5������ԯ���"�ei����&@x�Ldq����hq[e�͒�b��I��4׹lME�U�%�������.w;f�Z�_V�fz�IoEx7I������nK�AĽ+uv��'�B�9հHe�R,��nﵛ�+��Z&��ZtU�M�<U�AY�s��#S;y��b��:��	5�I�}q�O��1s�����66�2a[��H��OP0�2���Ð�j�!O�-��Zj-������i����[��n��q�^	B�O��z��
���R��SNlL���C�Aq>��N[���4|� �G�p�7>\�^Z�QDXn�p�p�G����MJ��֮��z�@_qo�`�'�[*Ne�7�p����t���J>s��(-��jҨx�٤o�H��7���:>���ŝ*�b.h����ȍ���z���3sM���|)Mn�8�����D����#�5>0�$
P����oq�R�m�&���T/�;Z�ʱ�e��J����I�3��\�_ ���\��h=G�hi���8�?�Nǲ;���a�u�)������=��g<��� ��iA���V�1������(�ϩsʡ��%��F��k�Sp}�%���\�l�!l�U0�9�X�bA=��Xm�Y9Ĉ8L����+�HV�5*�OI���<3%� ��^����(�9a{Yp��sIV�]Nԇ��>�Fgek��"��2�,$2�a�Q��O^I̅*��Op�X�E����Y$jcF�>���S�b�̢�X���rֶD��`jL�ݹd���⩈�!��⹟rz�k�`�2dw�(Y6�����;���}������3pZC�\��K/�drRX�l\��8��дfm[@��ۥr�
��/3J��$�z�}֜�3����(�vez�50�b'����P��!���9/	X-�Y�MO�b��0������Z�3Q�»���0�w��t�k7u�{K=�N/-5�aXM�/H6�L
9,��`�"�6��A�&�CB�����3A,YB+S�<��:��&y
_A�gp�`�nu	*YxuP7���*0�-�0�2F�/6v�^��wӧU=����2�����	0�{�[�X2 ��%���D%��`IY���s�z+[�ʥ��	�}[i&	Z�Dr�a}�\�E.8���?��ı��#�g�8�_n:G���9[��n�.��-���~R�H�;��_@އN���E�}��o)��&f{��������.�_n�re�>���,�nM��"�D�~,O�yZ)��>!���i[q��������'q�T��Ɣ�c�()C����7M͚�'�.���"C�L�nAG��B?+tA�������ߛ,�9�Cnβ.�0e�K�*�R�]���/���1��݉�&���,2(W6�� �/J���,Ű�'�*5?e�-�����(��T�7[�8~����6CX�&��~;A�a�%4&�W�ϸ�Ǹj�"�W�֕^m_��ݟ�T�"n���<�}PY�M��@ ��9����U����8���3�e3EPd�{Zuq�r�`xN��:��'�o��S��B��tC-�h�@,�$k�UZ���f� T)�5I�~�k� �Gq� �W��}J� b5�����0zG�M�*1��ʉ�]T%����%X
j+:`�.���9�$|�y9�nR�+���h������V�m�I�*��\w!�<)�0��R!��r��O٠�d^�H �J��Ͻ�\����/��R�-�iq��FXP���� +G��$��H�L^A��"��@�Q�ɯ]`������C�u��T%8�7B ��,��r�x+�d�W����θx0Dī��4�|:��&:��g�>�x�F��.F�>m��v�qa��!o��A�L��Jٚ�
���=��lPC���t��G �^�x��X�ԇ,~
�J8��i�:�����T�R����$8��<+v�kZG�� c�b�ũ{����5a̠t�x�s�\�j����~^�,�b~�;�����(l�oYg%JZ�<��-�붆4C�H�S 웑_S���"J_��c��f�O�O؉�2N���i��A�L�~ho@bh_\a��� m�_9i�9��j�J<|���>��$����`�4=�+�Y��+�^�o�!��\����XDN}���d��h�j�~4�Y�%_�/xx(}���.
L����)ӓ�6 nn>��h�p�Imv�B� ����T�؅9���u~��f�)%�*� J���T<�a���i���푖�f��L�����>��wvǖjE9�BL/�1u��k�����n�!q8N(�r������m�rX1x*/�����q�;�H�� ����>���I#�<\�4q3�F�Y�>l$�Xp����hw=2�*(w]2�b��p+`/&���8����f�l ������X�7x�^�YH�T/J�e�A�A���"T�o/��O��@		,���饼k�8����:E`�(�B8H�+�%!�z)�M�P�m��2T��tX���
d\�T����T�?l�����v�4�N��d�{�c��p�Vm��Zl��������v��"���H���"�ɔ	�����"`�� <���!4+�d� ��b��IX��㢩� >6޳]I`N���iƇ�d�y.3�ќ���ۥ(C���	���a�5������ͬ�ߵ)��&.X�9��B!.�����9��I�N�����j[i��B��u�]ՅP t]|u}x�X9�y�J(� ��=��w/b�A�i ���B9f�	wGc�%�"���Sa�t�_���}����[��q}����:�	H��O�cSƙ�v6~��ߛd���hFث�ae_�R��[/���9q"_������v����3�+�K���RI�y�n����^�ߋ��&�d���B3��n;�:]ݎz+�Ab�ᛛ2�{
rE�h�; |��]��u��B���7�P$�Զ��� �,�&�f�R���l���;J��x�s�����5�ܧ�s�#���{��d���O�ц1u^�g6S��@L�Pß�.a��qUfW��,`�sc�G3�i�P�� 'I��n�5p���/
L�Ni�Y���U���*��mfGs8�����Ac1�m�a�J���>��v/��_Hu�Ŗ�s��*�7�F��t#�u��ǌ"_jrM�R�j���i4C�#��՜�j��w��|4T�r�ɐ�+�a���lv��� �;�F`�3�Z��p.�wu�"?��h:ћ"
��5�}%�7xWz�;���щze*?ޟ-���n;L	�E��6�]Ĉmn�v�R:�!��.����.�Oc���c�-�ϧ:d���I�%���!8Z�@2��S�6�r��T���z�/4��W���y���F���q�^�υ@�VL�@�Z�����XH��9C�NY
+������� �/�$=ơ߫g*5eV����DT0*�+�����[خC��_1�IWOEh��̿���=�K���_�= �g�l���q+a��1�\�s�Ϩ���Iq�.X�@�i�1T�ެ�\Λ��gބ�2�~���x�J�^��S"(�+o�#�� ��!O�_;�~��I �4(K�x��Ҿ곧0���6�=�=+-��V˰b�y_��N�e\�C�w��$*��
�υ��w�fnI`�����L���J}de_������*��Q�_T� �> �ȧIw5����b|�S���ʏ�Ȧp��.e�h��@�V�tMmM���V<�U�rB��W�e�魟�X�c/[KnO寒|oD�h��8AЄ?n&?]�=Ɣ���l�xoe-|I}�n��P�*�0��b�u��HB2�Y+J��L�m+����}���ZJ�yo�k���M��d�O����;�{Sn�X�͑�@~}�!w+��2���x�ĵ̈́���&E�E��&�f!=���)aZB���-�Q��d"I���a��E�]�魯��"jwAe� p��bůe_�����+ �[�W�M1R�Q;o���1H����+�Xk���&x�����n��������[xSyǘ�x��&�&�d�.ͦa��+�HX���K	����`�M�\g�t���{����F�,��e_g�%J�I�z�#	�o�>����;+v�X�-{�KĘa���+s�I����k`��#�^ܡ�j/��������{,�YZ�Xx��*o5KB����"�
����!��-R�c�'d�N��B	���gO�Sw̥��^�yȢF��*]@(�Ȍ��\g��D�K��TNqoOL��ґ���Ѱ��&���q���>�t���~P"E�jV��}6�n�T����IWN(��d�ݺ]�� �@wNc�WH`����Q�[엮W<T����M���~4x���vf��Jc4AWe1,�R�5J~�NMlFq{�/@���_���Bwv��@x��9!��{��a���l>8 rQ=��霔��� ���5�`;w�h�E�#�H��P~QV`ݜ�������x��y�,���VR�N��o��\��i>[�L���j��vP��u��f�(��2�d�Hv�QE5=̮�1y��L��E�d":1�O+i~ @�·!�i�w����a��jf���[K�LF\�<�P��yZm���{���k���,GN�!q��viw�љ��}yٴ�LZ���>bd����;� �&<�ׯ�u��հ��^J.O����v>
���&]�WPӏ)�C���H�R����xmS,Ҫ���P)�Sp'�@�ε:��b���v����l�J��Y�R4��1��[e��]q�~�yy|9
$��h�&��$A'���f;�V�(��f�9@���R�?�c�O5!F���"���׫�B^��S�'P�w�O���^c)/OA�2"E�>��R��N��ȋ����AZŞ�$�}B��+B̮����5w�7̼��E6Pyx��ߪ���S�Q�I a ��!�>%.�8�dt��AFAm�YOk^�%[]�BN�(�^��4%:ɮj�=�Ŝb�{Xy�>�i;m�ƨm�U��dժi��G��70�ٰ�Φy�;�i�*���b@���B�'*���l��V���+�jy��ڠ�����|BW���`��O�L���SZy����)��,wE�H
H.:�g[��v�����C�c݀��]�jx�Mc�T[+�Z�oc�5E�L���m�@�^���.}/�5�M}��Y���pjL�"���^��s(-�yN��$�$T4E57dq�#M��;Hc��{��xڬs��[ZIu�|�v��@0��Ѽ*�ch���ܾ<���D
5��U5�)�{��bcf�ν$��}7?�@�MFx�-�v�:\�E���b_*��%l��2R�7/���[ȆE�Ǚ/���bf��E0WWmFh�,~��K!�5��&#]襦�����z-����M`�X�9�h[�R��+a$ܰQ�!f�޸�ܕ�VZ�[y6�$���}���ǖn����,.�xr����)�>y���	Ԁ�>���C�[��XW%2x	�;<5?���d���!�P���X�W���dr�հU2����kZ
�Z�������T�y� r1Lo�kƍ�����_#���b��!qN��8h�E�d��;i�Jؼg��y�L��-�+~z#���G�Vs}p�(r:��ݏe��9u�KdhL8ئlCk�/�-�b�����A��m��T� t���"ϐ����\z��f����b���]��y/������0:�؋�8L<��ah�K���\�9���[K}�&��?��(�d�[C�{�kA°�]����=2��^�`�Yv��������(�Eʜ�OG��	���G�W��ie�q����0�a5�x�9�|k?B"�%�;������@C�@�Py̟Ҟ�3�8���T�̊m���Z/ic@�j}��qq�׻x��A���H���V�a
 ��C	S*�|{.��p-�٧�����`�;c���K�¸��A1��3�f3�ŕъ��ٌu�00 �>,������H��6n�6_��G���	��n(��|9�`���\�Lq�v�oyE�H�ܩf=�����ò�5�����y���O������{7�)��c��źvJ�ϡ�y�5�&�_]j���<=�n�;3Ύ�`���
��X��o��xQ���{]&ü~w��ѭ{6�WCfs�� ��L9�*}>��q�D���Jԏ�9p��H����驭�&�h��L�_��.{!'�,�suK�_�.���մ�b$�2���@�1@��h��Dߢ��Q���BC�*�A)����Jb�>,���w�ҡ�ٺ� ,+'ɒՀ����֐���)���`����pd�L�<v\�}����$�ᤏ��ԊL���Y��kv2L�ݑB�� ���y�Ujz�/6h0)��%	ع����e<]�x�u�Rf��C�2���E.��zf�b{���K� ^N��'ca��G]l@<���Z�����v�csD�\	�0Z�X.����)�@_[_J]xZ|�(�DF�L�¡��.�/1�����I&IVNI��A���g���C�LY�k��Q���u�j�
t�5�U7؆�����7N����x-�m��紮O���_U���psC(Yt�^1r����WX|��{$5"��C��|o�ߕ}jr����&']�и��!���p�����Oq
�z���
x�g�<�Իk�%"3�@eVA䉞�k��,�Op��N�e��o�����Ac�E��.Gr�f�A�%]º��[����%i<�$=$b+JD��3RiE-�B��	������>_�ʤ�ET��o��=xGtTv��K�f��yS�J��'�d�6e�$F��c��Y���^�
t|cpE�&�K��B�m\�j
�ٝ\�=y4�^A�DV�@�8��r�8��������v�+�!{��0��9.vi �����`s9�]������t��.���\�%��q�!�ɤD4���wokQU�#V�Y�Vc����w8�R�VU:E��)x�u�:�DfD�0�'b�C_��!T��Ad�K��[��q͡H,�����w�_�j*�S��됳�վ����z�޲�o��?鎊���Y+Hb	/���g��������g��>%����O�UA��ڈhoΓ��w]����6]0�JiB��v�R���6x ��Du�Ͽ�;���tfi��z���A���~B���R�G�7�hq*S	d�;�M8OX|c��5-��0+����Ъ�"}I)B���Jajt!j��f���O�QCوCy5�zM�T�e�eD��>�0�J['55\eQ�����*�U�B{S^��3Ґf �?�D�����WveS�,�%�;h���{yܕ�vHG�F[*����U�ހYZ�O�B�n�b�S<��v��S�PMxQ�$9$��)�@@g �ew�d/oov�ɱU���z�+U��s��J�{"�A�a����
�-FT�2G_��3�.�b�+gw����G���)���$��	u���0 b��2I�x��1Q��ɉ��/�_/ab������S,�O>��T�C�iO^��h�>���믚v�>%�<�1<M"��ʭ��
b�|M�"�{G�u�H���'���7U0���[f�%+���xĤw�
�'X�5�П�ԓ�p
?���Zz�w?q��b3%Њ���j(�`q�B`;l=����
-���U\�RAz*H/�-�x>y֠ WD(=�~�u�&���^![ƛ2�'E�PͱA���$vܑuo�hڶ+�E�����h_9 ���r���������ۋ�f�� ���$~�Y:#�ʫ#x�2�����/�Yd���t��#�J8A�Q�G��.A�G�a��Ma�]��𲫟KA����^Q?4�M
�Ռ�����.�n�Q�ò�⪺��0˹�T� @��5�	�[3�|������D����E�������S�7$=�'��~�°���g��C�c�q�5�̹q܁�ݭ���*6\�����Y0�!����M�7�UO��$�b0���'�v��m[t�I���?����K~X�t�1����E)9�G��Y�r�_{��J�vXk�pps����ʴ	�i��E|��[Ykq�����aY̙V=�,]�E��q�G���f�	Bcv���TW�A�
 u�2�$��xB'�8����vYb��Z6�\���6�ڐ׊)AJ��J��q\�Hڅ�Uk��2߻��N�}�s���B�a�3.x�����,�T��.���>�EH� �<����,<&\ц�:>7��c��͠��]hE�- ={3��\��e�:�*��)�)�[ �=�U�	��%��^�8�(,���9)�m�2�L�3��l�_��|���R�u$�R�/�B��T{����C�$Gr�z�c��|Z#�3��C��1�^�ѭ�_䶄<����e��0����/��5�o�%SAt{��:�?���������&t�+<7����4��&��^a�H�{+��t���.��n���h�;��������d�o�H�Z~[�Nـb(������),�_wj\�Ā!]�:٧q�#P8��w �R�Y��<�Yw6��(3�mU���g0��+F�۬��fX�$��
��n�-KNkn/���ߧ���oA��`��T��(�������Z&#Q�ځ������0H&ުt���z~�:ÙL�S8�0<8e���o�SZv.�}�q����:%2�WL����h,���k)5K�L��<τ/�:U��c�L�kò�m!�w,�B)B���(�]2�US�L��'�b�,�{0E�Kec1��w��FJH�;�'�;z��c��Ld�h}q����f��˩�Y�g���b7�:��m�nL����lM�)�˻���;�2u����y��<z��Nv;D˰�3һ�*$yL�ᎊ���ٸ����&��U�e��g$Lx��yo0�r���p��;e�ɵE����6��u�?��"�ܓ��3��c�i��-���bYh
,�=M�U ��Ĳ���MzF
���|CA�u9@dv��Ղ�)��O�KNw�"�1��Ԝs���T��g��)DK�?T⺹���$S(�h�/1N���yaV�#�H��r���{H�Q��ٺ����I�c�~��Ӿ�ק�I�aȥ	c��0�r�ɉ1��i&eoy��c=�־�(��0����hHl����?2���0��9]7�7)-����&< o;|�w�?H��+ɡ��p>K���e�A�{�Hȼ��8J�E�L��dd���/܊/�PO~��8�(�!"��vE��\cO�p��^�h@
h��8`�JeJU�E�{ʴ�CD��c�d��������[|z���Ÿ�M71�E�<�}�hJ��
��zr��ߤ��p{Fd6�)�k���Bc�����!��u�[�>��ݚ�rp2I���*=+�Zœ�����9�\�?�O&�]Wj��Gg��.�։�NNSߛR: ��%is��N����T1�LM���U�0Uj�a����� u��m0#�bl õb�[�έ:�yP��C��/�S��q8j������q�)$q��w�=c�h���C.��ab��I�?PB���jӁID�"��.h��ӽ��ְK߬)N�(:���>Lg��ޠ�u}κ_��2�KOI`��V�f�����Ф@�ą£���,hB=8DR˺'��p�r�3����F�؃W������T�K$�ʘ�M#$�i����Q�:Ź��Eg8Pb��z0S,f`���2	�#��!�!Tp��
�4T#M*��ڎ�_	���Dr@wգ����Ο�>sOK����-��#���\���G�I��{j}sڒ�e��~� �7S�8�H0Y�q��F���D{&fA��`���Br�L��pi-D>�+9��1�����%���G&b��D��hkH�[�W~
�����]�#Ul'�K��#��V� ո��{�������$�LK��&��3��(Z�m��m��z7��VAȘ�d�^&�m}[�� V��ö�th�S#���q�P��d�%��>9�'���c!�#?O?uX�xx�&�A����G��׀�����l) 0;31hD���������!r=-CȪ*��Vk७�H�O�h��m���x0CҸ}��WỒ��P˝Ke��#��c�x����H�E�`��dkZp�vQ�˯��0J����lÓ�*�������#Ie &�P:tK�AvO��pl�te����WG��H$p\��'�̑)��Ι��s<2t�h����F�8�Δ�%*7�34�&s��"����t�4l���Pp�CT3��q�Vk!J���{w�@�Q<�c��{B�T4�U�jL���4�+�.�G��B�v"K�o�2�%� hzg��?����?R8��$�r�/L2M8(7%i�j������/RoS�Ù3������+P{��ֽ���.��i�@�![�/w���%��~%
��P
�޾�ß�)kBf��TU��'���iɈ<h@�4�M���\]b�W��'#>᥉N��/S��*��fCo詨7T?9	�A�m13Qt�Iߏߖ�F�M�����v��@�-u��M0z�e�ÿ�b.И�;�5]f(ޙ`�b��0��&L1�7����L�t�Z!������2&l=Y�7�&L�I��&�?_�Ibg��U�A�c�8��o8[P��|��p�Wb2�n�sB<�=ƭ�3�P���A����+_/%�ʛ}*c���W�N�͕j"��v�tFz+�g�
Of�
SA.�݌����Mpڸ~ +����[�3p$�c�?s�=�:�s�e��<"�ln���o�$�6���V�X\UZמq����s�J��*��k����*����T&����-P{��^��?Y� �I���d?��(�E�}��a���cD�iz����p@[���s���Cn�637�?]M��`���}��!�$�:S:	Qe�2Ԅ��h��_�B�~���D������hJ�$�8��r���7$��+���yZ�n
~C)X\�[3����6D���~����P�ߣA�����p����d_�9����/�~̗�uS%3Ϧ����Ao1C��#k�H��#_�ú�{��@P;���|��d���t�r1m	�q*�SK�gI�t�I۪� ����Ԁ�W_Ɓ���TtT�	O�F&x74;cb��[�O�'�ح���#ud����(��f���Q�{�~��`��VlTX��a(�iE�~<�;�u�J�hd��MtHq��<7w��Ť@6B2S��}�lXP6*���8�d� �#!h��=�Gi�85�^!1x��He��(T�*��H�����s�!%�B �jFw�]��H��YXf�<g�t.I�uW`�vl4W������`
8Z$�l������'�Qgr%��ɟ�����<���!�a���WD�G`>���y�>g�x��m1f"���$��4;�ኝ�)$�;0�v�Z�ڲh ��,��R����

)~���yD|�S���~�a�����Pe7IZ�C�Ii��F��2�{��c?o��ժ\����+�Mo���*Z"f���AX$�����\�9	���'۱�/ߑ	�T�y[P�'����guɕ��.��a}(Jvr.X�y���G��=��ٺGXR�3pe���r��"�Q�^G�6��97J���ᢄЁ�"�ATB1��"8Fg�U�o,�c��m�"�Y�И�4c�b7�T@��>n�7o�@~ f���o������Y��qn�Ձܐ����f�dw�-���u!�fܹM@a�Z����0<�3؃U�Ў	<��sS�y
�=eC�+��������S��+27�XAK��F�|T����5UZ����}!�$0Z�ac�G�q��a�%��{�u�F):��H�4�1��ޡ��?x�B����b��!���D��9��5���V��4o���A;��3�0�h!����PE�Z���x�"������Y]��sd]�.%5�;b���)X�%�8
��\�\��$;�����-#ʾ�Y���P���;�9Yw�)u���>^��8��emf�]w^�������+Q��	�L��f"8��[R��x�B����!��;�c�[�� j����.��D1�^p(���-CQj&�^�G&����Ό�b��n":����i$��'�~2�O�ϡR@
[C?��8i��`���?�b��z_И���@�}X�E�̜x�? s!K�6i�2��R��b��d��}Yy��&���Z��%�l�I��H�C���n=��7���������-n�'I�V��{�[��vIt���A�t�hT�f+=-ӯ۬�syF�S䃝�h9�?ɮ��j�>h�l��л�6�+$�`���F��b���U�
/2Et��'A��o!,QGʔl>�L&�Vfg6Y���_z� �}��0C�f�i���T�A��0@�W}G�%$�d�q�_`��I*0�܂j����<Sy�_�dmޠ��[�c�2��`v���'q9��z�pK���$��x��i��<E���sO����BF@vEL{ކ�:m���{��b&#;��6�y� \�z���[c-L��F�t r?8'�p^��z��~�e��-d-��v���	-����_-�c7C�LF��j�W�;��]g�M�Te�g�ZY�3n����	���7R�R�J>%;�&�ߙ���s]kp��&lt�Ű��7]QH���d�z�����x�']9�B���Vj��kA>{G�����v���fybը���T�- ��3�u�=k�n��'�hZ=бl�y�ş��h�"�1B���֧�-�B8*���]��(�>�Ug�A�_/��:HJ�iQ�)�i��׊�"���/O nRb:|FC� E��j(hs������Os���i��}|xi�t�?Բ�!.�{�����r��~�+&>�#璘B�ߒ�{��'�W�������ޮ��b��$�o�&�C,:V�������}�$�yXv�Gw������b��0q�x�(����!��Zz�ȠTJK�G������� ��nЊ1m&�b��R���m�<�I�z�T3|�g��?�b]<3��FIT%�n�Gz!k�޲k�Z�d���b�����2�GJ����5���됕z���.ID�*��@!�2^P��d�i�*����;!£$58%v!��ɑ��tY�Q��y�Z���0��֏�V�rȣ��ρ~Ϊ����1�'��Nn>[�^N~'��bG]b5.��|�*T�ї)/������W���ۇR9�=�5~������
�Ҙ�c E�Q-K*���C�����G�\:�kl$г�Ĳ�]e�Z+Zꥡ�/�`c-�����|�>�k�rRk�*��Mq��;I�x�nJns���+�
���3�Kݽ�A̰������E�C�׺3�_��=��)��cw���0nzq"'j%ϯ�ji+���l_�[%�զ�Yj��:�tQc�i��&x�����e��K:�Q�rL�t�����3F9ƽL��x�F!�''��g��-��,�)�J���m�r��̲�'� �+��B�uod�ȼPs�O���AD+�:g�~3��2iDV
Mk�j&����`�q<w"� �/9\�,���;8%(?1q�6FK�|�_��^Y���N!}f[�>1�oflZ�. ecC��:���)+�D���~	��f���y�\N��Q֘M�|O	2q���,�~e'�K�[��B��U%��*��,dR��:�n9��ݻ��j���l�Hp*m��������e��@��NH:ʧ��!C�/��Nz{�L�����K�5��m֚z�ς����3i��� ���$�Z��`����J`���>L�g��zrM��T��<Ԟ'����j�a�e�5	�{��ܕ���xGqW]�"/yJD<VNװN��B��e�uB{�έ�q�b�������y�B��RGY�^�f���|��7�V��
(9r��`d����S���\)i��sT�F��-$���A�vU���)6�Ӑ=lRV#���_e��U^��o�o��m�`��~��c�9��KkV��x�e�u+Ɍ�T$�m�ǭn�=�F��v�͖�lX�D֦UD
����D����k��X�x:�Qj@�hE2A/��V�@�=�$�۰N��%tm����Mo�4��ց$�!R�����~p�0��aj���Ze�H[es��p�͟Z-��?����8��-�]F����1��L��	��A�O����"��RD��y7�D���;��b��tMM�us��\���Qōu���NM�,������B.=-Y���y�j���ea�[?^���M���53��0��z�z����`�qc�WeߏV��s�Nfͧ���M��j����#92�(7�H3/ӻ,���#���$�/���?�?��#��:v)����^�p�cS<�`R���aJ(�o�]�7zy��ƒD@���o�J�Lq����]���+w��r'�a�U�;:fG#�+�<�o��[���Ԁ�2��0�s�,\�w4W&yT�灺)j�Z��.~b�ЯsNnpi^^���	$� l��D7LN!�6�g@�JB~P�H�Q��^]LZ��Ǆ9^�7$���"哊d�;Gv��w��nH�W�8�<��W�>�e��k�tϻ��7����j�v��"��>����j�O��g1����w�/*��dPS��Hc:��lNv�71��g6���2��|y>��8�������ª����66���J2�d��Ӏ^_D��"��@���zo*��o4�3�pʠ�HSW� [{��}-v��'�F��o���/	�K!�$���~�ƭ�]�
��|ъN��u��z�/K��S3������m�;}���^�̮��_�92ج�~�j'���`�!�I��3�|�Py����{ `5������"����Έ0v���
��'QM"�z-������exF�8��l((�#n���י�f9��%Yܝ<�~
3�ͨmǡ[$�VS$o[Y�I�i�v*�ZP���?��?j.��_HATֶ[�XP�. JP5�ɺ_�J5Wg�|mM��z���+�S��J��r�dO�"�KP���� �"��L
�q�:��! y�9�N������	��
��lw��I�Qe�^�D��~xg�u'8v;�>��>�����W�e�!!q��?	�>،�~��Vyw޴�5;W�Wa�n��TL�;S��_��w�*� �bm���e@��
'��J���x|�)H�����H��3�sF����-a ~��D��G�-��__��g���rKt�U��}!��5���qp`�
�v�Y�j\�Ò�����-����Ec���HHb�iTZ<���[U8�l0B�F�%D��@P�Xi
�k����AH�~�YB���ֹ��6k�xo�]�R�G���̦�����IO�@%�5�9�F��[��F�i���ҡ��k���bӚw�i���0���.�[5/k9]V_u6\�z�����H��vq���p���
�N�to�`�#��	.�٢d8M�bMJZ��:c32��Y�BD}@�ao�,wH���B�/�o �n�1�Ѷ�$j��
�-s��ֶt���1`/�Bnԉt����0�j�m` M�Ȅ�I��,蟹��?���YY�8�%���O�\U�]�t���T81�RyU�ɱ���	G�lB�Z#�B��`N��;�����V�e�;Z��Bh�g���S��E-�d��?�b��Gr��[e���Ǔ�NN��`�5fY�1('�|�]ԑw�"qI��ŷ�yʋ�Ip�p��N9��Hɿu��v��;Ɇ������c�Y\u]�;�x��%��_e>gY��-�ZCXO�Zy��3�����ӫB�G���[ܰNZ�j�&����'�Mn�=�[���4\�{���\Q�)L8��]$��K�l���%-�g�T�������P�S�2Oh!]���y�sgxP�ѤZWi������7���n��;��&�a��:�_�8�j�/��y;���S�DV>���5UAF��a�%G���MjA�h��w�4�n/5��19�~R܃�����c	$�3�����U���zγA��5@�Y��	���8�����\&��OxܥPzv["���K�ۉ}�����`�a����t�^."w���a�.B(�U���N�!�gr�mSU$�
�P�S��P��v����a��~�"�eRY>ŖlhRz��kf�bT�ۆ�f�ޓ��AN��W]���p��h>˖��� jn�_�� �c?�.��
6b����A�P��:Ag=�����{�V.fc��f��{S%~N���<5Ϫ��`rdk.�+����d�X�ǋd*�d��V
1�ut�P�C�� �X�@ �w����g)�_���
�2��O�T�� ű^��,7.�&�T�u��@���[%dr���O<u����'_�)_�.��nǥՒW.�yJ5�b�mf������#K�J+)�XV�qܹbʙ�$�%�N�ƴ���a,���V�yx������͔��X�a�rX$6�V�UaJ�F�th�V�1iy������L��'��9M!t�mPvA��C
7�C#I�r,�U�Z�[���?��K"K�.]4�Δ��m_v��d�n�6��=�3� �~�p#r"�*�v�ee��Չ�$t���_��t�S=����io�f)zc��.�AY�l��j������}�$�U����L꺽\�#şݦ?��ud�b�P.0�5։:�󣖁��|��6(ӛ����돜^�uq�R��|��Sxw*�䜗|X����p�ءۂ�Ň�33�%6��W�>���9���T�J�O2Xtvz��<u�ۙ�}�vo��P����� �]�8 O����i��l�� �ޏ�̊�8S7g���ug��ӣC��\{'R��1�js�Ef����V�ܡ����Bt����9�XF�i��������P���r[��b-v��X�$m ?�S��{]�G�&�}Zc��4����U�l:r^�wmq�k"�v�'q��Vl91u�	�v����Tş��%o���^�s��xi��P��_F�}Ȏ���|d�����˄��*O��7�IM?,]�������[��G.P��*S^`CH���Y��ҍ�+�w.-qo%��@m��J��)F.8���3��u�"�Y6�:z�]�}*�,q��E�O��­c����L H�̏�P�G2.7Ϋ���0���2p�¨��M$(�� �k#z�������o�yh�d��`�$��/��HxF�]�� �lS>����]�>M�ͣ�����g��,L=��/�P��|��H �M�K��r{�.h����R��gC�ͯ�4G�� M�8_�s0&eŷ�����^U�^�e�P,�GD�dxr������/*�G�r�}yC����h���o�����E v<���o@��Ҫ9j�۠Dm���BQ�+�[>�^��{y&ԔQ0������O��#;2̖����T��=S��-�t.|���d�a�S�����������F���~�n��j��F�<��*�U�<D�Z1o�HF5ƽhb(���OMae��~�����ӛ�[BǛ��Y��qB�cIì��R�j'�@t�;�( eݖ%PJv6@�%�@�dIu/D�E|�g6IA��J(�
*�F�s�	In�U���i�:�>M�V�b{0��Z��b%���
�� ����=���bI�(q1�j�j����X�O��Ew�a9�������1"��\xZ�v�����K��ms�/����I r�H���M�^�v%A��T
��q<�Xavς�(Ltz4�\������Č�*U��@�k��`&�%v�*�S�jL��9~�g���,�P�q)�Ą"�BL�~��ۘ��%��[���/v�EE1)�ϟy:=6w,�<R�����T�����d�8�i�ᬿ�~>��B��� �S�{�E��!�3���-|)��vCS94Sɩ��a�~��S��q�Г~��0���=�J�`��3�D�"�&i#Q,�Aȥ�'�o[a���P�L�U��j�)>&>���Ht����'�r��0��h+`�m��ʼ�XB�Ws4��}�8\��=ZC�=�`�E���1}�h���è�?=�c*T�o:�l�
����o�v�PO���~�Hlm,�32���"��h(��,���%�^�¾	�����b7�%�\"G��R�ֶ|ͦ�Q��ee�F�~_wq��� �x�[�� ��	���&#C��XRv)��DgJ ���Q�R|�^|g��
�$v�:�a-g�I�=��a=uO]�Q(�?C���[}zl2��'�(�Z��<k�����R
A1¶<H��I��v	Jҁ�O0_W�oB[���&�a<�(�G�_Hi[F�c�������6�Ì�%�e�$��*~��!���"�^Xs�_R�ʤ�]��}�EiX4�
�V�,��!-B�6��'�)����kq��+Ӥ��p�w?�^�3��F1Kp
���$�"��`�U�Ui9~a�	�mf�h�Ոb���	�i21����ϊI��=���0����y���g�uh�Bͨ��Ȱ����ђ$�lWhz�WmB�CTa�@{zhV�Q�my��v��y�?�����A����~Y1Q��=E ��C$��4��C�b�����[����J2d�ض�3Ӆ�T�}�.��"c����8�?@ Y�J����?؜�HCH�C[���&��ہ_� �J᬴�y�谨@C���!J`"릊�>6�"�9���	����c�,{N�y��c���}��!����K�|��Ǚ�d��r���r&�O���	x��Td�|�ʔ]dÔ9-�M�b~��?���4TW"�b��{f���8>�j<���L��{G:�F�3�	��Vp����>�+a[H��W�	����`sIHo
�ds4z��aR���Y!��͢��w��i�����&�	�0���C���yvq�4*��$ ����Q7�oW��Q:��Aپ��\�JŤqX1k8�Q�rU3���u@�������J��7��+W�>�z/|y<=�B�f}>�j�`�!���ʃ� )�^f�hv������қ��@Y�m�(��>�ss� d8%���,���ĩ���P��C��ҕ}Q)�#xRa�y(��^!�-��4$�7��A��r�d���}jg=�(���E`�#8	��"�.%�m囸��/��>�����'L��3}�*��~�{ ���w>м�n%���5|��w��?`e3r3�R�N�L�`��<��@
uQ���5�B!�+���M<���ݠB�&����(�m��`z�*�-��
���'�Z��o$��-�D�]f�~� }��g�O�H�s"�����l�T�S'��[ƥ����s�g��ZͷQ~�Z�DR*JcH���r�>��l�e��w ��Ԫ���~{M��E�Έ���fI2.�Y_P��	\��9F.�1�1Γ�W�t!;��d����*��v�]��H���ꢠA<�W�c8w-�`5�_��ޙ�����Ui�9�7l���`:G8��uth���kTm���q��- �10TV;���I�!:��x�*ե1 �b��E�i�
J����j�/�_���K��emj��z�m-:�ʑP��^�nC�+�-���8WTƌ��ѻW����O��\��sۣi� ��U�⁖=dpI���O��-�D�$��B�������t?f�g⽃���nCU�Y�MK�i�Ѹ�M�����ƙ�ҿ�4A�CV��"�>d�)j1hQs�w�{��o�g��|�~��̱8'v��tD&	��@Y��o�� -����C�e���[iƙ���j�I�=jI�cQ��L����걀%�_��'�z�'yX�@JöW�����X���R)I�O�a��^�Z�Ǫ[I�o��`AĶ���������4��"gï���QL�8�cG����]��_��bs��iTXz��+k�ͱ�D�S��+�j~!:;�j�@__)^��]�iqV�d�JSP6���&������]��g:���U��Gcz��9��f!\?KU��|���'����V&���EEU�%��E�%IQv{�߂��r���Z�X����|Y�7�n���1��'���|�Z$����Ķ$������ �a�F� ������9!:��)m�bI]qZ�pF��9�)�;���2�Rց1��N����n�w�`�&8��������U��G�)�;�E$�f�x�L������O��	���q7�@v��TS#z���x�i��U?~rv˓g�@\3wHDUXr�ܴ�K��]>�} �'ygV�/G!9��l��o��G;�(\s�VC�PtMN�8'�Ԁԍok��.jF��Dş8��3���e��[b�S�"������"�m]y�d>x�c�8�%��h�#xë,�:�`�6ڷ��%�ɼ\� ��+UY��J���:�c�{�eѪ8�䕅+�sq�wl�O���?��d�W����Mc�|Jn�m�� y��k����*�ehQ�E6�U����z����.q��C�;HP��*`ʳ��l��<�=��&룾xw�e���W]���50_���;���"� e
�� �s0�j�~�^����tz��%��hgo��VQ��b�>\��+�)1Uk@꘩i���0^M$�JA-ʁ����+�=����M�p�a�A�d!#O����O�ʑ�j�Ыa��-�.���_������a��j�@R��>O>�3P�����2�"8�t��z�|߄��1JS	2/K�.������ω��Zj��s�f�WWp���� �_�YwV5�L�+��7J~>7��(z�C�J�����+̂���܎�u���A�y#dg'�
Ʀ�&��ǟ�?w6������@�+�*���&�_�3+����]��C ��9����@^�&Ⱖa�1���(o��Y�u��x�S �v�x^4�	�e�b<�Hq����ׂ�`7�;X���v�c����kJ�l�(���S�:����,���K���]l��DW��_L<TELH���Y��\e��Y	�-)�~T��7�Q�L2�&]��Hw�=��4�tŌx��T��F�D�ı9�&�v��4KB�v��Х����-N�:}ЊoO�J��#|J|�Z��N��'oLǜ��zK��]CN*�F�-��w�DR�1���Y�Aӥ��|h4P�%�o�Eԃ'��Ӣ?D��G�X�хZC��\�W�J����x����z�i���-�&�������{�����g��u̻:f�v��Nf0�����8�����n���:���)~j4��
�V\S"��aX�3w�[��Y^#�6���$��϶(��!,�ƋZ�c� g��؊�������v��L�h�/�x����Ԍ|^6��| �����`n����8[���$�\<,�S���[�ʪ��J�hm~��)a̤dG�-S�� c����=:A�kp9��-��$�GGT1u��hZ�����\��z��`g�h����� �z*�g`H�D�`�k4����u���C.���r� �Iˢ ��_�c�hH躬�4�JI ���V�&*0�2�����?���s�x�B�q�o��JgM��M6�F���f�u��Z@}�bb��p;*`4��RiI�������ꩯ&��Z�d��M4uNΰ��5��_xkRF��Ybv,6�C�P(x�1�>m���T�)�8E2#� 6+N�M�?���;�}�F�3�������@��x�P����i��
�%��/~�l(,�����+�4 ��:1��rk ��+���p�:�js�����=Y-�z̄ߖ/o��M�,�LfJf��~m�@�*��ò��/��CI��$=�'��7�Lf�:K����I+>�ޞ@�������d~:OZ闞1�<]l��ې��jKK$��#����z%=�jO�v�Ne�=wv�Z��:��ݭ�
�r� �Yn�m=�U��Ŭ-h[g��#������Fk)>Rvg���3I�~L�0�uR�X��I��:�! ����L�A̵��g��g�&��$���S ��/�����\U2�ߕ�����:ȳa�$��&�~�pFlݮ�|��֚G0`#�V^�,�Ϧ����r�(nCq�8|g�Z*�V��������+�Qu���v~ɱ
޹�&����3޳�W���pV�-����?C�ݎ�����D"�!�ZD�2ϡfC���ۙ���*��03o�~��\U�\X�Ad�p�M����J.7�yu�x�ڦÅgCw �7R�/ɀ��k֤-M�	��d�!�j�\��X�c���G&[��!�1��	�ǒ���ܽ�m�Oh-��OJ��vR�{i9ߤOK9by�u}p�UM����M�FA��A�e�}�/�ߌ��T��l�Y��r�-F�cis��ǒw��$�b9�#KRJ�1&��i���[����o�ׄg��]�Z�%��Q..T#�1��!��Ni���8cnJz�&w��d` ���Yn���^]�{� r��$/��	��%M/��%Ik���/F(ް�s�-�3eC	Z�cj1֙6z�z8�f�5�K�4��XV'�!�^ԓ�r!Z�����ŏv��B$?�/ݾDn����]��0b��ؘ���S��y
"�62O�i^b�_�~%R&�7^�0�rJK�%��Y�߉��]?n1��q��X�����Z�����2��	5�V����G�hF�����S�T���[�7�$<���m%'��PڬY�����1)K�T�X"fA��՗=	����T�z����k�
��TP�2�!�i��Q�ϊ�q�@Y�x�/�f��ຐhL4'q�y�,p���X�~[��ۆ��~ۺ|���w k�(R����M� �X� m%^�#� ΂�C����ִ�)�lHE�nOx�47ѤD4ĺ��AX��BN:�Qًз��`1k��4�:@}���6}D�zW`j� TO�YT���"���������A���G���r��!]�}JӉ���O����t3�Pt �-7"L���-d�'MbF�����^��+s�s�9�r	y���'��K����x� �f�#GJ�Vs�����0�u0"��M9����KZm�-X�Nx�P��/^�2�����z��&֏=���
�n�h�x����r2L=���I���<�5uI_��n��3qҼ��M�<�'0�ӺC��AR�Y{1-��D ��C�vӠ���߆l˄e�Q���;���(��!Uc2>|�A��G��'�A.��n�Q���-�q�15�Eyw�5�w��h@�M?
.d�S��bm�޴�l��vs�̋H-��&[s���Օ"�;�B�q_�(����>F1$����
Sz��r��q*����0P�;�#��h-�ΐ�zd����%�¬�z����s^$��ռ��B���H_|��&[)Yv�E�\���&��,/�EQG�U�uuF �L=��%�c4��o�*~jr �i��xv�-*b�W�]N��3������2Z��vh�o��f2�f�n��'�v�����q(�2��a0u�-hҲ��tη��8P�8�t��x�N־\hB��3C�3 ���5g�{[.�u��a�!>��Wşu@��y�Tx'�c���b��U<�)�����[���'��K���` ��������Ǣ����X�>.���j7��_f�U8�}�.Ǔڒ�t�������N��>�+Ɓ�RT8$��ں�L��)O0��c�1�;�����`3ߤ_~Os�#{Z^{9���U+V�/��I��R�p��*]�n�PQ��{�*��ίHf��͆;�w����G�nLn_M�Vg"���H��B�D�ǽy��>m�s�1u�z=:g� ���`B�1����"Q T��S�)�v��J�CJ8N�Iz+�~q˳qio�i���>n¦HA�\X�2U
A���Uy[��<ȓʕC'�jT���E�_�����Y��@� ��~��~��ߟH��Z�����<�gV��Z!<���)a
d8�
K[�};�enc��7������2c���?��$�⧾ό��j�5k�z(�!����b�v i$��\�4�y� ļ��5���1ᙎ���򹽸��!O���V�C^���*��ঐ/K�_M. �K�9Wۗ��K��iDO��i�̘8xd�]������O��z��LøHʑn�^�yW֑�}Nn�{��M6�m��l�*�����8����j�i�$��g���|4��^�C}W�z�CO�]L
zY{��WJJo�ӧ�㜴ݬM�7��^[�y��@���~�6���^3�K�_�Ϣ��]/ۯ��U��sh�@tr�05����I���ʺ�}��S>��_ؚ�RI���)\��J6��C���[S/;�'��\^}t2�^sݔ9��c��p������'ˑ��<9�Z�w۞�G��?2Fj�bHMK\�E�K��(mv˟�������-�	3&��T߃��ҫ��C��Ⱦ@��~��%�υ�1���8����옠i����_�V��9��s5�G� 55|��xR׀�O6$���	��85����1��񿉔����q�c8��4
zM��nLv	�l��K)/X$VY��s��|=���������� �I/���<���N�����I-=�_&=�i7"n4ZVD@����|P�����9���lLh%� Z�e���ל$���Uq`$ʗ��&ϔ^!&��&@Q���]|���>������ك|d�p�X�/��\K
�m�dބ�Ԁ� ����Up����T�
5	^ٹ�K+m�'����1�F]�_eqC7� ўH0F�cU�� �_A��ɚ"^��gϕn�G+O�5�Z���2M�|��k�M��D-����̧9�Q��#j6ǱOk���ą���W�I���+slC̽�W��.t����jE:O�z m}RWÈ���5�{(fA����
�L�mŭ,V�@)�r3Ԧ-K�"�1&.S�Y�Z�������׊�����|�4�hN;�@��U�"wĔ��	I�I��y��W�j�ds���o��Ѿ3��Mx�����Jyks�L5_��η��͓�� r�4�?�]/���M�W��t��mڂ�qއ��֫(@(�,����Ij�ρ�6����k�^�,T�
j��7��-��`pk�">�.��+��r�HO�ʰ�0���0��p��D����o�>�8%�����O� �n���(�B�ĤR1x_̞�Tƥfk�_W��p�t�T%vE4�Z�z�Rx�<
�h�x������u��$����U�',^�5Ҩ�|چ���o=���l�8T�H�����-�c���D�,N��Lc�/V<v��$}�6�����T�[�!&�2����װ*��l�ӳ$`�{H(Q������\�I*X�����:.~���t��A��� HN�B-	���&�cՁA2�;��.U2��7d����,I6a�<��z.$J_{��*i�Q���h��B騀\_�W/�֢�Ie+i(��yw!�Q�vN�����c��OC��\�6�L;��u��Y��;J�K- K�6 fS��L�J�Z���x@]�?�l��I7~�����5aL�-[Ƴ�=>&r!��\>�2A�5�L��9E��71~�!�ꅃM�oy��'�|�qX;XJ�;�+p�~�qU�����>��xmQy���V�npp4���dY�ε;�:����e� �#��a�c5ֱ��C D��'P1��i������mU����$<"r�6��>L�kХ�괥��X���Y��cp�~�:�_�\�'�.�GS.�I��ɶh�+fBC�J-��V6��P�I�)�Mx�2� ���'/!p�S��ni���v���x,�����2t����T�&���f\����9LÖ,S��JEdNd�	U������̬__��T��У�7���e6P�� ��2�
=�j7 vG��«}] ɺ��}w5��V�����A�n$��`�5�����M흹����X��Dq��6��7 �;jmM�R�`����㔢ȗ��%�By�J�|0����}8����ll����Y��Z̡]b/��Av��xG#�)�[��	q�#,�T<B���g.�5uBۋ�r�λ���l�a���N�= Z�C<dE���^�+�p��EƬ�<�����_�:gNB��=��2�-UkqQ�ED�9ڭ����k^ߔ�`�%��-�#�Hp�@I�B��p)���n<��D���C��H��p�;��O��Q�j��?Z���D"�Be���|1�g���J��{�	���1��tq����e�|+�Ƹ��u���ګH#���LT;5�h	o��C�Q��PK^����qt���J#ԑ���s�Km�³܌h4��o��o�ӱ���A�2��x�ZʸPa�9�oF˫IX�� 0�B.=��H6J�oˑ�#��ŷ�d.׫0�A��4��<��|��"6\�дu���RP[%��י�	��ke�3��-�J�e��Z�֝'�Wu�x�н[�����sV�6!���=\P`�� ���?ϖ���<�>�5i��Y�li�sޗ�Q3�r���� ʟ'�`(���Jť�?\��,���Pm����[jRi1l�j���"�N���(��z\m������=(��P=��
Dt�x/�>����R�R���b�j�(i�b$9n�������^�� �#�9B�IT�_	ᴳ���:֙"���'j��^hlp��*��X%�]}w>�<���<6J�@���Բ S� �I�4�^�����_�;������닼�k½�#��҆���e /F&_�qUr���(���u{�v��~�	�n�:MS�Z�����Dd������CT7iy�a?�� <*@s�4�ҍ�0�f���*�9��2Z\0�Fg�����n�{8�b�9�w�Ǉo"b�
��rt�0�����`Q����Z�����2�%�tx�4M�1�N��x]��G�A�z/��K�Wl�P�'��Hk5�y�S"���3���'R����C\��w����cE�.F�и���S�Е�%���U��r���~\�f�r.o+I���k��ݽ�]��GGG�Ɍr�=ܥ�����>_��^�	0�䉻�s�2�`��p�|�1.k�[㞙b2�J��w]��*'3��7$�DҼ�qv"�d��� p��~S���v�g�#<j� ���F`(��GQJ��Z�"���b���y�X�_l�bƅ�u4|,kP�6ҍ�,��)���Q6>6�"���=qp@
K|�<�|��5[~��?yv���t2�	�Vg0З�[/�#�	a��m��d�55��q���<��W�0��d璫
4�"ڟ0nl(z\�C���H��*��kĵ��⭝�_8�⚍ ���'Z����1c5ɠ�C�'��%�	���ܩ=�Po��V���\�ӓM[/D�S�s|��~�)-�(�V󲍀T�����.��2�SuQd�5�_�#��,+h�&�W��֐�D�����??a��.��!�5#�F�*�<�Fؤ�X�a.�s>�|�@�I�Z5���XV��\T�� B����O�5��d������������9�R�_D7��b|.�h��b��3*$b��VU�΍1�h`jIsN���q�h�Ia�d�	�j낺'�7�X���2z� Eg@��v'��h�]j�my��[6f?=�~E�䘾�3���sr�S�v?��?�ڜɅ)���1�s�����ȵ>���b���K+���9�}�uuU	�0�b�-�h���mʢ���Q�Uf��1ˬ:�;%t�xC#���te�qY�󣄸4�8sL^b�z�E����@��+��'Q%d6%���͌B���*y���gn�qC�Ȗ���\��e���mK��w���:ˌ�n�uj�LbwQ�� �nP���'�v�`K�� ��3�j$!��o#o��}����������u��e��ua��#�\.l�?6
�r�ؤZK�Lri/�����mj`�~q dJ{fZ:*���V����z��.'����h���k�=��E>���
�/�xտ�����N9tU��-Cԕ&ф[��$fǡ��ő��z�xAR�F��m���zac��p<S
R�C�7���J�_n�f�N{*�A(�G+K�L�Z����D ��XCh��i"��]�Bh6�gK�L��̔���궫�axx81��e³������Sp���}��>���o�W�$�(|����k�(5�V�5ˍ��p��"�>�ZU8-�2���,��W�5�`�޾Z2�S�&�}�іU��@0�[?���[��qN�0d��9��#V��nR.���_���Gh�^JU��ɭ�Y�n���������Zh6��+���ߞM�lV��収���m�QI
��<�au���Obݧ�VDp�t�F��0�lS�Q�D�#�(�m�������/��z���;D����蠷�EpB�Z�?�x	w���8�Y�(�@q"h(H.��KKdg
����Vޙ'��/�<�cMutй�����b����=�60l"?]��Q�́.�JjL��A2�A�J5��ѷ��ɑ�7^� @�kj����궄ܒ�k�0 ;�Ԗ%a/~V��JE2eg+�������?��5{i	|g�z2��ftI�-�@���u͔�l�|F�U�}����F�\�5E�����2@��L�'�e0:�Z���@�S�P��Y�� ��"/V���6���kE^�0�1���=�����XKVH��]|���r��@~to�x�r��ǧ��rS�ee���l#�AѰ��y��If�o-��,	�<�9�MP����8�D��m"������f�H@3�52h��t$�� R'i9HL~�IT&����F���_ˡ�7��9ޟ�w����� ��7��9�/��B�k��6,�¶���R|��GyF2�RQ���'[C�Ƞ��>��"gȲ�<�����<F#6GuÁ(u�~�(�A�|����|5����m���Q'`+��xղ�K��:�9K��5w��ASw�<Rd����LA�TҞySeں��hy�8 �w2��d�9�Tb�lB�C*u�3��xz�
?HG?x��+Q��K���Qp�q9��yEn���W��*��UNh�i="�v�od��*5�԰� ��T5��v�1ִ�D��X�*~d��"V�m�з׾:*]�0jy}Eöu���7'F����9 ֺx����Ҥ�?��`�����G�л��}JՖB�##|m�E�՛��#M_ԡ`���g�i"���Y��������Q��ݥ�U}����~Nk�g�jO0���a�ݯ1Z\���p�[�ven�.���%2��5vL�Q���Ԝ\�%���ᥞd�jD'ɒ���-���ip�%Mx��͢^$*���w��pQ��{}�!/A��ePy�У�S_?�����:'�'m���lŚ���,��8׀�����&�ز��WI6AJdfSe�K�>�]�&X�g*A]0x.Nd�o���A[XD�9 ,G����e^���#�T�;�G�C�J���!0g�^bf�|��rF'm������5��Q(v�m2ݝmG: }�0��\��o�+����"���lҹIG�n<k���v!3�-VO�M�,{����z�8��|�꼘�>P�F����gO��PI���wCfWA~]���C���U$�T��mUc.(��7ꓦ�H63�[��{�d�TV�w-�0qc����%N7���Z���%b3��B�k��3�'Dg�*�@�Q�&~ݑ�k�;Xk�Mr�k�K�p���û)k2��f3�� w��*;NE��~�K��[lv$b�mR �����>�m�&B�@��AI�NqOr5��,���4����~��o�=I(��5[-
I|3.��q�k��y�죱�@�4N-�F�D͡�e�E��i�P�f^��ŷf[
gl�vw#SJ�t,6���g�6&��.C��{i�bД�����!�(���t��)�{%���y]�겿����r����H��(Pdԙ(���Z{�_v�����7WG����i��a1(�E�<����zj�Z���3M��>t�@�;�qUm�v��t^�k�<?T�ֵ-��7c�����|~s%s��\f�,<�n���,��7Hn�şE��槚��I���1�S��3�JAEo�Jk��}��B
�1�:T��ǰ((��۞�gy�=.}" &�����[�U~Qc]��&*�����q�f��R��pE~@D;W�-"�Ś��;o�F�ENs�a��$a��Vﴡ��Ǵl���8��6/4u�;"U�s�q�,�J�j��>�:���T��*�Qz�$���
Qlf�?���OPh�5��@�-w:��aG5�Q��֒U�?yޝ��z�A�֞�` {n��"i��7`�χ$�Z�{M(���\ \�x������I�k��u�89��au[��ȯ�w�����9G����ᑂ-���|�$�z:�ݛ�AF��w7�ȑ .=�D������g6w��KPQԩ
�Ur�1�c�[�>�����X'�'G�~��N�iHJָ����� ��<�V'����c�3\����~X�	W+[�J�UK8>�wb�x�ߋ���ہA�K��&Ȓ��
+���`?)�À������I��rRJH�b��^ ���F�9�l�E��9��mU��(G��(��GIr"���,	�(/��^��H��}� ��<0�[FE��c��tq駯��Q8�2�R,U!�+�S��GX+���d\4�+��˝}P��U��S�9(^8\�P��<��ui���*{i��oʾ�B�c����Wf���+���a����<~I;�習���D��}f3�TV�� ��a�&�4�c�?�|����ƟޭN��C.�Hׇ���8�!	��z���0"���5�um��+��*mi���o��g�	&�&͵ �d�ص'#\�?w���L	Nv/)����%2[��![Wozg�"1A��_(��~�� ��H?���.��Zl�^���F
Q�̤�����|�"��r�46D��y➩;Ӑo祂\!��"�hp�K�6�u� n9[�d�ɸ��G'�d��ii� ��_�d=���Wp��`�}��"���o��|��9���ʘ��猃g�UcM���jyΚ�r�� k�>�vg���K�{���L��䰉���Փ�0s�h�}`��G&� qP�8�� �u�$[U�:�iv��Z��5R��<�1N�  �,�M0�ZȮ�+�Hj����Ӌć=4ͬQ�s"F*9w��9G�r1�ι���E$�[�m
49�ҳ�Fâq�N��0d��K�%�h�=�"ح?�Q�shn3�W�/��.I��I>��{�� wQ�����a�̝�($9R�15��_��
S!`.���*�=-)�s��ζ�n��P	W�q;�E�>��M͆�Kr�����WV��?�%��p3��,�n��F��־���Z:6h��;�+���	JNW���j�,݅�M�W2��s�"��9��~�|�AR?ai�����X��4m��~�L3ލyN{cA�1*�"���Y�����^�|�aNχ�gV��|� ��I�t�a� =�5��Ʌ��H�;�ZS�J��i�E��$:�W��d�.��71�-� �1�mI �[��S�V���l�=�W�J�wB܃���nm�se�z�x��H�K�P5+"wCQ�J�ji�t��]�k۷9�1q(3�1�t8�B�F� ���T��+s�pdb�f<Mm���������m��{/دW�s2���SLa�WY�,���؄��T�f1���������칉�g�a�VEa�{W�e�	�B*������-��Ie��bg�o��r�����b�5+�!�I$ϸ���n����/?x CF��SI�@!�=��>[y�ѹ�\����K���R���޸ L0Ճ�5�*7�-&r�tNݷ�9�����é�	rn��$�ԭڴ]�jh|�����){Z&��Kx��j�IsP��Q�2�X>�!i>�N��"\x�����]�؞��@I���P�5�Sc���.8���u%�{��U?5^�7&�m�\@p��V� ��c�J�my�n�������oK���).�6� Fe4rjd�m���FT��o0�Ed�Yٴ��,�!��\W^g�zs$�鉦���{��U[��tlϤ�$M@LÏ��"���\9���fJ���}RA-	#�lе6{�"y�dk�C-8� 4d{�lQ�S�y���!Z�`ߌ�@誗OnP�pZ=�o��
X���gc�ڴ�B��m`u�	;�k��szS>�?VZ�5�r4 T�TD'���6�E�e� �4���w���t'��>A �@�ud_�ɵ�xO�q�2=�o:
��Xǐ�w*BSc�Ǘ�5@�� ���궼'��s�O�G�6��Ob�&��²����!0v�����Xջ�nܠ5`p$ò��ށ�x�ygk����P4���gW!�CF{��������P���3^�8��(�7� �`��zg��E9�6���"=��b4�
���\9	�(���^$�8!�,��dߔ���������m(۳����P�C�����E�Ϲ�B-�8iO#����S��*F<�WR���?[Tx��a,?��N*SZ?a���g�\X�bx��w��]�M	a���S3P��~��0T_���עb��Kw���y��{��U,�/�
g5���'s6"�+ґ��@��#��c?���u�?�s��H0�2&��W~���9:��a�B��eX��?�N�����M��"+~V,��'l5r����b�X�4_�}�! �1{DL2�ML���Pe���4��	�6v�ʷ~��~����Lк�X����T��d��%�q��@0�n��j��>�&X�5�"v�Ro���;��*�k��f�46`j�On�~C?�d��gԑ�vw�E1M�i�#8r��p2NF�r��ZOk���`t���?�H�
�d+]X��FQL`f̷0}�~%�W�V�ӫa�0�����0�Sl��<]MB�(�c��Uu�
�+n���X5#�C�����?���4Z,Ҏ=Jؽ ���D�煿Ƀ/�b�.H?^��a�j��W��9�uOY�4��S�t0�MK#T�7¸-�Ay�:5��1��֩4t��)�� ��߂�r�<�ۂ�d�a���괚�T`g����-�߆z�U��/�J�ɲ��p5{g���ޖ�=�7�ډ�92�|b� ��ϥ��V���"�3^#>�To�H�����ݦ��ݞ|�Pq}�^�Z����v�������t�h�4��G�ڧ�I��*�Q]�\)��jſ ӄuE��Z.`֨h�p($��-�"v�<�f�K2�v7,�-��^���j+_�g!G��i���_��Yl�)���6_8�8F�ǒ�Zb�¿S�,x:��sE��n��G>�Z�I�����*i�1gn�1E7 �i�4��v�F�S�+��]\
!���ͯ̂]����.)�"��O�=3�;�8�l�I�Ś���V;���	�^o��JG�l������?N�B�[}�xv�'�Jc����Xt,��/9��7Bq�Ћ��."k��+5GY�d3o�ey�'g�飂�i�	�>�=���g��艄J�M����\�bL7&��m	`Յ��m��&���&�^Wu��a'R�l�>�&�����%Fy1Rc�O�c��<��� c�[�]��~{�٭���~�mAʇ���{��x�5�H�| 2�{q}\��<`�����^�P[n�XcG4.4�f�:*�c�SNJ%�;�ZZIwzu����'m?��bb7�>��U�(�_Ҫ�I�����l�ӄ���j{�~�u�h�7�Rx1�=yӂ����Z_/%L�8@�5���oO*��ϐ5��E�U�c�p�܃&�j8=�*�"�gQ�Z��[�At*$Ǔ%�\�Qy�f���;��yD�c�ۈV�lى�����t�0���ʌ�Ca��Wb���������Gb�3���{
�G���^*C�h���4_���=�Dt���}��߆ϵ��M��-���Y6F\=^�P�|��!��B!홣�u5@w�c�Z�yr{7V��vQk�r��F.�����X;_����	�n�#�*b�Б�RSʵ�)�KT�����\�:)Kf�
0��@٪8�JP8M�~�� |e����l� ��s���k��A&0󘙟u6=�'�eo��n��:YQ�ĿJ�eZ���S����c%aQQ�w�7���{ֳUC��Vk�X�R�"�á��0E� ��,�����2k>���1��z�x�Z;,� 0~�O,v�m�oߗ����|�$ �G�K��[���j.�YG�5*e�����-1���$����R�\#��E����;&$b�8���{�NMv�`��$*�0sAk@���L8"G�.�WM�&�s_�u��@���z��r�x�CT�>����e��D�H�5�=L�uDOTQ���%��2��3�c1�ر�A�ԋ���&�K�J�����x���+�i���1:��K�_�5L^��f�fMX�����<������)�%O�B��E�/�M���)3��6y �d��a_��R!1�C�g%F�G1��\\ݳ�k��Tt8���6T�ě蠒)�oU����&Rr��������k"#��"�}]�*r
޳d϶�w�PxG���q�a�C��_і�[~ן�7�N�~���>Lu�g�ͤ"G�C�+��6|]7j�SB}ɍ�븅���)w�[��/���Ř�s�5ז�$�O�$,�*?Z��/ �&����;_8��xt_=JÆ�\;t13�*��8�xC�k���XM�8`�n������?���ϐO[wG�=��هDJMK�$�Ա��+���cQ���A^��"~8PP�}"�O<Va�}~�x(R�v!՛d/�y/�����s=��7��q_PU�=ۛT񖎦��ܽb��� ���̠���p����I�����IU��^rq���GwG1�E٘":v��R��?M���xJk���������Yiedwh�X�a��y�M�F�U���s��]��Y��I��ʼ��w��_l���5�D�͵Eu�T*���C��LIH����p3�[L�4LCަ.}���h5�S�K0�w:�ѭ��~#~� 
de�.3,���7��F^������z� �z&��~O"K�����m��S�O� �A����;`g�Q�>S���b��NK�y��62)�����\�GvA/{�_���J{�6���&�,/�����i���K��i�!��-,V���I�/%⸺]
�8�;/�5�D�z"�G%�����L��7���b\��W��B	V�́�c]��K�U"3��Z�5�;4��x�^I�z�A3����*~��سk���iѺ��2V٥<�[���%U�g
y���J-п�D�[w�P��d=`h�&���<�k� B%��.��!W�Q�����M�asHj��V�'����4� saqт�ƅ�Z��m�'��9*�)c��#����LP1'��M��N�}��4� ���}��"h�S�1�a�=��b�T}�F\��nXO}Dhj���Ѩ�̺�1s4�=j������H;�0��\>s�7�`뱊��J�p��M�j��>.zې@�<!�ƃ#���"�O�~x�_��w���qj���|XwRv2�Vǵ��_��W�E���8 fzp�5�{R�'�����.�z�h���f���+�)��o��Qm��ϖf	GJ��
��|]tq�v�T~_�g+�vz�k܊/�>�g�!h֟ſ��1����S(��o�h���2A'P�Iʩ��~a�������>f }E��\8]���������1���IB���e6�)���d���������**�����K���P�B?�5��`E�8J���6�h�gO�X�5c襗�eBu��N��r)m2�ǁVY�}L��q�Bx�w�?k�Sj��ס&DJ��L�i+��gy�T���#�dD�
���$�-�er����!�%1�W�+�q��m1���<HW�[�rmc�g�>D�Ǆ�4�4��A@��R^�V�qJ.��p�ɀ/�t,�!	<G�#u�I����}ʼ�Q���M���]�����Eq���de��y���Ң��ιXU�5��b��B���P�a�wF��`nF�+�a�%�o���Fu���W;5�!�pdq���ݿq�(��T��5�.GTBBZ�W�x-��T��\d���m��Zsd�rNu�_?ƃd@vCx���Zkģ:y�vj7a�N��ُ�Z%��UMMs��2��\x߶=b�RT��
;�W�T�)��X�\A
��צ{�<,����$&l<ƾT�щ�)�B8x�	xUq;j#KE&3ĝ��˖x2��������,"�X/GRj��og��%bp��Mv~ۤ��7�i�zg|�m�t&�ц�)��/}&�p�箹�
:
Ѥ�Ǹ��&�l�>ŕ7NZ5�݄�!���ˉ���֭W%̅�'-sL.�����;����'��P�.�Z?��&���	ŭbiWI��V	��"sj���3����G�p�=�6��8��?�L+o}�}�g6=�o:���ti�<["2Zc��N2������G*}�:Iڠ���2����i"�����I i�};��d��l�<v?���ٕ�!�og�
�n8��W�:���-�Wr��d�J�a�/�l~���Ll�=���rz
��c)
,T��UWr��%�`O���Cz=3TCڸ&��Ҿcn�Q���{��
%
v&S}�E���!�:�oC�9=o� �	���@w_y�}�g�e�þ�:�T�Y&�V����Z�� �5�jlW����g�H̋j����Wq�& ���C��,�L���B�3�����F��W��;�9����&�a+*����>��&)��jP뤼��.�Ip���H��6��F���	S�Pa�e�
����D�U+[+�Gc��$�gu�3^�`�J�>c!K��1�t#s"�om�/Ă-^U�<��p`�q�,��aK���LJ����n��U�
E�_�K���Kcϗ���ƱN��T�|�?:j�|�Z��ۛ	@:.��!y�a&y�Ȁk�f���̈�0�J�_�C����p�E�O��F$Q��\*G@�)$�`�% vAf��Ibw���.Kp�����j����z�澝��E.�'�,'�Q�m�R�����r��%'�꽭TA��sr c��,�6��)��`�Rq��n��G�����&��j�12����QM��B���[����B�eJ�b���U��Uy����s�RBN"�+�}.��}߰��(�B|P/��u���)���#��F�S1�ړ�5�ZT*h���e}�3��b�%�=Ƌ�;��,�}u��_+9K1���h�ߩ���.rOA|+w�5�l����n���@m�r���9Ŗ��!�l���Q��bg >%a�A]�Sf�H�?���t`0��U���_�Yz���`�Zӳ���OB�w8q��Q��e"�� ���M�8�����nۇ��V�!d%c��x��Y��(�D�O�U�_����);�γ�F�H���+��$|l����*H4�^�)�y �K.���D6���̻҄��6����i���~+n#_^���Je>؀�z_(b9ح�.3)����"�c[�+f�@���>"�T�ȧ�����H��h_��/$	�����b�v�\�7lf�}�ņ �b弡Hf���K~���K�B�������1�ն�ħ�b�o�(G����pu#������Y�'�f�@DTiڤ�4;[@� ��E�����p����L�({BH�t� �xU�݂� $�n��2F�}�J��ܑm9ڌ¯.^�~Me�@+(U��g�F�2��X}�W5�O?(�5g�>&�^I�3�?�T�]�Rla���,Bq�3��wp��"h$=Ac�8|y=*����|Զ� ���%���Fۗ@%�7�)���Ѿ���H�[��H��`�L��|Gţv���|���)�^&�w�<E��|�D4`s8eH���pX}�'�7& $�ĒQ����(��;3о�sq�Ȱ���$d,AF݊H���jpsE�X=,�o3%���F�B�����	��ݔ�$�Azg�l���&ͻ���fZ�j<��'%��]��q?o�vͦw͕0i���y����߹��"��.��r� h�r\�;3������_�>i$���Ό��Rқ��u�b�3��;���5��ÏV|֢���(i"d=.q�e���>�/����u���#Hy���RH�)����9�3�>I�<�&�8҆Q�0��W��~��`}��!O/89�)TSr�@��3N���N��6��J_>�>=����1�G9������570��c��1���̐3־<c�-�V��c>���E��1���7}�r�7m�/�t6��Xox3&�l[YڑC�/�����SҲ����)���c��_
�o�7@�xCR6�O��RC��[���#�u�O��*<���_�C?�T�w5��Vc��|�n?�4M��
�6��L@J��JU�5���1�8����y��2��Y/��������TYA���lC�-0������)X��5��`���0�\"�9Db	K�} ���*�xz�|�����҉Y���P�cd�$)�̗��������%~ ��޹l�N{#n��P[D�l7FnG��~���<y���jB�(����3$W��W�C'GmENw�HN����bȸ!��cR$�f�A��W�`���~��8U�e*�&v ��� 9A.���V��Ͻ��5��������E�qxW�����3�bz���	H���ҫ�ÿ�����f����D2��`�`�"G�A� `W_�tO�P\zD��PI9^k &��D��!OK���3:rI�D�પr��C�
i�����?�:�K��F;&��l(�ϴ.��og�Uu�BW��
"d	0�(fϻ�/:z�	���6M�����!xeS���Qڀ"n��|a����BUʛ;�n��3a�
�v�Ư��>ƵYA1�q�5�L��~[f���Coc��T�r�bO�z�h�ۛ8x�pE�%Z����o��0��~�#XS)���B�<�ɩBܼ}}z�3���3��
>���-qt�,|��AQ"KXo�G�������]�Gv�c�|�?W�!�%������m��H��y]n���F����B�bV��U;}��N	}��Aⱐ������qE�肬�x�K�+4���$�0�*��3y15���!���s�(K�@�"\z<�Y�Nx�[LP�;�2.�@X��}�q���y��esvҸeK�����3�:��g��߮�����`��x�PM]��Ç�Dq�&�Ɔ&��ѓ$S;G医`tB�4�v�%�o	(iOcJ^q����q��\w?�ʛ��$�y+M�X"�9s#��uf�x�4^�R�ݏ���3�#����\����牥��<9Vֻ��G�Bơ�h��J�C��Pcc�>~;;���)g��9��!8�c�|��^�86�b��)�9)%'bz&�v�V��L~�������L^�'"Ő�u��^Լ�+�k�i�|���9d_��/�혊G���2�����n8	��௤���3���k���2�G�۶��^����n_�����O�Ϻ��3��A�{�`�o�pq[3+lacA['.ge�Y��q�VZ'4QPZّK0aq�"O-9��8#�T�CF�V�P�+^߱��ԍ�	p?|���+�' �������x�������d�K�����X3���$��)�M8��U �B�!�+�"'4H��IIӃ%���u��6�9-a����2}����T������
i�����ܜͻb�;JE�����������N�4>Ҍ�9%�}I�rhm��x��)��a�;<�Wz{����]�e�?�{k�r]2�Xy��IYO�KL��	��_�p%�OQl���+�\ ��������		�'Y�Vt&�DO�H�<�<�~r�+劲��ע�"����g�D^�����m7'����r�e:\HZ�j�*��^S��V�:���-#6�7�8@Lg��D�SꓜD�Y0@�y��s�oo�U:v�����������z�@�(���v��bwS�
�h����z�8�3*���K7��Z �C�e!Z0� �&�X��1-S��g�OI!�o��į�� �$��b�qTk�7b�y,�	��c��c�Z}�Ug���	"�8CCǿ��K&���IZ�.�
����"�N��ܣ�NG��p������D=�ō3f��j3�
K#ﾕ(u��pU!G�vH�̽���E��g��~��xao(������R�K�VH�'^1Us�Moj����f<��y��7�$u_��C�V�׊���]�JD|ZWժ��P����䘺f���/����{�͌w�>:����"&��Z��nO�B�q�)��� ?�v|��e�d�|ӳn�2o�I�sn�hC������du�Q��w�eقQb�������t8Ӣ�u�Tmr1�ʟj����0�Sr�$������1O��O���3лUŮ��&̭�
z�G�(8J�?�wb�F:І
�چ�t��(8m�=��v�U|ʺuD.�Έ/�l��}h&w%,�̭z��`�m{��$��(@^n����ND��)�
�>p4�d4^�@��-��+�2�T��{�����N�N;VKXu,�e,���P6�m�Z��i�MXr'�
����"A�w�'��}+J��6$3M��o�,9/!����+����*�ڜၜ����&@�5p�p���l��+`��|����4 �a�#@ƷqT����%	�	h.�RS�M�X['p����r�$C������!�u�i�h=[7�9;-�֭Swy�t�$Q�iY�G�Ӂ�y+�s�}�v�q|9m\������|/W�cd��f�
����mj����/�4�}+�M��>AYs���B���?�Z��.�z����F7�*_/M��Gl` Z�(HP`8�s�L�������krA.�$��n4��<���*�b����_Y�կm��@�/W6n�y5���=�y��w!��gЇ���H-I3����	��f��XQz��Nʇ��-����V�P�%�9�Sl�lY��`1��� ��L9�vL����aSg�p�,j<(.#k!��XJ}�:
+����P64�'E��D%��X���m��2������pǌ԰���\�W����Zl��#`o�N��0�z>zBn;�!(��V�x�Z�_�.�1�]r��yxP���D�v�h*���I�^���8]�!Q� pls�o��ɊA>5a�����4�h�~��
�z{��]�pe���l��=�<�V'����jդ�w�׍N��a5pwy�5�p�\a��0�cp��fA8�ւ"�bt�j���^�M�������P� �����s��KM��YQXW��'lN>��Mi	�s���:!{.6J��Fz�<���:k�"d�m�g�wfDE���e>�U��ii�aǹ�2���x���j�|�!�i��洃��:��
lK��hZO�M�v�%=$A�Ӳ�&B�#૚�Ku ��|鼨C7v�L��X$~�i�� � ��,q�V-�7�d}�q�.�M>�`�Dx��C�a�?;�7�Xv�#{y'�I�G2����������\^��ު �'$�j��W��le�L1h#s/�U�T���y���P~�{��"���p�(3I�v����cd����ǧ��������4R���/���ura��R��!^\��]�Ŋ����WD���.�I���qN������`��H#����(X��\�%��7�����m���fb&4 �Bi��;Uan[����Jk�m��9�ݘo��V�]���l�,E����Wkݕ�_m���Z�P/#Ӗ��K�z=�}�;`R���+��~Ys�[��8��Ȩ86�pK9=dn��y�k��h����Sk�3Lƥ�o�8�Mfoה_�*��֓������X����4@vO���g>��!;}h6]W��X�9A����͡ĹP� Ћ��`�Ed�)ai�����������(G���PT���Yϔ;�>Ԩ9��HJ���֌��Y3&~[�k�>��L���|},K�*{�|�����j�a�}㊮�B�u �k���C�^���e��B
=-�<��S*Y� c���0��֖��e�$�;�Ê=d���"yZ���;��;\��-D��H����v��<IѸ��'��6V���^R������yȒy��Iv��o���SX3�����K���]�P)�-�҇�B�M�Ě���p� j��C��5��͠B]�){wMc��2��d��=@��pqY�����Z�,\�|�u�;��E��juP���:k����� ��s���7+����	B�G8x=�zI��tzV��9v���S���@*H��+D���0�XB�k��gei�X�"-�xxu��p��
w����v	o�H�4��!	���/�gb�����I��wqzn�j<�y%���*�� C׸$V�<+�K��L���_8���y��	%�B�{��kL�_�SK%Z&�6���EK�#8%��/�V��]:��i�-#��!���뎤/�^'�-ՎI:�>�MlF�KȨ��Ш}�L���jH��f
H�3���ˣ%nC�#m��0�J�q�_|����0),�k��.D(�b�5m8�{a����qh�� �7- �iL2�0��5`'����f��2�@��΍�?�n�'9�
h
�4�Y*�W_�UΡ��m(zr�>��M��d��*ûWS���|2�hԄ0>L��S���?��3�7�&}�����%#xś��`��@��V)t���F�x��Sm(mn#Y���gM�p:s�~�K҂��P���d�}�[->�N��c-���������Nm]�Ŷ?��Oq��+�=�{d�8����-[V����m����f9�X[������+v�?U�γguu<��8hP@T|�{c�����3���p�=������=mՖ���s�mlt�N�B�h��������cG�����^�i�TWT�\��`k�CA�c|���F���h��K�1��B�gi����2sQ��)�ir�Y����`�h���ĵ������b��N��h�'tU�W���g[�̾�1�ϸ��#7ǣ��5tSL�������x������A��EpJ��Y�F��i��.��D�(xPG��i�.�D��f/{��S色h	�*h)@T:��{�w�/JH��t7�D��(�J�{��U�j8�q����Ƽ���1��䔀h��-�O}��B��Bh�v�I)Ư�5��]�bZ���`��1��Gv����)���Jf0��I�"]��O$�7�����y{����Rj�V�㖎�60h�iem>
MT���V��zir������dA$�C!Y��&�Pu&��&I��׎�Y�<���;S�;�V���8C_���i��)�����c]���~�C~�ůƔ�yb&OL�ݣL����L^ܼ\����{���F�o8�P�����F������}D���<g�=�{��z��q!ͩ�B'L�B�B�Vb�� g�N��y&`���9�mHJ���ڒ�)�#(�=�5~�����U�����d��q�f2���k�L���U�=�D}Aڳi��C9�(��k3"mC~i*CD}pAI��E�8C�`G�T|�
z*5Pm�@��0k�q2P~^Aa��ٕ	V޻x
)-	n؛�����K���"� �I�g�w&7p<��e�:�a�rZn��'b�;P��aҙ�W��N5x���SI�.�K�����\0���5����SD���;6G�2�̞�)�䋙��"p�4/j��pq�Y ��`Ɇ�ɣ��>d	��0s<�{ˈm'�縣h���iv��&�q{.�A��.�v'-'P�.� �Cm�c�E��r�OLPԻ����������DN���<G�K���9�:(ν׊��v�b��j�����iG�h�Ũb"�I� �M]�nM�p�~���-��sg.���;���Yl��4/��n�y�vNE��OKH��#�ۘ��O)����:;��F?���#);ӿ��@�&ױ��q���f8����7Qy��U��ʲ���@�+�������bd�9��P�2����uh�j5���a������A]M=�3����U�C�� ꤆��r�0�wb$G����?y�4`�n�*����w0�>J®p��A�z)���gT�J��B��T�f�6K��",�u	ּ6N�
(K��z���
;�@����0���R�q��0/0��?������Ό��a�"`_�xU�t����:	:PaV����@���!��>�:�1�_e�B` ��g��f�R��z�`q���f�	��o�̖�O��U�R֒�w����:k�a���x�c�=���aRΝ�FEn õ��7����t3�� oդX�ˑ�Qg6��&lo�.4���|V��!���sZo��"��&��uB�:��n���6:� ��`�2k�S�n� Z����Z8�j\�E� z����--�6��)�g,6	_u]���D�"6��O��0G�����UX�����#���f�b�b�����q�N������+�\�����0�ԪBO]c�֣3�1D�.t>Q��\��z׍u�\w���1�(�w@�����t���������8dJ>�P=�
�f���?4���!��	
�P��Je�^���h�)�\4�-(�@fLW�#��!_�J��z�8@�<vu8��Jj��M<Ku�"x�&l�ϭf��-�3�m�>�����z��w�s��H������lϕ�䜞o���yM�Ј;��^v����c 	wM��#.ʦW��M	�W�r�gpPР)PU��K�1��妧���msи(��2f� M���A��-�+�I����~ӆA��F������bM��7�$��I�j�鑳��Dߒ���v4U�	���O�����"j���D]�h�r+-~�T��*�Ci���:֬�~���^�`�W����DU{!	� ��0��mM=V���	�G�kĔ�����q��ʑ�g�G<&d�=e�LUF���)}��7]���&�E:}/�8v����Ѩ��"�m�J�ʅ���i��U���k�u�&vU4�"~�A��?l|q�b���5�=��M��R�����?�5����,	^䃆�x��ev�	��,/���u�ϨS'��t�ye���d���}��c����}ڷ2�I����W�{J�9ȝ�~��q����V'�L����� Q�a&�*7ea� �1��.wGVd�pe>�x�n-7��ͮ�T��U�pg�ߌ������1��#5����0�ϧMͨ��G'$׮�`?~��QF��wp�:Ѿ�&ձ��н-;o�Sa4�mN7:o��Q�۷n�wl|��f1�[*7)�h�M"�%�?�s��ˤ:�Q�x���f�\w&�֜Cbm�ؔP�RȲ	���l/]����!��#�4f{����|�VYԛp)���b}2iPPJ�)B�h	4ND����Li;$��c%m-��<Y�w����ڇ<�u+;����v�7�׿�zT4F�$��gy>��W<�t�t�e��ϳ�8�g�y������~�B����5��A�p�P��*�NT�0�E�V!Q��X׶�H*���'i�
{�j������8G(��#�o�<ߋ-�(g�B�e������b����ŬT�lw��N�v�y+Bv|�y�l	4��?ߴ�EY�yޠ���?I���{)�F�ZP�SșMG`��g6U���J�0E�h�H�GQ�
��noȭ����uޣQe5���&=�7\��XѬ>p���L˽���7u���$a�<�A�4�F��Z�yO�3�Od�G�|�U?�!�!�2if"�]߇2C�����f�����21��E+Ȫ�F>�8ʆ��ȐB��/�T�#�"*�W����zd]I�p�2��GP$��/_,}<����IR,2��믎�����5�}g\Ò̽(�i��:�S&��w#k`F ����$��L�ykۭ�JnB�"j�e�R�j�9�/}h:̾�0����^�I��>�;�W��#���d^�����B��.�}����#�2E*��!W6���I�8��D�ו ���#*�$�n�qS�ɧGF`��W%2ڏ�Dq�.�(H�m[��Y�ے�t{�����n��pa��h�9A�Xx�Y����6H�&��wr9�,@H�<�(��-�����uMm�#���a�Ps9�t)iN����	�h��x��DJ��s���Խ/�� �0�E�,���ݢ��%z&^,���x5����j�
n|)��J;��C�BtS
��T�9@���
{E��Fk;=�2�������MP�3�,D�޻!����AWs�ð㊔,{ɨw�N���|�\�7�:㾛�a�/�:��lK�ip��+���7�:遠�G �B�Q��4�c���y�����ȇ�Ӈ�	�T�}f�SZxB����7$��56�-t�
��'+�
�����8�<_V��/�f:z:w�O����hC&�t������a؂)����~������Ⱃ$�7����GP������p#?��os�}Z`2���ܙfC�%�E KiS�ͬ�AO��\t>o��Z`D�t������A���ը:b�5��*/U�x1������K�O^ev���	x��>�d8[)���lL��fP��������O���'S�(zqi��Eӂi\%�F�{����8s~�@R7<�U�sz��*���޺�Z������YK$A��㋐�m~��mM�:gS�
W����>��`���acv��p������8K�(?Ά�r줉�}�&�JN�Oh��"\8w��mԎ_�d��v���^�o B(���K�~3���{�L�c�ޗz������Ͻ�(ʧ]�j�ޞ!3��:�am�v�{% �f�s#Y��>i�#o�eI;��+�u�w%À�E����C�KƋ��&Mx���6�+sC�Z�>t&�90U�:Z�H�n,4$��Rn9:�U���v�{;	�x?uߦ�����C}!p�뼺�(C��Y(+���2�<���;��+�L�q|bp�$�o��`�Q[r�B^�z��띾��}�E��`�
����銡��h.��eQX�7V��� -'�����BX�U�=��9�x�E=U"2ps�m�>i$䢢���K�xcUᝁ� �$��KZ|}i��v��G+��l@���2N�9�ts[�Jc_�!A�^����yjn=l{�D��c\�lS-t�'�Õx�W9g�&O��'Z��w;�Z�H[�[�n�P����1c̷�QzY� �ڭ�Hԏ}�С��&Sb�ߝ�4�D�h�0˞?�p�=?�&�^�c&�S�V�92�'�@w�-��^Zo�wxկw[��r����-'�⇐����8oA���#�3 �\d-��yry;�+�\����o�9t�'n� ���W3Jw��M�>��7��0��;o������.�q����˷� �`aa�$_)ri�O<�XKQj}_A�?[���:q&u�/2k*+��
(z��N�2�yF�##f�\�U�Y�O��e�
��:��r�Э���K�d���ue[ �D��t^0��Mj�l��h�/�f�4��X@�.U�sD���C� i)������4$�`��^������U���M�Q+_���N6׻8}iˡ�袺c�ӷ���æ��Z�z/\�x������E"�+vG����x��G {ҽ�3�k˧i�D{�FM�	G����3�Wo+CN��{��5*|b&�
~ڛ�}R� �����঳n��i������p�
�q�%9�� ̧�S6�����HQ���?�|��A���v���1�h��q�#uj2)� 2�Lε���P�YY��S�iK�><,�Q ��	Z=�Gx��%�x��}�-i�+޼������]���]���8N� (m�~�j������j组}OE	�?��/�� �.晰 z$�>����F۟���׳\��Ej�x�N���,��M�����!@{>����TXkE��BJ#m!g�h�@jb
ȳ�6�6e��F��d����>c$#��a���׺
�z{�;�0%bUlhTv�����z岩�FXia0L�wmu�mo�!�W�dW>p�����}:ZF�|�\*ç����p-]�o��z��[��|���}���;�iù��F�����hk_9����
�k!e�D~���c��@rK����랲��S�(	��Z�|:�S+=�c ���Y�q
s=�l3�T>���q���H�`���eT����N�����Օu���DA�>�V�̇f�R�	�}F�t���y)����w8c�e�4��=3F]�+g�o���J���J��`�dT">B�V�@�^B��<h��sh+U����Ð�fC������Z$������ߺҭ6hf*Td)�wB_t��^.ш{�e�����k���骸�8���ވw"zB&j���^g�EQg�s#�o˟d���Y�u`�{4��ͫ,]�e<L	g����P�5�o��bhr���6��~�v��y3��)��K�b��!zL����Yl�s@hh���$�vS��w��W��(�{�^7���Dx�|#]F�=�5k�6\쓠9��U�T�?6�zl���4A��?WL�{E�-��A��+�U��������t#/
� �wf��˧[�#}��s�^�	Z�;�
�<.h��'����ު^-J�t��&.�S	)䲂x�	�����yQ�\�X>�Hcw���=���6@ơ'�Y��]��`�ޞ�յzݣ)�aW%p�$��^k���=��6ƲB���X�݃�u��)���뷁?֩���S:m���v�@��!4���آ��>G`"��)�Tk]�D�jV5Wd�}y��wպ �ȟM�C�&��
�u%rK0A(�sXm�o(9�º{2�+[S���)�vN��tb��2ۊP�QR�@� ���!�a�vO�|�V�6�	�'s��W���&$H���𿷫v�;7����]=�|�R,xH�1i��1hнZ�q�in���3(�-K�'��S�~˞����g�&O����R&�@1�����B�����t���Q�V�oܻ{�3�^cI|V!H���H�`�!��>T� �}k4�Jaa�g�L{���F��g�6���] �$$��cXϯ�rR
�;r�S����֎�|��^�7(t��������O�`hA2�����^)~�Vh��/Dq�V���h�ϕ����t�y3�';�A�o����8.fJ5�"W#A��"{����x��oC-\Nl[���nHZٿ�Y�Ӗ<8�� %m^cs�5"5�,b\�a�:�Y(4�=��[�"�<��#J�[r���NU��u��NR{1ۮ����'o*�Nؽ(hb��5�d0���V�7�S�L�.oQ/Ƙ}���#��1�M���ރ��:����K䏱_5<��HC��dϘ�C)v��e�f�C�Ԓ�]�J�׃tj�	
���v2v�<zbmݚD6�#L�~k9���8*�4��c�^��ڠts�a֚hC�o��s�/�²�k���3G]��V�Oۙa .QISF��@���3�H��H%&�ܖw�Ȓ��p(ī����6�4J�(�Df":88s��9����iS�^����e�T����'�Bc׽O�sfQ�@7TB��r������?SA��n�C2�6�T�:w�*"�c=�d��p��N%	�+Th��F��d u(z�㶞�4,���1��7ߡ�eM4��ܥ���C�b���i����Iʮmd���hHӥ`y�v�l�� *�S6F���*}6!*��[�;^+��8�}t�~[�fY�tx�=�"`1��#)��!~nbu��q��5_�U(��h�y�6d3��╶R6�!���:����ucf5�F}>EV�A�-��,�8�}.Wo�+� �=)�+�.C�����x>\��t���z1�p��D��(��q�9MSre���1j�n=���6����Ӝ�6{��/���E-l��v[H��6�	�����N��Y�����@�%�tY�� ���v;alu�?�xc�Ӽ�*0�H�j�V�q��q^�!/���h|α?���"o�%�(Q1�o/MA9wi�4���p�ԙ�O���|�_�Nѳ����O�-2]�Խx3L9b��⧲�D�y9���:�1�1��D@][��"�&��� m�G�,ۂ�E�AKw���k"7=��嘑���11v�l�"��8��%�<Ty:t�����VC�3�����V�R{R8N�"C!��-��+�h����#��i��]�CgG!�q{]:��6���*���,��1x�ym;�ƳbxjB�6�o �V�����9 �G�8_������v#������{V��|���_�١�=�%+\�u� c���t�O//rV�<FMp��ԝX|���p<��}?�W�@����'��)�Ӄ�mჁ�d۰=���>�!R�����|>���j��������0�|�Ҵ5��y��e
*�͒�T�U(9b������b��#�*���B�ȓ�ݸt4��T����
}ۑ}��
.��X�E�w��?�Х�����X�C�Z�
q�uF��aq%��h��f�h�-�)ڗ����>���N��{7(u���+�M���v5��Ļ`c�q�m����2Uf١��ջax�y�6�d��%8{0��U�b,?e���H,x��mt�>I�7<D�a����!&��Ȯu�z\���9���
S���K�E��$%4��)��Ⱥc�����ֺ� ��L���3��@}�O�l+�HJ��b��4M����ݺ������ڡ�q�a��߬7���5/���9_��8��v�D���u���
���B��E�#y�#��ajf\�[��e�?�B�e�▂~�=����q�/����妓X4`�HA��;-\�)��l-W���3��eT��Lo֙4���Ŝ�x*����ߣϳ�e^g	K�)��a�ç��t&^�`���D^�ر�!�;F+������B�Cb	-'�EH��Gwδ-b�6��9�` \����@A�	�F�=@���[��KR*�v�����%1��r��c$B5�_}5�	����kjv�����|D5�-ܿl�|��D��{��O=����E���0|�S���S����CIJ�稩��4�䥾����ݯ+[�߯L�3e��oHI���x�[�
��`���E�a�bf�J�oGR ��X e�:� i�v4�8n���i!���>�/���с�E��Z�hJh��N26�!�n�&c1�f;�J�83���S9f� j��]ݹi� �Z�y�骡6��B��9[����[��o�D���H&�c`F���	!��Qb�y��߉r5L4�?]!�ݵ$������5\����\xO�#z�X-sR�e�0�Zo��PP�k��Y���3���su�p|�ݗ���n�<��'ᷱ�h�Q���!~nO
m�>\x��"���6�[n�Κ���_��,$e�!�8-g$O��Z�I��q0,�}�oxn�'�G��y���?LJ�n����鬔����I!�텱dõ��O��|b$�])n�p��\�Y�X�d�L�c�V��<�Z��WϜ(I/ͳ��%VD��5����4�>6	��f����σ��䫋p�jJSn��v�=(��9�*��a!�?v��Y�0䙴��e����~R3�;N�	�{�=H�4*�}�ӑ��]lE�.0,�.ͺ�og2z������td�!���\�vG� 1rϏb`�5Y�ށ2�u7*�&��hoF1wٮ=��D<��rk�p)��& �����{^c �.�i���;�>���ץ�g6%�q-o��7�s	d�-���}"Ow���j�R��X��m�K��卩
�Z�G͆X�X�H�w#4���I=D�bl�Ix⶛:JPf�HW�aH�aU�o���I3��il�Ò��!K<�QG%-����h�V��I|�NVt]Vf��w"p���zy�"��"�Y���@g��$O���)�b\[$�Z���S^�Wz���Em��&�.��G�Y��p��І�/lnrpBˉE�mn�`Kc\FЊ���CM<&����Q:E���]ѽ��;��44�NNˑ�0�Wy��f��	C)B��D����2γ�'\/t��N�������(%4��Sѯ���8�sIKS����Sm>;�rמT��'�jO9��o����#���kg�[.0a�7]+�l�L����G�ng�@�_(�@{ � ���d[W��7������XR��_����� 9|��O^o�'�^�=M	�d�гX�`7��*-ɹ�&v�\W�c�vMg�,���Z䄭�d[��J(Mh{}2�q�/�6b��xpu��:p��V���?�6�_Wz$h
	-�j� �����8���)�?0��7�H��Xl��I���Q�B�I77��d�g�F r?��@bv!g�)�a:$i!/��$��z�i�œY��5dA��:�̉�F��������n��4���s��>$W������м�~S�m���Cƿ��+�0c�]B�9���҇_i�{����\H����ؿe�5����2�[r8��(Ol�_��ګ�P�~k:ڦ��L�d�=s�[�t�L�@7����]s���3���ٺM{�z��Q�Ů�(�n o�T�\:�7t��XܔBu�e�f��Q�	�jt+�3	������hz�N���<d`���s�-;\|k��9��,�t@��!*��$�N�#obş� ,Y�z.*lu�*�F_z��i�^�r�s��Щ�A�ʀC�Dö�k2��o�t���E����Hz��.R����Kt�������.�[1�i'<��՜?HsM{�r�����Q`v&)�e�-B�J�2��MP�;[�࿗z����b�^���֊ҕ�<��L
O=��3,��c#W�dx~��J�l���-	�~�j���3���S������ee������`�;NKo�j
r:���ۉs"�8r)�ep��+�M�OC�+�s��H��kTA%x&<�VB�t��7V'��ݠ~�SUA�#f�s�L����D�����\ZX�2��H3އZ7q�a�J�{{� �w�	�v���#�C[t�k@�V��8�+��G�3��=���'[;ϩ�FI�8]ڂ	�ʵϵ�UfV"^Q{�����Ip��W��0��R"����3�A��>��Q/
�][����� ����`��e�S��M��|r�C���fk����x�����`�K��]��6���'MLhk��u�p'-R&6��v�,��;�&hj�!��u���jK�y�ۨ����Wj��n6�y�=W{��q�����RG�O��Q�+&@�/L_Ƞ[���o�fr�o����b`L���k�=��k�� 96ƚ���j���~��:U,�aAf�����CQ	2 �P��B"װ�
9a��z��Re'�ކ��(�6W��GO�����!�Q�V���EmM�ҺK�u�uʉC�Vf̤�j��#��x	Rz��s�P�BYg�u��Q��Xڕ���0�:֓�ɎM��.��AV����*M��������Q_�d)�~G	��"��P�\W�eo�"���7z�81���:�VKg��f�J�ɔI�N�����n��#����S���cz�L�LfEO�"�:��`D��$ۗ����"[�oۿ��Ƹh҂���ޡ���D�b� �ڱ^�*1�9�)�q��{��n���N�p���烆u(�F�9��ϼ��䨟Mr�# �>�}_�B
��Ha�!��VQs�I��w�]����DO�)J79��#
5BMn<+I6+�l����-�z{+��fL�j���6�KN�(�\���f�;�9) �Ό
q����8�Qo�{�Iӧ�
E��|�Ȏ
���� ����� ����$e���E����<�'����:�Ʉ~h�p�����¦I�ߟ+�s� ՚F���)Ѥ&�M�w�< (AB2a:�G���ƴ�ה/�*�x�gH��e�F��/ܯ]�8r"=��!UH(��aQ=KT�3P>�a�	L��3 �v���ͳʈ�Jgh�oPoH�i9L�4A��je'��)��?vXET�'�o~��C�3�|����N�kF���7=�h3�!8'T�i�f>�52߳���j� �I:��_-ĸb�g�M�V��'x�r��Y�ʄ'��<:��)K7��7����W& ��'*#@�9��_��[�qP���>Gp �,]W�	8��Q9Pr9��7ز�5�����%�s`��4�\H�$�<'�c���+�yN�)O��v<^(F�V	u��u�����ŲR?td���k6f:�i#�_�p��4#�ߴo�(��E�12�,�Qg"��D�bv.�)wǵ��c{��yJf��Nv�'Br����c���|E}�kћ��=��`��ܕ�QsjtPiJ�YGA���H�;���[����O�M�N���`N�Hn�75��T5��]�^onb�Ǡڊ���5�C��)õۭ}�%3��`�r_����̲#�t�94�ְQ/�L6g> 'D�]�^N����{�Z��˜H�ꂺ�I��'$�D����ݡL�'����j(�p�J��`U�i�N�Q�(_�a�iL�Ё��{9R����a��	k�`m��WՂ jPM��h]Ɔ��
c�ҵJ���<��|�&�9~�kpg��m��Q9��]k�I�0-�G��i8��o��O ����*��|-��V���J�x���ڽ�)��`(`2�ڕ�+枂f������-�d�5��\*T6����yW02	%��b�ϛ��E(�7uъO��|��;$�8^	�U���g��e�'�Ø9��K%�Y�K���˟�W@|,^H̛��#���- گ�3��S�<�ZO��?a����<U=]�n6V�Է��F��Q�8w�����O�Ϧ
���8�k�2�S�xu>fOd8t��CS�ժ=/�!����#�%8�0D�:�;ؐ��i�|z��	R���ﾠ�R߰�����ЯMI&�^��c�#���)�-]T����<0_d%}<�ݵ	gd��lVѧH��ɗ�n�0}��Zǔm,T�@���o�H0�4��sa�3�V�O�Y�l`I2�1��G׎�	�aX����	�O��V���ܶR����߿�B���.��!���	+���^0(��
̈́H�B^g�*{���:i��n�O֙�v`��wc�a!����H�=��T����#'9RG�6%��<ˆ��_�[�ASEj��׿����6f�ه��d��t3ƩTH�?I���t������q�T���fgf�`��Kk�C�0���*ߣg��Ȭ�~�]��<���
+#;υ�Tw{�BL����7t�T}��Z�c��Q@Do�nRK�Ù��f{K�8�B�c�1�6��9�:-	�q�:�FfF���_��5ě:>�X��i�Me���K��>�ֆ&�u�_U7|��k+P�쯎��E��.j��J���5Y"�u0��nCۓ�YR�~`U�+��\z�p
Hq{�� �]�ǴĚ1!|�S\<G�q�D�TO
Aڙ&w��Ȝ��;�+˼��Xڐ8)��=atDw{;?�W�Wu�����Ն��G�U9㞕��Мh�|N���u Oڞ�U/)��+!��y�lv۞$Z��7CF;�t�Yw�(K����U�t4�D�ȿ�so�o�h&�1Yn����ʝ1�b�Y�}k���܈V��x��֥�K�[��l�P�6Me8}���lh�(�dOU�~�����a���x�I��{q793��9G�F�Y������1�o�]�?r�6����O��n���5�x������Y�~~p�l���)��E���h�o�g-��g�n��V�%���3�{��O)f3�����L~������!B�f0�MF�����j�6I9"�Mk��ZC����zi3&�f�Hg�yL����ԕ���E��u�b�c�����vp�u��(Ց-K������5��r=�a��P�Q�ħ�gǜ���P0��p����Ȱ�Kj�]�9 �-_2&Q�Y�?��-<q�V��� �<q짣�b������>�^0�|�>���q�c��8\��w�֫�ؗ����2O��Pfl��6-%_~͋#M&3�O&��F��[�"G�W
n�>����7:f�ف��a��,�Ǵ��ӛ�Z���Bk E]�.�N�k�?�!w^�顀��P&$��?��>)��gyȽp�Ow��p@���E��ӈ��d�4Gt.?߅��$�R�������Uđ�8ɽ}x��Qp��n��D\.��TK׳�K=M�b95,�	YH����p�WkF\��+:��
_��Mo����Yd@_?B��T���C�j��$E��ڌ����;Ǻ�E����%h#�����-��3��@���'4���'O᭧(�B��p�
ځ~6ʡ�t>�8'�+fb�NC�}���\�%5�g��7HO���Ă:J�A�������SS��m�,xNe���<�*8n�S�ђ�uc*�q��w�rJH���%�� ���_���F h{�@��hgכ��|Ω`,F:��n�&�[��^�k�}�}y���{z�i���$�aM��R[M��4�MY��Bc������8
���j���X�GY� ��~+�nX�`�dzV�{�:�ݭU ��>ж��!���o�f�`5������p"�ͤ(�iy�R��ðge��u�a�p�Y�2��P�8��d��^X��򧠶�(~�����[��JZ&��(�[^�RAD��._�[�'k#�N���n*R�(�Wq��!�I��}l��@�,�LP}?*�·e鍔R���P�o�R��B��]#O�K#k6+z�]��)���{�#�J{mvn�Y��U =��:�� # :s��/� #V�#>z<�bk�`�Wb��ނ}��|{��BcP_*qޮ-�[�|�ɓe\�8�˻��Y�G�s��ⴥ��سǕ�����ŏ�٤PJcCG@JLs֙��Y���r�^�I��.af7j?"ܧp�=*-�H̛!�aD��s��`�$�2�߷�� e�apf���K�J��M��+��7��*����\ƶ�0�^cD,���?��>��s��ș����?����K��['�T�+���,�r_���c��]���.|=�:����&�DCG���>~�iu{��V��@TlGڄ��!h{<��5�������̮�p�q�ⷐ��#�V��S�IMWG؊�C��@�a������i��O���0D��O	��&�t��?�;�����޷Z��RաGȈ����~�~����:v5Уe~@t�;�K�w>���!cw�k� �Q�L��)�'���t59�j�kFq�I��U�ܐ�Na��o �ۛ0�?Ѿ��މ?���};^����
���Q��/��g0d��ڱ�S���O��݃�iS�I��]���d����wZ��=��	m��XT����x�\ճ�e�'F���&n��p�_��V<�l��1�i�j�i�W�5Ȫ�ѿ��0J�R벸0�k�[�
�ocZB��k�J�/�<�'�:�����`��1�&;CUHc~&ث+}rӪ�+��_���#��i�����-(��*����!�d:����.H,<��|�op ��5)"�|�L�1���:7���X�����4��*�Oc�*NL!�lpk���!�5ʹ�M�-�JcԿI82��/���Áu���fꩡ�veC�������	[M�����R��Ox��l���I��bp��|~9� �f�[�d'c�9q����4=`y�v��|;����1t+��u��FG�d���j��@���&����G�����Td�"|=��O�?������~p*�a�L4��J���ˎ�LO癮jb�[[�ן���؛�g���o�SZ�kY9�H��/:�̣�/ū�3jn&�=6��lE��|;w��O�mB�e���n��-����R=L�E���g�����o�_	]+��F�Y��ɬ��N�|��G~�y�ڊ��^Č3\�<;�4�Q!w��S��hw��-���#_{��$�O��h�����م5~kaH��mW�-�TH}I�QP4R�԰�L���m��b�)f�MD���N��)�-񻅸0G�GE7�;�� �N'�N(�~*R;U5�j�Q`�&x�?x��>2c%�B*��c�uQ�PƆl��z�v|��u����|���*�)����%#�?at����E��54J쏑�Q� ����\�����~w�K>��Ţ��X��up��=�U�x�XΛLݙ.6��q����(ic�@�jb7]����Q�UH�ԟ
���OV�>���N���z-���:�H%�[,����CcX~���
�o]��B��J���X.�.+p{���$>���5�LZ�;Z]g/L�l�v�~�7��!�7_	��~��}7��|���ȟ�~��+b�@�	����<����
��2�{���P� ������ώ�Ӎ�Tf���(Zȇ�K�4�l�������+[�9A�� �EPϸDcUЬV�z&]K��KW�lN:�w�w��^� ���F��i[/��E�w�a�Yު���������<<�Y�
��m�|�a"�>΋��w�s>؂JD[?�8�J-`h���j�V1&3� ��Ew��dR.���[\�9�)Չ����޸�6ǈ	*��q�	��R�IM`a������x q�;p10""������V��a����2� ���ߙ��ǎ�*l@+�@�����`;�r!��T�2	���=ѩ��c�V} �je��X�1�`4���)�3��c0b���ϢZ�[�jɉG����~��ޞ�+�i���`�Ƃ��UAg�P{�oa
M���`���pq����2��i�6j*�T��Ǡ�e��Ț[7E���)n����S=���,�{����`������0�I�}�$�!8"��a'��-�H
�\���0}
����8w�y�(�����8C9o<ȑ�wg(Ux�S(mK{�?3��B+��a���p����}R�E[(aW�q��|Ȭ�A
��ܨa2����8�u_J�NJ��S.���RA��Yl��d.T�j�6����6���>������t��U����;�r"ĺ?l�W/X��V�����Q-~����G��um��EB�po�1�r�ޱT�Ŀ����4u��� su,�����W�52f���h���B����e��R���$�79u�O�	'H?���N��Q�;� �!9��	�%O@��r�f��K6f ��/�#Lk�k��С��
�0�j�[����mo�R���p�~�O׳k?�pK����k�p��]�����c
�2`����C�R,{Xp�@�T1��
8_�갫��L�b+G�m�`��6�P���ac���!]��M q��,��d1-�)��\�m�n]Ӻt��}�ޗ��"3!p�ϻ��V��u����?4[龸�w��r�[>�5?��`�{5�)����Q��/�^�\ϳ���pGA1S
��q֢̮����XwZ�L��_Cr�Qt�{]~��!��Sr�aW��5�te]���ѥl���n����َFc��݅����!Ѩz�K܉b�ot�tӭ��K��Êhts^�Lmt�� ��@ ��F3�2�u��eܡA�E��CvK�6l���&���0=��]�k��Y
�fw~�g{�Y(ԫ�$�#�j��-xD�`cG�^��h�n>	����n�'���o�m�I���ô9�X�mo��/9E�v������^�������r����M���}_<���Ɋ
��**+T*�G���w�To՚����c�B��-^��p�q��k��1F�}��-��c��mY�X�Ae�uQ��nt�3�Z�Rv������y�SD�����HW��z}����%xrg�����`��ˠ��U�Q�~"��Oy*���)P~��+j�5��f���V����WW�[�Ԅg1����W!��t��4�.Ү�-_�< a4��8�a?&�w����FK�#f�Ę�[�\���~�������� ��cюi"J�hȴ��z{��rDڜ�r ����^*}h�q0��M������S�a-矞��|+;}�Zм�.=����6Rh�C���#������e���iX{8�8�;�R��X�x;���/��yNy�\�s��R�_ �@ �(��q��;e|��t��ջՍ�9��T�k.�šD�/��%����QA.��^�ۨ[�w��`&���b�E<.��PP�ϸ�n���H��g�
���i��kZh鯪�s[� �[����
��E*���t�s���h��[E�}+���'Z�mԅ��c��U�ұ-w����ݎ�\3�[�6���$�E�l�-9A��g�wA�h;d=a�|:�j�!DU����:�u�D� �˞��%��ֶ��Mղpw���
���Y8�E�Y�^D�� ����_j,�zΝ�I�nV����?<q�c��r���(HN�d�������|�=��_��jt׻����PW���ǫD�z�%D�E��+��U���Ԗ]>~P&Nc���^IB'�0%n�%�[z��m���� �e�+�蓕ǀD�꡶����s]:��C�E?Ҏ�D�e��}��`:�Ęf��/�G��k:f =�u�7fs�R��ܶ��đxx��7���@!�X�(��or#��=�1p�^�ْ�,�tJ����.���vK������o�h�1���x�Ճ7,cl����K�_�K�d�+Z��~�Z��\�C^7�g��a[��v�+4��,�"	���gN፠|�[�i�C������t����ʄZ��L,���(k��v�Q�)�Z6�W�|!x��JG' =77{�ϭ���kQ@�8���CkϏʗ�\����Ҧ�M��`[�45~r,1iTd�<�AF
�̞/�Ab2�(N��K��jS/Ċ��AG�K=��	�F�b��>Ü��M�b�� 7���7�K����}���Q����q�u�_�jQ no#�j�1)��G���T�2W�p�26!!�Z<���)�����p���'su�X��H��xW�F��8+���M�S�Zӣ�Z���(�o7�CjS�`9�(�7,�q&�."H-� 6�f��a����+^i-ݕ)�$��ʬ�e�-[��1&���Ǐi,|s&$,6Q����/=��d&�����lu���r��E�,i���gs� �a�� pf�6CTw�#{�(q���_��
��<������xm�Û�+��?��婰���d�(׸�Æ{9^mlXֆB�w/	+ה��!�U��t~ze�4K��-��f� �����ȱ�/�����C:�ڝ��t�}�y"J�y���<2�LUr����C��4�]��뜋�h���\����ݛ�k��������+�I�iMý���\l:��xh�P$:��ؚi�[���X)�e������c����*���}|RZ�N��4�ta��'Qт[5�FX�]��r������+n� 4����a���&�ѽ��/z(��9(�qveF��*2+e׵^�u~Y̶-DS��A@e�[_����D��Gh!bP��9��h�KK*���`7PU���פ�U��a6v�R�8�P�!�n�[��Uc�����&
Ÿ���E�oa7����~|��$�d�DKd�6@N�r����ϻ��U.ԯ����	��g�'"�-��lf�����JF��es�loNQo��/�o0
P	��)wMS=S\.ھ�] A2⓬d���q�������|5�K�8ݱ�����۱P�_b)3-������a�������^ɩe��(�mF2`�'������<џEI���4�!r�0���
�1i���]i�jnU���n��؄X[=�C���X���]��/�+�'Ł�l>�`x�}.5�Rv�[mIV�S�t�Z<��L,4��y�n�/k��#�&D	��.�k�ۇF���Z죏m��w�e�8~�r��Y�!fL{�5�Ii6���q���j;����l������nf��)��Ђ+���_�7Ԭݐ�ԤGom������b�� ��D��=�kT����Ip]��K)��M
��[&Р�rf ���|ݒj���ȮwK��D��j ��cL����Uy��� �n@��mw�Ppx��#Lj��*Q���P?x�u���T�(�;���i�57��*�V����c͜'oj��j���P��#�*`�z�e�u��x�o�ǀ�֘]��E�b˟3`&�	N����j/d��;|P�f~�UO�Z�)u-����
C��
!�����﬒z���#ۻx�ڕ�'���^�57g��j>�Р��x��t=l3sSh�7����KZ��wK���.� '+�K�Ce�.�+'>�W ��V��:=���z����L����>��g��� 2\;�#�:mO��#�!h���}�=������E+{�n�Ѐ{'΃��tC����\�[��`Ϭ��
�Y��lnbz�:�mT�H+�V�����9�	:�
�&�A������;R����C�*�$Q��
�]s��3���
�J�/��dl�
@x���!�Z}bm|�6�d�)Ҥ��v�܌��u_���u��4��1�@�Y=O��nD����wJ���k�3?G^�|�-%��'sdh� P'v"wd�����n�^�P�~��e��-��O"�q�=l�s�S��V�32IwAD���?�=>k>���[��͛�ZL�;g�^�$�&��Q��SE"T�]2kw�J����W����G��>����vR;̘�̢�1c�9(_�ع�����⃋L����X�h�����t���zWٸ���m�(�ٓ$ fץT94 �m*'������V����|ΐ���v��}�o��ά<?@�Uٜ�p�|�:j���Z,�X6r�@�d��:���_�[-S�O��)6y�'�3L[B�F��t�C/U*V_(Ƃ�� Y��q<�vX����G�wJ��5����h����BnH4��: �8�.Z��<�ۃ���ߐ��_#���-�7�96�B1z"�K�-S��./u�4�+�O+�<�ٰ$�*��#����4���mn7*JF����+���	�T�;������S�!qc��Q�?�T�q5G��9�G5kq� [ݶ⸴�1�}���ZAȎNyT� ;������Z�9�°�>�H2��FJ�u=H�L2XH�6��e&.G�}S��7 _� >Q3^{0UFr�N_D�y�T��F�~֎�)E8e��ɜ��C�@|�D��Pm�����8��� �N���B�
4��,M�g{Tc�J������������=���۽B�$:��FRx[����2�ԙwU����͙G��T� l��ıZ��F����G֚��sb�C��v��q_N�-�C���xQ:=�X�]�P�O�''����/���:Qib|�A>�����Aă��z�𚌳�A���1��)>Ǵqr��.��Wa*Yh��H�V���(ӓ�9�q�^0V^d��_@";F�j���p�0�g����س�A6]�YT�����!�S�I)��aV�t�eH&:��8|�Y1ы���V�B���,H[6��^�n#����>���-�~�&��L��Na�c>�j���E���\�!��W�ݓLQ����Ae'���&�����=`-Y}����k�䟰o��������Rş3}(�����6�y�{��a�]�8��������1̯)��)t���	�'�Дi7��î����H����t�q(�"��m�3:�l�"ua�+;�6���0;�/�o�` �+��g�!��o�W�FEQL��ʃs�j��@�i�O;~�h�C�X�/u:�Í���&�0�w���ů���ן�粩,��APG�kJ�ʔ��A�YR�5�)�����a�(�Q�g�kv܂��!Gtkuj���Fy�Kܾ�H�7r��cvԦ3�]â�?���ԃ����/�m6N��,s�a�"�h��L��Op�A7^����͛���э�{���g�����(����vc�D(���?2r����m.�!Q��_������_௷�]��3o���E��7üH�VI���)ʽ��@�l�ET�'o��:�8�o�� Diu�k{��ɪ�j.����6�1䢦�Ы�J6a�p�G���ssi�˚['�D��a㖊��c��ƅ�m�������?�q}`(�7q#�; V��r��-Ap�WU(�����..���Ճh1Thɬ�l��� �D�t%�H��ֿ�w���q_'�|�|��kaZ"x�ܠ��J^�)�E	q��C��$m��7IU���Q�^;/S�\Y�\�p]e��^+���!��:'��o�Ϗ$Fj����4>i���h���Ҋ�}��Ŧ�91PW��#CyH`ڬt�%kF�O���e�V�6��� �Q�љ����w�����Q�he�x	8��`f+���4j�k��I5�^��I;��d�dE1�a�#�_��C���T6u&�n�z�7*ɚ�Lyē��x���T����U$��!\����(c��|v7��bNTљAr��2�~K�id��C�r]�Q�����*��j�~��7M���m"(+U� ����v�MƇ5�W�\}X���
e�HR�m����K���A� �煮Du[$�5B�8�A�l[��,��G���(��W0���k��<�����d� �hOec�'䲄j�Q%�u2�˱#�����a�.jf����'�Ցecf���6�~��� -����d��5�S!�+�Eֶ��Ǐ]췁�wݟ�)�9����~��,��� ;�}A�����&��~%m]Y:äJ�I(��a���T��˒����Q������v��#c`D�o	����8 ٺ�R}������Ow �p0+s�.	PJ���y��.�������������QIT�G}/G����qqA�MI�uC*PY	�
G#7 ��ƌ�d?��%bu����8��7�n�!�b�ʥ�YΊ �jC�
����O�&�
F�67��w�B�3��|�<;�O;e�RS���62.�m�;j�8Ǹ���i�������׍/�E�u���qfc�B��ĚP&�F@�S6��S(��T���!���#t'pM|
�B0�\�KC��F=��֬�N�3؀�@".�9Ac$S�~(���Eg��ݸo���66�Md(����|hQ �6eEt�^y&�ù�%|�`���Ń`��k~x(fSQ���F������\[��O�]�/ҕ����Cx� jx�MH��k|�df/NL���H0�XL ;�����	}�T�����j� Va���y+y��{�I�.(A���h�+����1s�������x m$Z����͠���G�m.-����N��i�?�Р|����)�5��p��C�"�j���)���&p�%j'�����g8pS�������4�V ��'ݞVH�z�L.��^_����I�� %�uJ���τP���_�XFw��BT��eGMb�$�k��\=�=q���t��u/�G챔�' ,Lr�'C���3,��"Y��q]��|_K�t��4y�b��:�~L�)��M�)���6�W�6t��9�⽹��n8�y��c�3���͡���-�J�$(MesH>���-����mF.�9�j���{F�Uү�}�y�(V���`�_W��)M-�āD��s*��@�hzp�$�P�}�u0n�\���e���Hcb
(�HR�)�aBr��v&��Ă��W�R���3��T����uE%�b�?1� ۻ��)�7����������W�{�����n=�y�b**+��X[o4����܎�M�t�Q��l�}O!�3(�wcY�4o��3��1pc{j���������;�T�=�Gf�OH2M���/�O�mY֢�^c!�&��dj�v5֒p!1D(n�'�\����v�GN�qb�����0��}_���V��Zrm�1F��b�9%� ,F�E����jXq�^�ĩ�,���3Z�(4Rے�k�%+��[������v���W2�J���	z���|�*�4��7k8j��欥�uQ�Yݣn}�1�/��-\_�}+F+�|:UdB0�����}�l�;B�k;NlZ�-\�=���s�D�_U{	i��ٿ*:U���v�Ng#Η8M��x�Z.|�J!�;�*厰 �ru�X]ޛ�Y��M�3��T�E8JitE�M:H��@l����-tL��B����i��t�?�*6���ڞ2*��'��Lb,����[���Y"��B�p���E�5�¡Ia7���/�zA��z�a�A��`�;}\�z�Ֆvkt�B�o����׈4�5��$�pO���wQ�&s�0�K��	���\>�F�E��쓑��1g��-�>����J�P���!��OKŅi�+��HfGTnl;��;�eA �<��S%-�*�qvU^$,�C�	��n]�6����9�{׶�%��^���<})�Y��O��`�y%�o~i�@?��&���D�f��rAP>vo>+	�]�j7@��$$Y�"~Q1�w����mk����v��E�K�+�ws@��b�I�U|��33�ɻ��I�>�Uз.� <�t���0�ݦ�iř�ͼ��gt�8l��D�L|5`�>�wh ��U�u�"�$�����.LWH�s�6n�p=�x�~�ݍ����!�MHf ޶��RRۑ*!��o:B��l�����(�F��e�=i��Y�����8dŦkU�����1:�{�mڤ/S5�n����LYa�I��d�P�ٯv���nޕ������T܀[�k��'鞯�q��)wZ�L5)�f�fp�ю.T��in�?�Vz�L�~b㒩eQ[�M'�wy����A�^���li�����az�_#��mi��B}���"���;��d�n!�����k�^+�륚B���S��ڼ��%[�:S��X5�[�dϺ��#�:%�]6}ni�Ȋݔ�&ki�����s�����Kxb�7�Zc�[?Y�d$�Y�>���&��&��Bnb�(�����r�:�2�\��G�a=�J��n�wt��W�t�uY���C�V��s(2�%]���RL��hY�oK��u#?��ts�����%Q8�|��WHD���W�������Bd����-oLӻۻ�@�� <ŀ	F�����0��P����YW����m��SΕ��%��5	�,FL%�Dh�8OW��juֲ�V�i��|�פ��
�6/��f����K���%B��ۄ~�9:��]�4�?V�X�c�I�]`���Y?A��]�������:����T���Nao�`��2f>4��X��0"ϔJ��/;67��G�5rõpଢNۈ��z�.T�3���)����
L�y@_I�0Opn�׹ްh�t7{+'�U�׾E��������8F�H�=t���^d}%Wӷ�U�2��F��\p)���ޥb�of�w5�f������;	j2x�@f���V1�M��l<�OV�Gl@��FSbW��Y�/d۫��Ą^�R5!�₰�)�D�~���;�c��_[�h*(8�^�*�y�v=S�U�_OH�'?��-0S�~晳�י��
z2+������ȑ ?�æ_Ф�p���z��P�q���[KS7 &��.�1���	��{J._ݝ!��m̀���z�1�HZ��f�赛$D�2��S%�Ԛ��+�X�'�&�WZS�**R�.�o~-�
JLzL~-W,|�.L��Wt�i��r�]`�I��<�G���E�,�!�Z�Z�k�Ӛ�p7{3f<$KF�#�!U����,(�
�D���6­wY�[�^��D��w���UـF|�&��c��0����8�Q�d���Dv�ʩ��@�,�ᇞ����ԡ��*��!c�����Nau۲&ð|�=7A��ɆK�����W�3�,�����.�" -�rC�"�"������l�#_�a�� ��+�Fݗ�:%�ą�i���E����� }�ԍ��9�D��[O�R��3O���'+\��X���ԽZ�.�>9�1g(��У�Z���0� �,閌5bhk�M�IQ0��b��j ��j>Ǌ��hX-����`���#�=b�A��m�OA�@|��풴�!�쎍����zg�+Շ��_}(c*��ȸG�� �>��G)�;�-v8_1(}�H{h�V����Ԍ4��];�-�Tgʨ��%��~�ד����p��������4����t�w���]���R�y�D�F��hA^k�u�fR�!_՜��dQ�	��ܓ�J� dYq�
��z��n���|�<�i��v�mX1{���^�� #��<Su0Zv�7�`�<3O�
U�f�x�hE�`��n������� �A+��TxK^1�bgȐ���3N��o�;0ԯ��Q�d�^!F�T.�9Yhx����C��G�>{�ߤ,�������vP������>�۬��{��o�{��́�L�I�T4�V�V��5�����h������*�)�Qg�	�vc���#ܫ�_�j]t�QD����<k��ֵ�,\/�;쭫�5���i�ψ�W�����J�,O8vw;ΐ%|9~ѽ�I���I��7����pm�޴�Z�S�e�V.�z�qQG�Y�������xR�]����h5kh>��p)ќ���t��ې��r�U���  ����}y1N\E�1�a���X�v)��Ŋ�85u����h���y�<[��1��c�e"9��tXn� ��s��m{*m��1s)�p��YSU�'8kN�B!�c�R����"���y�`���	p��t���f]�ɬ͘��Y���"�D�D�ތ�.y3�M�Y ��l4���S��U*�;�?+/K��蜯sP�BXAy��W� }�P��D�3�=�ʊ�l2+��dJ\>�5��8.�Y��@	_4Ҿi�6�3+�;3�_�ɳ��#m�"?����Tl��t�gB��]O���17�����>^�M��9Ȇ7����Y�H����NM�d���ք�c�
5�F�4����5_�w�Y�2����	h5th����Ez�������[h�L/�|�S�5V�}S̷�e-
���x� �CZ*���kx���S���G��Y�0 �^oBb�W���J��I)�Mi�[뫥[-Y0V�uF�׌ݪ�m���PJ�l]��,�|*`�	����+�ݪ��J���=��{��ч��R�Y���w��+K����@7e`����z�x�pXZ
�5p�8?�;��M�}�������k+����&�%��M��Nr�@�G3�8U�sU�,e���{�1>�Lt�G	,��)��6&�sr�9�-��٧�j6�:��J"��q>�L,����B6{w��U����ڕA���Ow�k�jj0�$u�����$���;�����I�|�e9�aP�<���h������j���R@��^���X�:��thT�a��Ql'�e=��W�߱xX�㩉������ڼ@�����L�z̄H�t:1*�}a&Ԑ�8chDo���,⌽ 't��.��R1�ht��j��x�"�eKX�LZ[t�#횏�����W���s��r+�V<�솽y�cg�!�Ƨί���i����)������Q?N�y�n4 �H��˿=@_�����Kd�L�d:3������'��x�����v)b��FŅ�<؜�غ�����u��1_��ލ�LJ�z������3ʙ8����?=M���O��AZ{{�Y"�����93.Q���Ü����L��^�W|��k%;SN�1��
1m ��̐YT�P��tu9�<k=���e�ϯ !ئMiC�����t��������{P�"�(L���'�Q&��Fh�$I̓H>{rnƭ�]�SY��-f�@�~{8�^�;]�伋��������8��� p�1�g/��c����nM�f���<�q;�V�;�%�+	􇽏m��wϮI� �At��YC��GJ�(;�Z��O��t�@���`3��í�:����$�����c�sP�nS���,�&��u*��՛�y���~�lX�����@�w¨qTP��e��+H���ϸ�*Th�A8�ڰ���V����`P�ռnq�g��y�"{�Q�j*�DFٌ�.�]!U���<�DndW�$1�'��	]'��9[�}JI&q�������µ�8�)�uTH��R_����	L/���0��
HC*S���Z���:Xv��A��)�3BՉ������"ID="^G�3��'hQr�����"m�S���	b��:ϐ�.����i�m��Ql��L�>zQ/<���H���������V�Gۋ|d�t_��e�[�&�C%�a} �I�юs��h{�r���y�����ѸmC����1��=@1�hmxlO�3K�Ư��y�ѯ�s�����C��{���]1���2�����8�����c&[����u%�O j��2����P�j�����e��(�U�K�S�ZT(����������ّ1y&}nˑ��0d@HVie��F̼�Q���}���"yݦ�Gf7�X�m0�N�6�ڌM=`���φ�����P��G�~�yW�GW,�7�O;DhE����N��=~�{�q�����E���\y��ǃ����Uo�Je��'�a���?��@�␷�kC���LML�S�H菝t�s�6��en�}��׭�j�)� ��y"P�c�.��������N��.F�:��p���#���0�%lrp�C�elT�HH�� ���Y0�rmu���yƻrk�EH�:��rA��^���,`�=�Io�k�<��ټ&�Xs�(��,�"�9$H��ي�į�/rvp��6�>b!�06�D���Q�$�����+�E��=~U5y���p#��ַ'�fTzI�4�{�kz�&�9�kV�&A��nw�Q��!�j���&��2ğ /�����:n�m	?�f�G\�=��2)N��S?����� ���dh�r�t�x?C�Fhkٯ�=<���	����N��eۓ��SV�o�{`7��]���ˊ��ǈÏ��>��B���.���9'eJ�^ B���F�r���^��Ȥ��3~W�Z�Y���7!U�o�E�ܔ�f_� �U�㔹m7F���Dc�	p|H� ��s?��@rq"���t��}���"���?���=����ޛ�幆C������i���
��<6O�4�����03����������&���]Z�!ݼ[��X�
7{'?���ݯ�q��&W������hm<�`�pO���P�R�@���N�EK�B}�>R�tKHT�dnM̈�_��W�XoI+֓t7���������U'l���(�gL�"k
��&�sN�?M���Jޫز�k����3Ox�
�,n�Z*Yq�|8���&����C�j�G�8*���53�c�'r~`T������"�A����iR8�����I���S}�/�.5�9�>��g�A1O!Sӥ�)ņ`4�r"p�����e�� \��j������U��DH��g"Cm��@�<%�y����xrv����D:��Cn�ȳ�-X$O&l��4�#��43���&��� 2S���^�.i�z��#�u�(�^�N��O\^���b�����VP�_+N��&�܅�w�Զl--;2*��F'ө��P��26�YY���+������+�;D�:ޱ߅��$���A���!��>ܷ�ke��u�2�vv���q� � ȗ�e�H����8�)�3�:*k�c��9�~5������hj`�lK���ѯ�b懛n�����X�
���"������{�F4�FU0�=yi����^P�Tڛ�z�[L��V��HG"y����Z�Ӈr7^V�K ��?��2��ب]'��@��M"mԕ�i�w�7Pת�kJ"UZ��&^�	����T�h��e��5��]ƥ4ȕ�L]{Y��eda�9�]�D��&7M�Zd.�b�$�Q��Ś�V%�
�V��rQ�H߫ܒ��5%6�{xFRˈ��\똃��sh�؇.'�A�+�b�<e�#6(l��,,~:�ƎG�N���4,���r�X���ь��ͤ�}�=�r0A��C3�ܮ�~\��:X�?]�3/�K�㘆(/����H,\�u��H gI5uJ�Q�^wV�ט�*�L4�I�~�U�xc��?�m!f�������S�e��sÂ�,_YA����� \WMŒ^���Pʣ|�*�>uz=��ɗ�թ���6�d�HB�T�-��:�8UB܁w$����-׿4;���c�.7���WZQ7�3�����>��̯,V�-������2������i����!�ͥ�4�=N��>�Du�{��e\K�w��������"����}W��3x��%�i+�l�o��_�5�=��eK	��Z,��WdB�t�
�?���Om�y���E���1��l|�t��>cD�E��G�ug,��Dt�TȮ$��
�Zr� ����B��%�e�xֆ��L(�7?�@�ޭd.�5�fڸԮ��42�t�v�-���?��`$ʠ�K�+�b��501	�� X�H3H���A�9�����^p?�/7���;�?�w���#�o{����q�C`eȹ։�P�U��V�5��ƴ2c�*�� ���P��:��@9�$�t����`Lwyy�ab�d��,2��nR=���Jr��h�T�+��-F}�o7PI1r�48ԣ�D˵�8Y�dwJ�i����/���a����L�aB�U[��������G$�^�$wIfCs���%��N�]bi;,����`��j����+�#l<>�T�|����(���A�\N��?�+.�A����n�^�?�>Ϛ��o��T�%���}|����;��J*�x�*�б&��o����n��J]����&qN��|	���t�n�1o���e_�K5��l~�`^d"s�p�s�0�g	x��h;�'U�o���1�����jBeҊ0��q�R{��O~!��W�������{7V*�g㨮fncDO��dc��^a�n����Y��4"�o���p����R4XP(��iSԺ��}���ߐX�֪���������)�GH'o�`0�,+TG�t˿g���L�Ś�p5�c{�;Sr�������pW���#����Y`*
�JFc��qJv����-������Q��H����6� v<ӛ	��3�ja+m�е�v�p�F�7@���Z@�$���S�r�^Ǫ���APlǄ��m�-|Un"���;�G�">��:W�$2i6K,��1y:�3�w����4����}�P�O����2��/�i�r�hu�9��۟3S����bQ:Ɓ����lTC���0�.�J��C�;��;�̾�;.BIq��oM.��N�u���f��!Ys?�-�b�g�-�!I�B�A>���� t.����Y���E1��h�d	\��y�fL�Λև:�rv�����@��l5�B}���kp��n	O��[Z���Y?���*o㞲e�V�C:��q2n���z/����\�����*��ہNNQ�-˄��C;Z; �#�c�ӕ��2�/!�֛	�{%zP��Ү���N8z�����G�ꓼ&�5��.L�;+,�n�?g��wH�3Q�؍3�=�(k3���d�f
��mʟ�'����.|Q���ay 9lTo����Q3���4ڋ�Ob'vn�����Y;��E��P>��@:+G�o�m���5�&�n
&��O�"�3�>)�VV��.(9<4�-�;�e´+i�?i� �	/�ã���(��d��N��h�7�p��d2C�OL�D}�tU.i������_�qr��-�[�p�sN�>��k*�����R!�f������j����s�����b��݊36�� ��M�ʡ@qy��Y((F�3Tx��5�)~T��7�=�P#��OkV�D�8aE�z��힘c�wEۏ�0Y�$Օ�ԙ�p+�u��F,��;��3"u[M�6F�������r�32��f{��S	ELW�b>iT׭��)'�-i�6+u�����c����V���U2���Z��@�LC�컩�'3�q�;u�Y���?Hrݐ�kr�Ew�.�2�r�|.[���A
4h�_W8���}�m�����K��Hf<���[TD�%����u��# I^�rD߷F5ʼ����Xܘ�5G{�b��Z	+�a_6WӍ�	ϫ�b+^a"�=q�K~��2v���0/��^�CM?��󔒚�0�_R�(?�MH����80�"��TG�;�髷V�r���i-di������@A/O�R����f��5ĵ�da�s���F�<����'�.�
�i�K���P����/|�֫aځ-�l��*c��r�.߆"O5T:�5%Ze�\�0���֘r�G���)����q0˨6X���-c<��m�:k�o:qrF�5�Q☨~��G�\��:�T��{�r�O�B��m��)�,/�T���IO�(����#R��`7���E��
�KU�EG(ߴr�u�3> ��罯���X�����u7��I�PZ��'�@[/��g�|ӑ��w��O���������9��W�4�D���]��!6G���l$���k����[��+�ʒԮoLMdz�����	T�4s��V���T YO������s&�ޡQ3��hħ��1���#%_
��핬����O$�G���Q�Vcc���@��O�/aK ^WGCu}�܅�k��6<-���kK�fY��bGe���I�WX�i��ǣ�*����2�7��(�d�>����|yXd�>�z���,c�ͮ�Y[M�;��9�x�
�����#�ɏ�0{�+/��J�g�;'DP}AU�r�Ù�@΃����Өo��*s��Z���7�g��ru<6g�i*n�eT�#��Cv	$i[{���-E7K�0F��UC�9�q�������S����+������_���G�I���ʁ�īv�gZ.�:m4S�ёo��w���O���Ǥ���k�����RZ�x����[K�����!%��A��ީ�&d�����7;`� �{�g8?h�>�́
=�Çbp�nw�d��bB�QO+�L�񫶚>�:�֤޻.!!c��&�X���9ʳ��h#���@�S4������b��FP�a��ԘzCs�W���٤]�j�4�@ f!n�n�s�O{��Y�cD�/"hû��RsG�|�O��^�,*=��&� ���S�Ec5�כ�?L�m��Z(�Y9��&.Z��k��(�jx�ʧ�H�ؑk<5�vXY�q5�@����3~6��OC�峞��^�P�~ouD�[���H���a�g�#8P2I�g2��^��X���dq�o�;�*K�5>�_n[����v��'��ȯc�G류�i2��R8�����H�]��KĤ��`Mk��!`�IN�Y.L�? �B��	lP����Ѐj��a���2�����X�8��uF�O��ƋSYn��I��J,�2��M����3Ui��ω�I,�h\��l���,ǖ����?�ֲv��;���͈-{K�4.�F(?+a����CΞ��Z�s�#8 )�#���5``���J�a��[�z3��D#�vH��`.�.�'���������B,�}Ҙ@T+���Ƴ�e�e��r����������q�Z��v���Ή�ٸ}�>�rS�4c�(Pf�Qb����uQ/O���]��� +����z��2_�5��}��}�B瓦TZ�c_�Y����~(-XѾ��Ii�B}�WAzbGb���y6��4t���(�g�$̠�r��C��+{*%6�&qk
\x���3/f� �'��N]�R�
bW��qd|U��˷M��HnX��x_|�Ź'�gEh��.�Ģ����ȹ��x#2~��EK/�]lK�᪙���Q�PG3h�M�l�J˾'e�K0).v�ҝi�a���@�ި�\���[�e�H����B��Ǘ�����*�6��q�j4p�ޱ�[b��8�։ �����r�waR��m��;�6���BD�[(<�+�����U�<Q�&GbX�˞^�ϊi��#?mr�E̟y�G�xm�M�����$�T�-Ї+���+�&�C��eo�;kzw���Hg�m�IwC�>��0�!��o�������JcaS��~�s�����1>?y�Ĳ�e��d���w2��m��\��M�3�G��w�V�����nL�rf��Y����KF}fx`�*:B���35��o>�N�o���'p�Ej��h��QU����9<<kSH@M��Έ�����F��%��S��UQj���;��EGݞW.�+�j�I���ݟe��������i}58X�z=��1Z���"7g�۞����-�Y�A#_���H���O*
g����߲K�a=� �Ed���B)FxKq�o������zQ��a8Cf6R��m�X3ɫ{0�hYY ���T�J���'_Y��*�Y�Ë ^�䑰R�{��r�!���h���"��I� �j�~�0���1�ީص�9�UOt�oB������%�+�L�-���v�(OE�e�(-/4��'�$��>�5�_��b-͐cJU������b�'k0�ȥ�����7���k�߁mw����F���͆�Ϳ��6��Hu��up.:�RѦ�C,����#����x���<�BNf;CP��q˃�IЧ��_��t�J~'�2��I͇Wk�Q��?���@-Y1q%�g�Պ�*�%��V�}r�x�R�RR�h��|rY=�e���T9�[���1$x�PЯ�obJ�g�&+\ha�ɼav��L�����o��Y�,����b������Г|aN¸���Id�Z���׊C��e�I�
��p�QM�4'�4Cܳ'���52�_Ve����&�K�d�"�,��v-.��i$h�Kg�P��^�Z�� �<-Vҏ@ �re��k���>ri>%Q��b�ψ��'�@j-�y6�a~9���>����[��6�˞B[EQ��e4�駈�
o�i4ۗ	 ǭ��Փ`�{������R8��'!o��d��f��a�;J|�d��d�r�*���ĈG�w��~�7r�|WcrnH1a?�0�ge�܆ī�`�P�oִ�ǟ=�����j�+Gp/�DN�l��]�{�������a�(�P%�M~ٵ2*�zocS�j�\6����v�$T���}&ЄF��u����AW�t��fJ)Ab���������t&���~q�e����Y�R�.+�������d�����wIK�Ӭ��ަS;�����SH�[���:k_j��<,�,�/�w�{�(I�f��w�guE�â�9,˝�^k,+=X�[}�7�ځ�	�UV*n������H���u��;��q�D˭�|Z��cF�ͭprUHg�N�]�z�����H p��,�8���X�
�L�9�ȉz�]������#t�?�[�6���u��w��p�8T��5��3�lJ������a�5Z��Y��N}���g��G! �
@u�]aB4Э�^*ߔdߍBp5g"�5�كOd�[#8x�wQ���&���i�~�#\��5�Y4��,����^\��ɔz&��n
�f�����ic�d��7j�1�L�\�Et����<F�W�c"�&0�Ъޑ����M �h��`�5A���gce����%|eғP��,R<�* �v��[��Y0��a�V��:�0tq ha���XY҃����y̖0ﻯR@���{=���7���Z����E��mG����ӎ�8O��~�� ��E��)�ئ}�}���	��M6*\���'�+xݘd�lR����_�	�����7�Bd�e��Q]W���=%g��O��L)�ie⦜��S�b?-�ր"i6�v��8��?��fJj5��f�m��T���#ܩ��+v�]���wD����T�<"��Y��xy����ӬjNr.ؼѭlFx#1}]�~?�"�^��B��8˘jQy����ph+��1Q�~ċ^��G�x����S��^7�4�(���]��1=n�����Fb��S��NAN�,z_qKB��o�0v�a���༘���&瘱X;S]�L�^J����� ?[]C���j��v�4��b���x��Tu�96�r�7�{tO�=�8���s��� �j�z)ʢ�����s����V�Osg"�NnQX��ۀ�:��P7.��i�Q`�)D��O)��T�H~(ް�=4փ΁Y!)\���\�t�u{U�$l����i�wڸ�����z䀮U8�);�8��A�R<3���'K��K����b��ƐN�|ڸ�h�n��ǝ5�ݼ��6��ʣ���I��y�9
8��ZW4G��.��1��C���67tc��g����@ׂ�r�׼����N+���� �4^���,fM�([d(Fr�l�5Q�Luȃ��ΣW)L�����ss˼�=����t��^�m�G�<N�G�>e�,<�;�ˤ�d�q��*��͗���쒬�ӶpL�)�|@���V��Q����z�g2!Cf�C$����rAsQ{�6��b���¶E	:�K,A ��ªM�[E,uVef�!����B�m���U�{�=N��)g"�䱮��r�א��8�v<~�T���Y�%bx�%YL����w<{���}�%��m@��|�U�]�-��� ��2�Qz?�?p�1�*�����x;�]oeſu������ș�X��U�o���9��}mM�j�������_u���cy�����OZl�
��@��W*r�Z���A���	5�M���I��<[ ���Ǣ8�ho+d��=�E�b[p��{������U�Ԑ�����f8"K�@O��n���L�㧼�okK�#� �JK�a��*]i���g��ssH��k��v���.g;Q�)�_��U|9�/��k�9����[�I�A��tiP��K�-�V���K�����;�|�Ī�UL �.p�RR�?~����p�<'|����/�R�G��$��`�0��Z�4�$��v�RȈY���kK��j�Q��)/��*�\(DH/)�Yմ��lL��ˍ0 2��RI�/��CL2~�s�v�L0��w�?t�Qhf⥙����;���4>d���)�E�53�~vQ��Q�&hF��ͪ�Nm���n�ܮi����P�(J�柪[ђ� ޳���� �,��z�M-�3�wb^�^^��wG�\��x�u�6h�aFCŞ&N��y�������DrF�^��B��֯�9��)�h��q��n�j�E3�*�{c�A��J��E���,�G(}�F����m��9ʺ�P�
WR ]���^v=��%�O	����Ti�����_��0Q8y=�rh�Ϝ#n�מ�f<&��\\S�����G�Z*����o���q�Q����j�#̮�U��U��غ��FVlA�ҏ^��M]��b���fbZ8�$>�	p;����c��>[���ml�9x�㞇�~{�}Џ��7���<�S����A�B�SF��!˷��h/2-��Y�o}�� �W�/"߻���6&����b��������	��-�ɢt�ڠ���������dU�l�E-�*8��
zSj)�F(P��'�$��:���RZ���;s�/T)�/�c|��FU�Xm�a�P��"��2�)Ƨ�P��Fpn�˿u���Hp��!��UE�;w����6�K�p\2�)�pPn;����^�Q� ��i�E�lW�Dg!��	%���?���nj����[)�"'��f�Cc�6_�p8U�(mA���>�Dׁ�7���8�|��D�����g�A����ݬvP�%�;6�B�W�1Ņ���5�T�*��*2۱�r15�j�GM!:���a4�5"�濻Nh�������;�}8y*޹]S����t<5-�/�?��^5�Hč�@^3���E���r��.�d�F'��,d�V"����mAg�0��f��z5'���t"�����I�7MP�u��at�J�C=Ս�,�4e���n��	�;O�$��oly�pF8k[�|���խ}nG�̰���C0�U	R��}$�uU:L[���AqB�#1<К�8�?�+"�84W�r(���C�������.V���n7�'�N�aH����]}���أ���oo��~Hn�m��~�m�q�z3pr��布I������;D����T'��~����i5�n�Ki��7%	5m� �V�����US�T�k@%yC�[w�Қ�?�F�L?:��"a���&(3H-[r��
g�������H~B���>��;���`��z>��/�$��A��ٸ�t�"�)��(țk��F�&����K%L��g��;4� 8���:��R���;���� �M����{G�����vp#i������%4���L=B�3�b��yVK�9��Ӝk�2Ԫ_�$�S�p��R>&A���I��zΣs2�zLՏͷ����p �I�:Fb�C�ґc2N�}����|Lx���.��I���K((��B�1+)CF��-��(W,��~S�%�bi�"�����\p<�ZdΠ�z+�hG�=���ע�q5�:6n�S
MX�/LL��$T8vR'�l�a�5��<Ӷ��;	�>�ɁJ^��(�1�Y����zCH�о�@���}L��c�����+�%�0
��J���zޘNK�bU������?�|Tfz���I9�ا?��Yw>����J1��DM��AÒȬ��2��۞}8T1���xIJ�x��p�]��i�����T���(�w��K�����[	�-#�Xvh��&w>�������?ר<{���Q�6n}�}p��l��0{5�=��	F0j ��1������f��2B��\�*���-�q7�.q@s��c��L�IZ&[�䛏�Ⱦ˻֩U�fvʳ ��J��4& [��N�q�8捬�?P�r.CM��$
9�&��G�fG�P�wf��jwR¶�
�� R�߹�Lh�E��N�gB��d�]m50j�R7��ʄ��Ր3d�g�>����z��*g%"��ʍ�VE
dwKz@�/f�*�f�ܰ��/�r�U/Z|��迗$�l��#�r; -��BH{E�s8P���Ū�(
3#��Ԉ����蘦B�p��h��Y���0H�H������c�<��L�6.��t�'���q���5$�LǼ�6|51�B�'�AO�j��f�q4���z�}H��>���d��~� �׭Y�m�KIܙ��cd6����,��+IaE���HD­� RF�[��\��
ze<2�D��ܗ>�?0!z\��4�QDt���Ite������f���  FO���-�vዜ-�KL��dET7XĤ�y+�EZ����]~�o���IfH�β�٭0�������W`���!^���D��j���O

2�B�2�r�y��6R_�1����ߥ Y�.�z׷����O� �Č�e��"�����k��4kj#�
�w��E�l���[�!0��ݷ�"�X�z��Ca!���ˌ[1w��8����kҬ��߼�e�^�fPy"�d������`�HՋ|?�G�+�9����a�n��0$t����c�H�|�U:ДYjLb�7�Y�\�U�������@]#��z-a-�I?X�j������p ҕ�V����J��`R���>n�]��Pk<@j!G� �i�"O"]Czɱ��v��!��e������"7~�������I���ـSm�+���1��쓗�o�/��+U�[���_k��2��t������w%"���w^�r�<��`	^l}SC�	q�
N��ɧBN��O�Ǳ�71�E���/@��೔-�_�7F\2+S1��v �#'��d|Va���f�cF�5c)�G���y�\��_�B7a��P���_6zl}Kl� 'u˗�"1���HKS7�#a> (c=�A��~@~	p|`3�u.�5��MM���~��&�/y�d�)\�X�]J_��(�����z��7�tĉsj�޵c�O�|:/q�d���	?��
��q,,�?����\�k����80������K<��� ��r9i�#ȫ@�᫧��ZP�[:A�wP��ʦ������8������<F��*��)�(˿��B��w��`���N�/=?<��� ~�tn������A�ҭ�ܒL��_��'!�����=��3���uܥ�.uo��D�L�:z������b�`��O�$�Kg����V�:��n�7��HĊn�q�Z�5�<�i�9�U� �CDT`N�k3Y�AlB��ա+�$K�8J8�5�̍W�:��Հ������Z����:K�$�d�e5�ZО�vpi�9p)��T���5����d$�2�K�׭P��h˦i��V#������d�Q�-[40t��8p-��m�/e-�7A��co"�LߣT[&M��zO�����@���D�y��/]���aS�P�[�'ϸd'!IC0�"W1��"�� `ݕ�G�x��X��%%i#���U��~7�-|��QJ�zVŤ(jQ>}43���䷭�~(�hc�����r�b�:��Ms���5�|�m50��h����F����X�v�X��Z��g��A��0Qg����c�><,_˽$	���Zg%�7ଢ଼9_쮵s��r�Z�4oArI�1غe/FSJ�a��.^ �^��9
b���N�($!O�kE�y"��:���]�g�E�r�����G�D�2������9���$�&k�L��w���4��9v%�����y�+&-�^����S� �4G��E�M���w2_�M�z�E�!!�QEU9v{ۻ��(�����T��]+�YE�x	ȣ%��$���pԃ X)�`����������d�ez��Om���f����cBW���!Q���6�VEb1S^�PuKH�
e.o�S���|4�c�E�r��TJ�I	��14V�^Nᑮ��$��J�?]��2�k!�ߨдd��΀�E��
rĐ��6ۘBX�?���,Itysew`���֦��w�"��ӱB��A&,����R~	A��>f��H��Kcf��q���+��&��R�q�����C�<�>��	m�Ѵ���'K�I��a�|��F�C�y���o�qm��6��tb��)Z���j����@T��w�9;���A����7)��4���A�g6��l�QX�V����e*lRj�]��`O�-�01dñ�"41YI��[�Ye@��1؞�S�i� ?��E�l��ov���\:wZAN�:����ߴJ��3�l�Q�=ks����B/�4���W����*aMC��t��C��Z�ڡv�}��p��J�t�R)���7"EKI�,�TBNS�p!D�{���댊AM���@�AՑ�	�6��;\=2Z"��<?��[�O�/B��ho�g������.�s��o��OD��e����?��"�Qޝ� ��0��4(�c$���$*�ű�T'�O
ǂKAw��\"S��ʑqEB�=���F�g@`�$!V�"&�K�SIwyr�=c�}X�k��c�4�uBy�RyVǒ�}��+"p>	�~�%\���	�d�zx��r�>x�z
��%�K��E3`�Q�4���W�$����9�9����HE���]��n��f`���`{$�u�K��f�a|i�'�e�s�̿)�	I��:����K��j<b�אʒ4�,��aݯ��=��Bh�=���<�R{�)OC���d�͎MZ7��
ϾR��r���5�mM���nJ�!p�쐴kE���7��#�jf�x��x	���h������l/��i	:�(�ۻ��<}z�T�\�
O��J&4�񪰋��B����/AW�z.S�W�ä�ayͣd�"�>լ9Yx���CI<�M��c4�VQH�����s�L!��X$'G��^��$R*�rU�H9d6ͬxmjR/�h�h$P�_��Dx�{���cLs�Yɍ!$y�Y��a�`h|�2�Ϯ✒/-8�-xg7ʭF
Ə�_;�0-I����ƄF7�6�w�4��Q��t��!�S�Y>ædz�y]�;�����\����哢�¤X������T�H#�&>����G���g��S	�fsc8�r��G�=�h��bd��7���Js�n���}�	-���-�h�?qvmoy쿙,s�[��Gc���0ő��4p��%+r] \��Ó��_��.4��4s�}���/e��W�_���=�1�����Q/��<���_�'D��?HR����z�b�:Ri͘��:�rW	�it����0l	���ن�$h���Uh�)W��N���#[*ҽg�s�c���KF4@}�ɷ��YH��2u����+���	��bUH��e47f�,�
���m��mYx��&%�t{˙3d��-D%uI%�KaҴ��3���������e[U���xT8�Q�	iB�|����՚��B��<��T1�Ƅ�r�'��rզ:�)�y2.�'��+�{��O]o06:��d�L�PF�`�5gvy�e:�%��ʋ�����`jݓ��%���圠`K_G�4&��� O9{���ɏ%=�4�E��m��}�:���tƉ���̼�4�$���c�-�gk9�p�.��pZ|��P�Ī�o��Mݭqjy��߶�=]��
�}%���M8�&ߊ��D�5�Ψ��U���qd�y�7��oI
���-��vf#}�3��&ٺ���o��|����y��ɨ���5j�<S�ҥ8��'fĻn�5@N�;�	&aM�I�J��ޒ�>�a��/��'����:�n�ILb�
���)�ڴ�5<��	��XM�Bˁ�GH�gT�ڧ�9�4�Md�|�zq�/���F��&��}����oj���e��$9:7�[D���Ei�q|�6%c	;��K+��5�c��Q��N�d���[@���H���`��������Nᘥ�@d�Si߿Ͷ��@����94�I I�H�g��=�ha;��e�����h��b��2z�
�+��93�b,	�qS��F��V���m�s� ���^q�٣^��8��c3���Ф�F��u��`tD���j����r�D�z��m��ͺ�h��m̠���I_��f�oS�^&��R���NeR�w����l+�I�@�C��g�	4�Ɲ�^Ǧ�0�Rt�� �T�s_�QP���Sw_V�"�����3�w�������?�D��p�ǈ����?��~yC �mu9����]'��!��.i�^q-�Ӎ:c9El#�7k%�T�m:�@@����==g y�A��C�=�N (�HIZ�ob8�B�b�O /`���9���/5�,����_ y�[��<p ���|������;��`�/D�܁������r8�Ya	��X���A�����f��m�s<�Z-�Jʑ/ͧ�l=�ZY �>�߉%k����U	�U#'����$���n���jr�4@�:�X8aF`�պ�k�ծh:��3y�ȸhE�E!��4\!Q��ܯXu��,���������U ��<�D�9�T_ n̓����d|��S�����o�]��,��|�p�ĝ��x2 ����y%Ԍ�i�����ќy�,�xW~X��*�(>aݘ�ێ�Q�-,�.>f�hDj��m�͌1XyLPss�!t�B�&i�,V�V�bƢ�ȴ�{�B w���� �-0��N��WBo�l�׵`8�t��0��~w>D9�|�Q� �i ��S�;��dW ~�K��B��|T�4@��d!�\�A8�B�T1[�
Y*Q�rr3��/a�J��H�[&�$gCiW*%	�����J��]���}��H����%���a��J�������ٰ@�_�Xq{�(a\�$2=��5��;�J�Gn��xI4�L��L
B���s�V0Q~���a�=�{����QȚߘ��[	��%{�n�W5�e(;+��k�d)��̻�	&����*?x:��-����=[�w���}�>����d{pUP&����e���.����ײD�O@@g�P��q��!�L�SW��TzC��G6'�G�X-0ͦ��H���[�ݺ��6��?��F��l��9�$���nR���s�,����D���=mҖ����OGa��Ҝ�%Ԅ4�6�sEG�80r@�؋!�e��������5��yEץ���q�c�8�-Hד96�f�?_�+�Y-6� FǢ��V��M�.���۵O>���\�u����{%"|>�'�d�m����@Oʍ0z�#���`�79�'J����:��H%?�:#�[q�y&�y�"��֜뻕<K�Ę���8J���+I��U�!�J� ��ܩW�	�$��p�J"Ln������BV<n&��P�D?�x-|��i��[v��GY����b�cn
�K^���V���ڸ,񦄑5��v�I����d�{-�̀)�@�{�����!�[H9� �ʤ���`��e"f�Hoܐ1��1)����w����
g����^�o}���}�;�I�������96��¿�tr$E�\�j�N�� [�2c�+�8�N�0�R��
�:=c#�T���j��Vw�i�ͥG1޳����>*�d���"<�l���6�.����bͣ�>��H�w�D��fXxE�é#����&7��s<_���s��]���ۻc�  =Ä@7��N���_�����]���T�`^V�=A�8=1��҃HB&��Q �Qi�{e�9{�	���t��?"��K�������N�v6�^��t�1Q�ԛsh�=�F+�D�9�U�+˴�A�33�I��_�T���z��i\�ѭ!I}i��ln0L�^p�y�B�(��}Q�t���)!y��lJ��܋s]�!�}��HC� &����M�/��
��I�a�4�����z��z-q�����a�Vp:6r��6���0U7�3�+��렽v��;�.���d|ו&d]�պ�/tvmw��Ċ�%̢;��&��L.ZSX}���q�Q�EW9O*:�0[|��,Vp�La<����6�%���-���@�����0>�\�>��ɘ�9#�oM"���ۨEߝ�Rk��J���r����T3옇	h�]:�3L�� tRS>�8]!��%>�<k�d���ӸP�KJ�B���!�Ow�����嶛5�i���p��/�9���3k�m9����¶":��}ڦ�q�>N7(������J9���� ��r5�n��JyhiW���"�$��E|��6x(���?+"��qGt����0I�$���b������I�6���B�Cf��X�+�p��A	J����*ÕM���B�>����V����O1��c�<�Ҿ8>�>}�4k6[eZh�"	�ZZ�Xj���>�^k�Gj�������Au�O����}2zvC��"�����y^lg~6�8,���	+."�S��]�I���[�M��<-�vV�޺>�>l�ݽZ�z���My���x��ܰ��U��k��>��<i
�oo�+
�p��ȓ,D^D,C��8+{�f0���`K?����5Lѷ'_�Ӡ�PU7#B��-	��6`1#�K�/֎�Y��ȢA�=|�Ym'�B�G�е˭~U�]��e�%���v>��}� 0d��P�hrZ�
��sq��ۘw���l��[�ãd<��fCr�ٌ��{M|l��Ai��Z�V�
B5m�б�
�܄s�:�9o�?�b��{)
!sl_�H����P�, 0`�� jF���V�A�u�ԫ��O��|����=�x�2vT�a�%�1��y���#��"�k�Zw:�g��r��J?�t��q��0yG�W�ǯUs�._�>���q�N��M5�X�A��%W��3�Ū'_~��P��71l����'��3J�&�6)��V��t�R�>��-��Z�����Ľ�4oJ�L���i���j%&OQ6!�Q�K����R
)pS�jػ��ϻA�̓׷ 8T�<n������q_x�lG�*]Qч���K}	���@[A�ߟ[;�;Ӹ�'��!�w�0�rz���YB]-�T̆����xn
8��y_5w�ѿ.�e�����fBI�������� �6�����ۭ��~fd��K�h>�p��
��G-��Э�qvίCj�DY���Z���R]c8j�#'�`*9�kD������[���~:�@G��
��}\g���1�Qq�y�E�B����b��KDS�?!�~�'?��O��G<lw0���C�O��\t_-�OSH��#�I�����0�J�����q��b� ½n�'z��� �Ny?�5j���b�1�?Q���v"��5N���Y������NwA��o�������d�&F�h#1!���=��I����^�"�V�����0=��PE���պl�Id��C�9��-l{Ӵ�����̠<�FO�Z%�WJ,��8���Y�
�Ⅱ<�e���&K��2IU��Π�V����3s9��M�=��YMY�iOV�t#�}�r騟l��eEj���gW5����QU�wЁn�D�������Y�I�w�^w������w����x���$\U���b��|!�	��j��sN>H^\?]�C��������&��7�o�s���ƌ��U�>)�#���D��}�s�:����E�4ھ��/ݞ�,*�00�I��x��Q�����P�� �H��W�LsխO`:_�h/�O�	��G�)�S�-�U5~�L^
��>6;�(���Ym�F�[�{�N��ȭA_�s��;�w�/�g~P���X��֚nMy�H���mBlWV���M'G�d�Jw5��؝��IoZ!GT����Ff���G�����Ɣa&�=U�z�U~	�f4�=�<�sTN���*�~��N~����H�����h����z)��>�{I)N'�����b��<3�.|���Nf���KYj�\u"	M&?��M���I�{������t3����My;j3�h�u�n����%B�d����}L��D7R@pŦT�x�$������,���8;�:���A/CZ"D�d�+�e�B%��v̘�ߩ�|D��>_$��Ð�5�MdvD���D>�N�)������7�=�d���A�;:mq�w tM�ߠ@���j��q��\l�Է���W	咭�'����m�_:n�~����)���\/c�E�`��C.�n&�3�"0sP+�����F�e��!8yu�K��{.(���d(V��,@��"�I��K΂jüB���6���U[�.�� w>9�q_�O����b��蝳�}i����:�H�7Z7{T�G���q�X<�����T���Jh��_��DZ�r���F�B��<��P�Y?b�e��9`��yh�&t�{ے�U�M�� q���)�u�(���ÆD��n�(Ѿ%歹�w�H��A��#y��G��TJI�����3wD���t�O�ĵ!�Z�ʿo������	.1ᬣ�����t���4��XR�W�}���}�{�c�MD�3�p�n���
�� ��}y}/7�룬[J���Id�]���+�b��~�Im�1�a���UHdL�_T��G*����L���- 'V�Ic���{�D�K/�]��ב}ن��fԥhKL�Z��>��NZl���E�90(�c�M�J���I��)�ejVj�?'!ZL������ �dl�H��>���}�F8�:ŔH������ɳ�zp&c1�Y�o�Ssf3�I}�Z�0!u���L��n،��GǺ�9p"�3W(�y�X�^���m�h2#�.A���rn}�e��	���y�H����L�d|�\u�\;2l66�H�J�5��?�kJWt]�XGoX�p���2��q<�p�Ҙ1�b?��X3L�j�EZJz�'\��s�>��@�o2��_.J�+����x/v�k�w���g[A��t�S'�q9���x�@қ���u����+e�=��Pi�oX���"�;	q=���P+'|�oh�6�"P�FP�v"�^&���ri�^�d��y�CD~�t����8��v��\��!�"��Q����ר�U�"��<�X��w`ٓ��O���%e��ͦV�O>ܿ�F}W����*h#�I�� v��dL������ѳ2���Y�i7���q!��A��-乄�חQ�ջG�Ž����t���݈
ګ]�(T�E!���s���]� ��߂cM��	����׍���Z�)� �O6=�NV�7p:��i����TC�<`���V$H�	�25V����Ș�{xw�|��@�6���ϴ���a,a67� ��
��߹;x�e����M��<�����v2�6��I���I�;�t�b�
�F(�,)X��
R���|q8��"	���"���I-q�j7��WS������9�����б"����z�圐�s�؛q5�6&�� &6�oXQ\ճ���E[D��xA`>:��gX��q��`\]�B�
�b���mϕ��x |>�z-���$�t�_���o꾢ģ�,��
o�n�T�0>��I�(�C��o.�8�-ɂ�8�݋_���l�Z�I�1����BRvLȕId+��9Z�a냻��{d^�l��S��̕|Hp3���f���R�p~/{�@*v�r-��@���!$X���"	H��o�j?z:"3N�{Sm[�kS������s�c�^c��|_+C9Ns��i��{�f���?�9S��g!����&�n�����Q�5O!�r{2��fn��� ���E��
*bg.�f�vk��u!�>Qkn��XG��Q4�C���l��0a@���S�S�`�W GT���}/�򚉹W��g��`�:4U�#����iw�:�� �h��AӬ�R ( �ț5)�D"u��I̤ny����`��d�|��0��?OH���c\�����<�k����� ���ڡ?tRӤ�AHʔ�%����;#Vc���FmĀF��wh>KV���H��U�gÊ�VlT6(5ˬ�!��)��ښ&��d�1�6��o3<���Խ���M�v.�g�&h_.�5��u�Mc�(� ��-*�B�\�Xz�j�~	�����qь�{.���-o�K58@�[`j�A;���%�Ud��b1
W�jt�0�Hv��c�l�1��Gf��A@��k�-�2��N�~�|��2w�|��pyfPRW+�*N| �J��#���v�k�u�ϟ��R���fk��,�#�NRECϜ�hn��:W	��Υ���f@�/��`
]��>��I{�&%�K��|����ĩ:*LYu�O�UIZ�L�喫��HJF�~��Z�z�� ����n9	���0�ӃF ��]YK�.�g��p{�ʬ�0I���qū�m�������|�-%q2��:[�tΉ�hQߚ�@7��,b��FA�<V���8��6����6���F��x۞����f�X2�n}O�a�Y$�xF�݄W��ҩ��ZR��Ve}�̾n�>���[!,m;Ԥ.N�<�$PD�N-��Uz�b���DO�(�D�%��|������J���J�v��V^�d�w��]�/�Ra��G�]�1�
LIHQ�aרn�HZx+`T�|P�T
H<�њ����, 5�z����>�v1%l����|��������>����
DE�7r�n�cG���;��=+�20�ŗ�����E?=j_N�uvvˎ�F���.�t���?�9baFu� xm�!���8.y�_.tr�W7c�7*V����Z�H���a�J�Լ� 	��ϕг7wG�#]oP �`���#3��b�܀,����YN��ҍ�Ew���ԇ�uv���}<�&�.߻Z*��}��CJ��2�P6F��(�G�̂��S1#5�2��t��Yc��\&� �e�r�d@ο��!3��Y+�XǓP�#L>�Z�U^�Xq���� l���3��.���������2�<���[��Uj�p��8��$��X�QF&)��`�8E(f�r%T���R8�(-튫O�	H�A��P0�D�vm3o����}K���|Nݫ�w��b��yЫi���lM���_�~��L�7�ӏ�S�zD�/�i��;�e����Hĕv���j<0[�|���-kh��X��c�WD䙽�~\�p�͓��v/q]�x2��Z�����sA�G�L��x�6���h:Ί{����K�A��-��d��N!873��+uɂ��!�w��S@��s�ic��h~���PR��q?����� Z#5%Pa�l�ZƗ��t�������U�� �T���f��p'�(���V�Q�ݕC�Ϊ��ΐ��r4�	γ��U�H��t��;ф7;a�|�2sE���'()_��/���3���j-�4�|���M,]���MG��踲�
^3������>�>�5
��I��3�Ӕ?�[���ڱh�8���mc"��`��!KL�B#4u'i����9'A.es�kn:hAts�Jr�ˍ-���kf�/�P���n��ۖ�&\dL�ݥ��Z���!s5��<{6�&q?�d��&YTE��~��l1ߡ�~h
x��LM��i]}���h��M�.-V�|�.���a��8v+33��}V����a,���\�[�j��$�U�@i5_=����6T4�X_@������@ Y�?�|ј-����`2�e���4g$�1-�K:���&�����˧*��"Qߋ�0���j�����c�����;�4H�}�~�n$�t۪�)J���F�X�݄:w>Vz[�R�5�=UPs|��s�I��(�!�$��$8H�����.$$Pe�����~�l���t�%���E�BE�3NG����9)^q+��C8��h�vR�٫^Lyz@�Bo��P����ċ^H�N�����Z�-4�7��|�����D@%�����t���&'�i7��ky?���xi�p*bu��e�%4����@���nEZ�o{�=US|E裱+�b���3��B�Be�jK��4�Q'�_� �P5j��!�>�rt����"<����h���o�Y�D�c��t-��JZ1�$?��˶���ٟ�����>��-�h���z)HG�j#T��<��� �]=���/ �	��W���$&n!Tj�<���U��s���Z�Cʝ��Kqh.N���{�Dըڻ+��]*�޴�5�RKW�pRWhW��=$<�I�܌W�Z�/'t#<�$|���M���3���O �ސ�fަ��i0O5����������?G���@����B��p�T�xK7����h�(���%��oP.-[��rKptcրs8���È��x�n
]n�׃�u�t�cײ�����}�v`��B��[" ��fHh�.xET�&�VaV�3Zݗ�6�M@�R���Zȇ�v�r�å�6��؞�9��1$��Y��JkU��\>?�U�N�u���\�P���t�.�ʁ�+.r���e&/��)GP�Z�Z���)t�ĄeP7����<2��ѷ����q*�{/Ίų��-|%�*���dL��2n�p�Wْ�~�T.s��L!�z_�k �@�*�������pq:��5�sgh[�~���Y��F�q�mD���y⸎_���+C�3��[�8��)5��`��
,�����`��\P�cs^0*�@
�z��m��E+��"Wgl$s´~Q���ؚ|�����<T��n���j��UV�'�����р������8��1��O6���*�2m������^+�Uu���Wyw��z�:�~o�oz��e���O���<�n#�=�L �j~.׾J�"ߤ)[
���I#��-��!��aD	g���kS�t���+zT���z���r~enu�}}*��W��oF�3�՛�KsVΊ���y��ߊ��)�PbW�} ��%�*�^���G�n�.�2���o�Y��� �z��P�����g��j8_�۰+���k�6��s�+p�O�>U��>}%����5�)8��Ĕ�f���F,�|7�pĢ�46b�z|6�yh�����7e�W�{�����z/�c���ar3�V91�;��j��)��hS�r��0�'0���he8�-5ކm՟�f����*Fj�"�u)<���4_�aʸOm�u��� ;͒�A�F�x���"��&$����<9��(�j�IR���B�&IS�a���^M���:����iǣe	hO���֧n����-� �D���C�D~�%uR7���˚���L��~<�Y�v0�/=��>F�X��E���H�H>���P�z��:�Q���:���_�c�B� �z��℻�#�h��+^��1�S
t�z��2"*�!*=��:T��˄�`��]2��R��.�5�d�`La@
��[j��0��0�9������t�UލI���#r=
!���R����Jǩ�HLǿq���������Tm�9���u���o����C��ڶ�E炢5ME�)�����lbg~ôq%P+�jL��B�]9�0^�$|P�1P�c��G��gA^/��o�:Q�q���Z���4��P�uzEyt���0-|yA��x��@icF��C�]���G����������M@<G0�|U�X�ٶ)$դ�����g�>����݉o��AE��Tf���]a���/��Ӡ�f����U���!��W�2�}w��(��Va12���A�c�������V�j���i+��rd�X6Dg��Im	��f}y��U_l���X��l.�0[Uy���mA��Y'F��K�P� 9T�H��D��㾤��A�X��2��(�9�h	�E^Fk�K����E1��8ZX/*�/�	��Z�� ��b@&+X��ݏ��q߿��#__0g���\pP�0��7'��g#(���ip�P@LؚPI�������d!��� !�2C ���8br>qt�
�m�UA����	9��r,*W|��-=h��*���`S��0y����}d�y�C�.RJ��Нĝ�-�"��5b�#\�Ih����^�XDp�NYEN���0Zѩ&��ˬZfe"%�B��2���9�t�|B�*(�e^O�D�Ux�<g���4��)'f��;�g���8��I`���!L�qC"u��WV1���i�R.h�|ژ.(��HN7 ~�B�a��dA�fpH��_��a�Q�?s��&��@�A$�m�v9�ؠ>}=�@<a�v�~щ�0�Y�E~���� �&�&�'&�V��vU��DRF#hI�k���%ErM>���OinQ1�����Y��J�J��P�f�K��!�V�B�e5�-�ɧw��G[�vE��V�_���汞����BTi֝{>E(N�������]w�~B��iK�x�ƦyK�}D��
�Ay(.=�]�$+Qd�q�a9ěA��%���_���	�'Y @M�r�D;���DDB�G�{҅ZӒy	��9��>��?$��pz�/�U��N�XQ�Tn���j�=��5���?q>Pt/�6jH���� �2�Y�H�s�Y7��u��WC�%�[�C�/P��d�3��>C&����!��&�3܈���-�Ù�1P��v���z I�5�Q�`�Ჲ��Y�"�Wі�FRP�Į�sF�dd�'|J��t�c7! n�bׄ��V���F�.{\<�:��#m��,���~��{عS[F�ֵ�M��Rk">��ީ&�-/7�"`��ܸ.���Y$Fŀ��m��б������ �8���)�Y����ܹ�2��wh�[O�`~�,�{�W�!�������.�	GBE���@��*q�\��Dꛎ�d�p(|��cr\y���.�L�>@�.p�3�KR�*�Y���Z~���qK�@�dt�;C�zMأ`��c�y�/oֹ�6�M�\2E���"��F���o��lVWc,����b/tPh��Ç�J�h��.;�^^���/���5�e�)��٤��+�Ƨ+�'�e���ҏ�& Y�-,��]bf3����� �D��$�ꅱ^p������8�B�4���/���p�fZ�h�j�"o4o�̄L*�P�� �0n��d�wu�#Y��l͊�N(s��J������u��iJ6�?I$8qTG�`��#��2Pw��2u"�	��j�>�o���5ן�Sش��Y��\G&=y���s��[���v i	"�\uOND�3���D�p�qW����g���u�;|#�s�9��2��
�b[9=���Jq�[�]ГY�t$(ײ>c�^sq_v���:\3��V:����o�n2���s̐�5�S"x�0�6d	�:?>����G/��X��5�`���GE���*��/L��{�J�4���Y�z2|S6X�ш���Um�H���4=/��QF���"�FwnUUŠ�����Р�ʵAe�P��;���u-��#���_9�#� �m�9+� ��g���x�r���x+�тR�CF��=(�ϫ`d}W�xp���2I:�^Mq�D���)�K��(]Q��E���`�eb��A7��8��~�	�5K���^=�8��l��ZL� ��!���t�C}��X;8f�%,Y�����!z1!�UKN���J�?�$�f����8)8FN�^�t�ׁ̰Q���	\�ʮ=��5}4��֠�Gd�����s;�k�@M]/L/��$�����+��$����q�$ �j��O7
��6	�o2��݌�1��������Db�`�%��q���g��F��.��C��H\��ϔ��j�K�8��:�5F��`S�G�8���:)W�u�&H<k�K�ʄ4���q��0�D�(G�<	�l��
=�m�����3���M��4W'H�Y���e �6���k���뀒W$q�*u7́�#��:���O�Y�-q��R�$��ml}��]ZQqsD���d�z>��{�
�ݹ�����!����Y��#�+BO��Ua�ɨ�Ej�;����1ݳ��p=B�-@��R��tz�,��}F�/-��zHxa�1�Q��:<NƋ)�N���)x	RD�
(h�̄aF6�f۴�R ܫ�R㡫>z�NO�+;��I]���� 0T������VT`C�Ub�,V���7!9X)N�+����_���EZ�xn^5>6���xr����$���Z�]8�s�a����$)���̥ؤ�r��4�Y��.�dn�DT�_'d>�"��n�Vb����%���%mL��\%m��t3@}�rP��7&����H)��okx�cM��(L�M����˒�-~2�x�Ћ(��U}���`x�Ԕ�Z�^�C����G~\�v��`�?��E���[�$�m�vo��U9O�E���{�m�����2֩�NN����O���&��~�NB�"�_;�NX�<�W5@Ȉ�����]�%LT�y��=�T���Y���Ӑ���� �1�B,k]���Hx�E�+�Z���6�_d�(K��l�0��7��kNV*����}�W2�p�N�c�)�c�(��H��oBdW6�����Y#	N�?�G��`���\e��j�(���I��g����{�F8�k�^���O� *�+JܞK���]_�b�T��:9Qn��GH1|��p�}�z�90prH8΅�W*h���0�]��Ow��]�뭢��r@���G�S�E�`���ubbc�UX�h�_��r���r�V��*V�s	��������;O���%`�� D����ĠوE��bZ�`	7�����HD�N$c���
��2㜥����[yZ�sM��L\x��* �0oeuZ���k���T�������l9>��8���t�a�%��x+	��϶�_���<��8Qy��#�c��q[t��\M6�/똨����G:t0\2ZT2���,�г\i�
�3�-�����F�]C����!{��(�֬6gU�k����z�줨v!�,��T�G{l����*�=������%���7�2w�j��<��#k�!@�/;�e[>��RnLx�8��	�zFD�!���W9s�C���É(�:�bK��n�xu�~"rd&����_l�o�!D�G8�V��Δ3��L�6���t�A�u�����o-@�.�᭦�.������vj������rQ��uǾ�6s�����W%0����b����a�n� ʚ"�}L�&tH(��v���7]�b��76��ǚ���@?+;I׭��w�������jGr���R���g�x�����ٙ�2b e�O!x�kS ������ʬ��<A�h��2��Y�>[4�a{L���5!cP{`h����[՚�#%���u��Ak�k|K�2%4�H�:��d�VH�1D|��l wp`��_���//�Ŝ���`PE�E�PmA̞x�ȡ�`Gփ�Q�]ؽ�ψ[�;'��Ci~�7Q�h�r7[rg�+9M�x�EC_�_7��/�v_rԯ���8��7E�=4��Q �|A**8~��@�l|����U�7 ��A�S�n�v����:":8�k�e\0��-~`�I��F[ݯ���L�k#4m�ψ$��.����wa�ή��Z�(DU�O[�&�	mNh�Տ�ĝ�=/�EJ�"�c�4f�JOy�!:��2}lJ�4Po��)�V�v<�F�C�"�E��,���̛�C������B��O�&L�ЪI{���"(Mwu�)���WJ�;�ȧ�f���rѡI��$����i����4�W}�-�'���N5[�� ��?yc�̺_ۙB2�f����nl�M�6m�Z	�9��B��,��y�6��pgKz��c/�h%ԘD��ٷ/�"����Pxs1@|d&��HvuA�%�����s�j�����fj7v��t8=�}k�&���h�����Ǩl&��a>� C�FtaVx�:�	�{�^q�,�u���B�Ⱦޭr&i���CW�sw�&G_c����Rpl�"�,a���'��=���:3��e׬�1W��#�X�g��$��k����9���X�#�J��j�<��m�Q�#��fl��\��ۻ>�����(_cYg2����}+�%%������?{�:�U����3�/ qr���Fb��x`�S�wFQM-�5%o6�z��b�h��/Թ{���?�+9�P*7�%�؟����S!��e�W���x�i��V�DW���@�+�ܲ��8�l���a�P	N���,"�y"���͞U�T�c�~�G�C8Ge]�)�J]�w2�K	G:��se����"s�_��T	#,'z��ė@bw$0WS*�>_�(�]�6�[�����@�͙��0G��bH���R3�ӹN��}��p�E�1 �]kI��i	w82Ъ8:)�/v�=����{V�/b����*b�Ę<�J?eLl�p���`��L[�G+ �l��:�M"_%q����
wYNߌd(��;�y���쳹�E�x��Qo���T
R�]��U*\u�D�]Lq�9�6��H(����M��n�Ԡ�h��n��`@�mT Xc�. �(Z��a36�_si���`�F�e5�:h��[g��G�H��E�$��1�4/S�P���32� �)f�К#F��1����$B�;j���w���	����o��\hW��9)Y���}�G�H���㡑�!l����逳w��]1����'��� ��O���`Qj��|�yS� kɤ�P��礜'?���e�g_"6G���x��,�m�MH����IX�((
'��2�����s��O|'Q�x�k��x;h&�)�?��.jyPm�j�{xuO�:X:[��S����!	U�ѳa�~�>�¶+uxh:R��,��� YEK�����zd\�"+w�Fۆ�I�>�m\�-�� @�nm�d�3�H�����w�$g�}V8�}�Vc�3�p�_$�!̺
��U ��5�����r��}�,�vH)׍ ��{�L�.��*��l���?�%E�2�j����K�sq ������}�˩['�L��u�J�u��70e|��@h�%�*ʱld����H��6��]�F)�giu���e��@�q���"i�.�~55_�z�e����B��J�=�S��rw�_���!��?S����&�i�@��e���H�<�J���{����I�m$����xlo}ح
ǲ�w��k?SMbІ�w�c�T��t��� �W�`�]�7&̑<e�=��C�������ql@f\K	|�0��l�]*ႁ��J�x���`���1��8�l�e@|b��݋>��5�ڔ��-rG{}���b���+L���ĐS�*�~�Z����I��.��z槯���i(�w�	{��f��&������@#�8�����腢��9n��?Z{X�C�p�$(Q���X3�xZ�Sht�x������IO5�y]��'ā�qǞ�M��i}ڇ
1���䂕�p���fI�ς-������5��~�~�y<v�J	|#�6��);�=	�w����c�[]c���d����y3������@�=k����G�q���<��I%�����{��/��/q!Q5�rT�a��?{&��խ��nŶ��i���c�@�=�V1|�w��px�`��&-�5_�k���v��1�q�����\�1���72i��4~����-c�?����
��t��Aؗ�����VR�$��?�)���N��A�)$��f^Ko]��VL�۳�P���[���ቬ'�~ǪZs颤�ڿ�4%G�^����
�ktRs�x����N� T�MRc�D�|>�&�'7z���ԅ��o����-�8/*7%��y��}���$���8�=����P4 �ING�ܥ<Y�uE���R�;z$�%��aB[Yq_��L��+�p���'���Ͷܼ��<���&ɕ�Dkb{EV����g�^�5(�d�<٥"�c����[@��8O˰l�%�G����:Ou�k�x~�ܳf�,�g����_�q�R��]�ϥC�Y��e�64��̭�Y�+O��7eb�Bu��d����C�*�}����Zq���v��@�6�F�0��[�4��K�;j��TC���RFV�V_��n�ge�R��i���S/uXna�V:z(a2�䘤����p�<} 6z@�����e[�fGsNj�|V�ԭGtd��p~o9�@��]�:�{�2k�]3�ڹ/RS��~f4[ɴ��o�,���u�z����2j4�ac\0�!��Zh��]o��y�}C>4���P<�9l�e�\�85w7h3G���$G+��\-4<rLGo��5Q���Q�R�y?����������E�71r8<VIH�n�H�k�Oi��iẂ�X�j���ͤ`błF63�OB��J�:��c32���G�2P���.#Lr�k,g�U�z���U*|�,����.��2��\���L�f�nǉ]�$�&zE��F��� �i�n��n�U!}����L �Ц�O��ˉ&���k�,��O@���S��zDi[jzq�p�0�H;a=�m�wf�<+���3���劯���F	�����Z�
�ҴE2,�Pq&	��4�Bޫ�>����+]�G��Y�$�N.�1�P���f���ky߇��nC�@Gln�ҒGj/�"Q
�li�J�m`
� �u�T<��y�/a�V��9Bˢ%l��v���x���\	ѻ�נ^/�ɕ�ƴW������[�|�w%���|�t�x���Ö�(ܺȹ�f���!V�Oj0�7U��7:��gy�A��Z�$ޗ��P�A� |������ꄕ�����b��� ,��#U��F�=�%3���-���Z�Ǫ7t1��ySz�gV-���}�P:ފ/�=���Z�$XPߩh~1r�,c�SD b��� o��Y�d/君�lR�C�2�h��g���l[U��;�ͤ��nc5V�o�]{h1w_K��<NB[D��~����Ms��vo/��x ���:9yn��%�t�'f�|`�K���4U����a?�<&�{�ʁ�[��Q�C� O~������O�i�iL���	f���>�!�|�Wat�
�y,B�@h�v�����)��~��g�W�A�݈�q���q�s��`T��n��I�����D[�r����V+M�a�:��-C���v��(߈�[K��k�@?pϽ�+�Tƞ��\_G#��Ob��Pߩk���8U<���p�l,��g�����S̆��.`ڞ�q�fU]�Z�"X��8ek3���0z�ט�X�L���O�!��L�1m��v�~P^�}��2)����TC@��5�B���@Z�Y�Y2����Ͳ%���;_&�E�/!��9O�-�+�!�@�X����r
���j_PpV��+̭j}��D[���¥�W���dP���r'��]�L�~�F� _@IY�U���Q�f�9ªh����%g ��M�\�X�-�Pj���u�F�ڰ�@��]��.-�[�����8�<98Fa~���>�>��j��}�PW����� 	����cU;�$6Y�&?�䗓�U#������[�eȀ��_Jf$����5k8t�;=��H�����l�$7�c�&�O�,���#P4Hx)�\)q��8r�8�U�Yk�,n��O���%������ݻD���bG��]�����^��tp�fe�ͣ&����������N΢�'w�8��9�K4f��},�Y!P�^��v����Q!ߠ&�sM�+�RSx���拲�	;_M��D՝Ln�/�YB:$0���bD�U�Gk\Usm0�-]���3ig�9�w��(�4F�~|�,���0�0&0���V���,OUS��=����J��f�P.���"��gH����RF+��o�a���Z����\Ǉ�P�g'�.
���Y�E���һ]�s�O����Lt3zY/3t	0�.����i�q��a嬼^$�3 Ւ�
z�P6������Y�����{�̊G�-�q���OQ�8
Cȃ��n@3���J��?9QlP�q���|.�z#�%y����n��ጢ�y�~oc}p����|�鋝�\�<N�톫����U�-@���
ی�:�7�>T��-��į��.��W�AcU��uK0��X��#�?� 帓j�����f%s5r�ZS�^u�{`̹o�_w-�u�F�'�N����=�ʳ('mh��!�FL�����'�b��~�1�j�ZN�v���Pk�o��ϔ�"_	�5��"} qWw���#F��@���\o"B*_<�ϱ 3CƛK�Ф�n��i�}�$��5aS�!n�}��S+���~_�����Aς�1N�d�V�j�`��ct� ����n�,�˧��	��%������P;�S
����֚),�R@|0fe��RIݏ�.�5�E5w���q���Œ���*����ڊ�~S��1�&+W�x���k	���\��?����e��q���1��'���N�r�|��LÔ�滀b��I,w�0��V*��i`I���Ql��_s�"�f��_�q�Z2v�Og���C��ǅ� ���#�Jka���?ﾾb|u{㠿�1��H�jǗ
E�
��=k��i��p�A8�cڏ͍Pl@#6|�߼f)XYn�(�w���c%A�P׫�����s��]�8�#��U����|��#Q��E���r�-E��ֲu�*�o��D1�Ӄ� '���=˷���;�ŋၐ��_������p҈xn�s�}�ܩ���������^�0	����E�ǘF��
b�Оx�ME��	&g�wuYa+�$N����(,��`��;p���٭�����5�pe��*���z���A�(�>�)��kij��*��I�d�&&����G��5�e�6��8��H�Lcȋ7�����>�Cj�S�'{�Xw
e�>���&���#���%Ӆ1�x�q���0S���9���K�P�o��{����.J�8�J^n�%��V�1r�Hӝ�Ca�x��OP���A��,!��uV:*���P�������_�"	?����Y<�c��j���\����c׻@i�fQy^�S�g��گ|�ש�7.9�U܀����eO�����x�����	�X0Ji����ӊ���Q�E�pŸ� <��7���f��H����h�5G��tG�w
L
U4���K>mT��U�wj�#�>_�-�Q�}"��*��TsQ�#4�]��Hky��{`�����dW�x�^�k7!|��"׌��	�7�$��{�9ќƝ�-#�(8ʄ�iѥ�<gZ��6�	��C.l^M~e@A���a�_au��t��r���� �d�~�������~��L�Q��ͩ�R1MD�g�-,��m�G�5+�!é1߱���~�k䶆1��^/C�-2|���A�X�>�e��	GM�lS�3k{�B9����4o�*1Aց27��?9�W��$z��ܛ,@3�%
渽[��_Kg6�N�����e��3� mO�G(�KTJ�!�Ŗ��J%ms�"'��s$, ])]a�Ww�e��Ѿ,���?�;� E�I\m^�m�uB�IO��4LU���\S	MnT��ғ~����|25����ݷ�0W�\5�`�IS4�|������v-V���q�>�H��U*�!�%5�=d��Nv��:뿾(+"�[�R�.O�>�7Z���Q�Ò%����ˌ�>��'�)��)%�X��ɇ$l/��r/���vi�b�e�4�A۟[��O/����b@=�)��J4l`ݴ�.,�����̡E����Ә��9g�4}I ���qT�mI�nO>�v��R79����T��|��|��*�s3�I�~Iy��{+�v��v��������m�1/
{�-;��Y�Z���&u �n��i�}f��kd�Q{ͪ��0��0�d�.��#����M=�a��~�6\�"<��H�M,O�#hѵ~qY�����v�w1�-e~˺����n)��|!�q__��B˫�{�� &+�4��uft��%1[.����>����ʆ�)&�,ɜ��[_�^���j/�	Vl�y�ݽz����z��J�U���g��2�7�8��U�k?:���)����c�B[�2ƽ������:���xI����ގO
���ȗ��^8h!禓+w�Da�?��2�;@�rM�����f�\h���w��f��T#�%6(��'4���Pv���o*�jM�Z�Y|�v��FRL=��9À�hd=H��s0Q�6�<���0�$�����F�"
/�-R���<����B;q>ҳ�a�"TTux��8��\(Q��Y��p�Z%>9T������m"m�0�8������ڡ�Z��U��2!�G�rOa����[D�q �5�Z�x��&4^U~��(�!��N�k�V�6Ya����s�^PEy��X}~��*_�j�3ڞ�q���0����+6	h&�R��#��3;�
�����WΊ���������pnŢ�n�9�����gw�$���N{�j�SCx�O��+�(�=��{?�6��|��_��M�n�}
����K	��#�1�59�k� �G�@�B�������@�\����T������֥1�H��'d! �M�B�L�2_�8��]n���1ۂY{
.@|_
g�o�5���0N�)�3����Nŧ�Fj�/6��nza��#ɀ5��~Z�������ˉa�ړ��o����q2�yڤ���3��[�	W5�YN?���!�ZW�ZR�*�����X��i����Yыݴ�}F��vv�pzX�����cy���H	���fʙ���J�`1��K꽢Fn��"��b�g��Dh�D�p��S�V��ְ��k���ե�*�J���������l��"ل���ze�E8��+E�6o�h!	�x��P��0���$������h>���t�/F����v��<�s�s���]B���ձ϶c-��v_C�&f�v)l�v�I��<P�tE|S�b~�\6�8�_Α�BX�l�nUK���U\?�-(7#<��_�7�_��u����HaT������q�*� >Y�x>�2K/y�2FE�P"�,�ԭcl}����t�S��ςZttqQ ��XPw�(YmO��I���rF2_��������]t�prl�e.�#b��Ԭ��F��ĸ�J�>	�'>�E���A���P����-5k,�������׭j�Rw�g^p6^�kE�����i�0�Yg3Tt������5�F��Rv2��{Q����l7"�|e�T[ �>�m'��i����&�?��Fɋ�p{n��Fzr1�߹�rT��΋b��]`�����ؘ(h�#c�zF�ԑf��ܩ��'��O��� ���G��k)~��8�I��?C�}qcRC!Z9*���#&��aJ�O٪d�~��G��O
@�[��T���G{�}۹���t�'I�����L����G��d�P�c
ʅ[�u9����~j�)p�x�h�����O�7`�W�&�p� E2٣��W��B��-E�
ޥ_+�o��$pp���m�P�Q�����;�ĭ}/|6Ah���XH�[�?V���$�jH�ee�U�^�Kʣ�F��0�5�zFjP�������1����,��$Mʃ�fc4Wn��x�����;�}��u���`�=��B�&y����E�a�ʪ:H���L|m����yt�\M�W72���`~\�(�C�Q$z* ݼG��Ra���	�"<��pE�-�t-w����j�ǨD��w�{�<	��!d!Υ�)�^v~)��/���e�yA]��򦡶�����<�~���C���4�Pj�P��%o�L�a� U@ĩ<��W��� �V���JO�tM���b���nv�Yt��&�e
���օ���*x�J���W<�):�	5<6;�W�B5@��9b�P�ݍ�����k�}�kH��\�U!Uoi��l�J��F�� ��)6V4��2���ŗ�+��"y�!�w�*;���i4a;�8�Z�
�j�P��j������r9������T�ӷB6(���?�+��ŕ@�kN���'��6����g�����L�吣e&UO�'s�a;��J #P*��hâ���[��di�_������l��������(��F{45俷��V�5G������<\v�=ӲV@�tY�\܈���1��F�̼�-�m�_�=\\G�{��0n�[C�H>g�C���eA�.�X�`�ӥJ���g�p��f��;*F`����$�5Q7��@ 	e�P�x�	v!o�V��i)N9��і%���z�2@�)Ljt�K��d*����W#�	H#a.tGv����+�]M჊����5�͏�'H8��&���b���x$�� K=/�� �>�^\��r|X�L�GQC�VkZ��D��6,�Ŷ�&Q�!��t�DHޞ>>|�] ȼ��5��{����	����9��_�[|��%8� ��9�Ϙ�{��e�jT�=H.�Ǡ�j�P���Z�C&��'�m��o�d�N�s�L�ƃ�?_0=}��w�:
�]Ǫ�&/Q��^���;1����{���Kn;����iн7�[�c���Ú`#mC�w�$r֐�[>MX��q5�I�Ǻ����x�d���3r	.�$=5z1!�%�!��҄��'���?#Ã�� x�{���	�W�=�խt���O�F���c�=)����*V�).5A��3�*m����*��5D�G%�܊�3C�#\��X�`˪��U�p�r�����)�4z�#7��J���],����e=�:f�_T◒k�7L)��Kk� �r�ϡ�ˬVXp���|fN�~�C����P3h�7�$}WX�T��S�����E�������8=Ut\1�[b~$�˫DΩ�.�@����}$N�[�{��[Xƥ8�F&a,��\@|�ţ�I��`����4��I,�M���(�?���a�$�.�X��"�����κI4��F�[��[����Ӟ<���*�y���{.�}����p�C�
u1�2|�mT��o�>T̋Eܜc@�3,#�l�{�D�o���ZY׈Bos��U
ޅ�.�H��Wp���,���iM$?_�������P��]�r��.������>���ͳ�kù#E�ᲈ$Oў��+�ͯ���-.���C�k��gv��g���X���?��D�����+�X��A)_K���z��X�78��.�����O�ƽ�v�ɮG��>;�Բ���pK�c@�Ϛ���<K;�� �����ջ�]&�����e�b�%5�p_�� `ږpX��AqH���n����;��J��T5�1�_S}�V�د���>���ʐd��	��ݽ$-L����O�tk�v����;�7��B�(�.��#=�[�y���/}<��yi*9�+P<�ͱ��
�y~=]��[;��j�2���E�J|7�!=��6J��~47���E�2�sM�[X���,�� >�@vg��hDU�߽�������O�z�M���P~���7��#�aR�����-s�>�&�%r���I�0�9�ۜ���$Qi�a�vmK��#��"k�"��c�����:F��Z�3ɛ�����	϶~p~s�6^�%��nZ���j���v�1��P5�j8�IbE��({�9B)S�Ѩw���q)k�K��<e��_���$�=G=c�|dC��~���
6��N�H��U���q�a���K���򏫲��/�P?�sŦ9����~ K =�ߏ���㦒�e�o1
���r�˱��ӫ�Q�y?���a:�}pML/v�|�d�mK�l����s�bY����� 5��5�F��G28J�n�Z�y��*��;�9�5�OW�:}Z�m��̌ij1�.���An�Ģ���͂��3ޅ�������Ih	;��XA��/�	r�i�C����O1�uY��/S�H�9&J�w6�`;�'�t��)�җe�d=s"�mV5e���Q�AH=�0�4�M�p:E��u���Yp�� ̫i;K%_���<t"��A���¸�[�|e@S��c� l�{+��}�?0&Ij���c��(�PlTPo.r���@0r��ҧM�8��@s�v������"]aM��b;�1��X!��:5� ���G�/�9���#_��n(�V���F��aXD�L����G̯��'r2�$�Ә�,�8^U��B�����W�r}L`!�v��R����&���`C�
L'�l���Mydݱ��Z	#B���e���<��)#�p�y�(�X0�膱���3��&��%����ƚ�6n����j�O�c8�w)����o��-�7>I�-��i����۞q=���-vK��@E�d��c���ԤD�.������V������k����B��v���C�w��R9����x�y)��l'���I�c����l�	v-Io+�L����f����B\v�1{��m��݄� O���7B��e�g����Ү��A3�i*�.s. �P�4��;G��r{[��Eqs [T�0e`�����n;C�k���4:����a���S2Q%�R���ze��9�@��\vvWvF,s'��(�AX�w ��^ٝO�m�^/Y�}E(LP��P�$r�p���ܝ����U�g��//a���>Q\8�Z��Ɓd�b��E�]W�h�{��	×�xl�ݻ����6����t�1cu}\�ݾ���כF_ѴA���֢��Tt�����\�������1:X���}�o1�g�궔�F��q'�\�A��M�HD0X��|�C��F��p�����u�����h�ќ\�}u3��(=.�)ey��,*�q�+��*e�T�a+Z����'%A�[�@�R�e�+�O����]:ǘ��?+�g�Õψ���Vq߁���0m���Y�_���1녲<O�W�|`(�3�;-Ս��e�ސ(����tX�N�1Vi�w�N�u��+w)���F*��m3�NAMB�!�.ƿ���X/�5��+���u�c/ua��=��=�$�q���QX�n\�FY���zN�_���Q��M���#�d�S��n��SFL@ºUP+����
�h�4G��Y#h�],J?��t� igKot�.�ވ`��\��'КYd�����N�ە��6����9�!�Xi\�o@K��l�HtD����j�o �k�Z���a�c��>��&ӻ�]��ȌP4dhck}b]�7�~�o��#e�tON�ztFU�0�N�톥��O���`O���-"�p�!ީ�����<���(��ѱq��2����E����2�>�"u�}�;#���~�����ʈ��#4!̍Z�^X�ￎ�9����n�'� ����`��Լ�2�� 5˱�n(s ����!���a���y�;z%�*-����X��M~��r�\�-����pKjJ�dbK�N��Tx����kj���8bԯGFs�	ABteYL�,`��0Ti�@ٲ�0�G~*�Jw��t�H�U�a�h��l� �ȫaU�A۪I���t��,BS-e�=jTd��T�+��h����N�r�kͳ\O�QJ��	�F-�!ЎO6-�G���r`ƹ|�'��R�iQ�b�4rxJd��`��]��ֺy���_:�*��T񩷵�Mɤ~W!7b}��)e: �`T�<(؀F�K����V��d��(�.���o�2?;1
��q^�f��ʸ���{��d�icS^�	=��9��è��g�k�MJz��:t�Q_��n�N~y��o�q�h Gk]���ڧM*hHLm/�a�A�ᴸʼ��G(xt@#y��Q���'�Ԥ[X;���4=�%߂��XA��$:�<xL�$��:�0܁���f>�@Wo �\}37R���C��VJ�]�je�q���s�Xk�x�	�nB(�g�!w?�޽����x���K(��
O�3`�d��&�kdﱃ���puX�5x��T��X��gk�ޡg8û�w໰�*���� �;��=�g"9�(�CM�u;��C�q���@�����n$DE�����R��5��U�b��D*0pےb{Ơ��bDe����\�d���h~��{��U����몥�������d���q���p1R��BWp��7a?Gb�Ӻ1�5&E�F���e�|�:O����(ͤƒ�E�U���z�:�*�F
�C���dod���>�M������
G[S�hK�b�Of�-�g%��KZ<v� ��6?����oA���G |��1�R�{�_��c�1n���~�L��TMg�*�b�v
���F�^F��ʿ�Q�b�=
� ��b�8�+d�iǉ�'�Ժs�Ot�E)�,����6��Ď��u��0�V���k�1M�6��	��U�Q��SL�kX�hM����\_�S�XM��7��'Ֆ��Ru�R3�ke薐A�@1���ۗ{�Z�UI,o*?$��]���B2��}�S�R���o����<����v�������n+�W� �&�9��C����R�(%_����x��c	�}!�w��My��Ӌ�?X�,����C^� JF���u�{�!�M�V��J傺!�+AZ�PW�R[�Y���[�j%P�xRm7� �6�����7��n=��"����$m	av7V]��n��{�����2k߯c얊��S�%�m�^�������R�b��6m}�f���- �ӥ'0+�|�w�����������|,�v�A㢫e��dțZ^NK��A�$���F���xV� zRU�>W>$�i�G�oOH�Ѥ>���<��$:[&�4�*��s8��1��&��X<UB����>񶯞ƌ�Q��i6�ٹ_�~����PIX�(&`���g�MY2�?I���"%9�Cg8WC��6�'2�>x�a�&�l,�O���V/�*`����դ�/� �)�':� {��M��f�BXu�p�Qʑ�x�y�*��ε���{�F������% �7�ҁ&u�x#(��Q��]�wT롼�>	�,�v��pY�g�K�z�r�TT�^��2h�E}�J�:X�4���ϥ��J�'?"���$��N�X<�êXvY���m�\��N_7M�߲����'=���{aW�!�LK��ޥ�<=:��r5H��t��Ӂ�F��T,1�"�T��2��a0��";I>�E6�Cu]���0QD�*�}�ޤRDt~�^&\��ط{u"��.M�\��W�x���c'R�i�_� l�:��8?7 �=q8�<��^b�J^h�Jϒ�f�4B��ӎ$��p���X^]`Ո��N,�3U^,�7"��m�sd>��B�J��}�a�Ӻ�����*h�
EX�1Rgm^�sQ��H���c��>;7�t�ݝ[�3)?6��?z�:|����m��f=���\F�\�[/SS8x�\x�g'��{����.ʮ b�LWM�4R���&a�q�{�Z�즩�-���;Zs��LK޳��s!���J{��L�x7~6߰���������)U�� ��>X[�g��Tzw�l8��&�@����£,�r�xaqJ�\�ȟj�q%8�x�?"x��1~�Ӻ[�\F,aQ�����4�rq�ӓa��d�Щᐿ��CM�$N=�N{s��Y��D���W�A0�O�2З����F��B�R&/B�F,'�e�z�$�-4̎�0d���'m��
!��e<3T�`���@�����K���:�CA��qtB^3K��Q�*��S#gj�E�P�2�ڐv�]�?���I���"�c�p	���*�r\��ح_ oY}6�78-�/���{�:�j�K۝��c�мA 7���ٟ�Q��lDu�H������J�������U4
۸]�D3��G���h�D���:/Ls��+�);S$�e��j�����^����_� ���f-'��L��iw6e��Fw�\�;y	�gm�&��o$q�pۿ�F\{�T�h댱oꄔ@/(9Ϋ�wr�P�B������u��� ��x��,~�t��C޴>>���0�N� j�ũ�rpF7��SaZ�˳���(�>(-���g�������*��om�'2~>�1%Dq.g�
&x.t��Ԛyx�#bI�v���� ��E��5z�?.m��Cpa���p*��j�Z����g^z`]��x�ygxT�9�v��\��֒��Ր�C�gqU�yAKb0�Ȑ
��M�Q�&�w����Vr��jxq"��Nt��b���X[��&b�<Ή8�{��O)���w#qj��pk1m������6Ӻ����؎�'�O��|PWװ��v�awR���WO�]�#���ҭ�H�~�?�y���2Z�NL�g��� N�������@���hY��f�Xi��%\�Q~�x��V������V��[+�2���L������_����?;��۲����$J�W��F8�� �/�_V��`�����=T���*X�1T�`�/5s_��c�&�~�92��������l_�?S������>����f���&M^Q�u�D��Z��7Sfν\���`��0h�3�h]=�M�lG��i�aJ;m�3.�EV٨<�N�4[��	Cyflt��N��́�t�h׈����O��|M�%A�]�;��+�� Y}Ȟ�@���tm7�[�Ge^\�2����I/����V)���D���m�����mn�����I{C��qFj�����ঢb�[^1��vuu���^d\Ȅ�=�g��&�����hx�G��O���C��I&����>*̠��L�Ii.C�*5�6�����烱l{h1���&�r�&�kH�/��Ζ��S:�p��?f�݁���ANH��2z��H���=9����L����}�%��!3�."s�_8���	��.K��R�LIg�&�
E%/�<;��A�P�j��=;t̏� 1�6l���'RU���N�J<��@�z8��	��zSb�'����闍��Gz��y|`��?�ơy囓g�td%H��u�}L�P������;����E��(��'b��v��~����&o*�K]?���)L'���� �Ɑw��*�����r��g��8�Md��6]O�jo��*�(�"�mU6[�@���>FZ���>?�P!�s$��F��B�9�s-'�U�v	��0� iړMm`��YTy��u:�3�$c�0��7�Ln����7������"��Kh|�^:��r8�愛x$�a(�nL{��ӌ�?�����F��~�)��~�8�oHSs�����dl�J�Z�90̓���Z���&<ߛ+�4�V[d|U�޿Qxc2����M24U(�W}j�N��p���ʐ�K^Za.�R=L�d'��o�]y���-�	���x��!řJN��p��/��!6�^��/?G��=�P���ؼv�F��~W���$�ӊ�'�wg��n��Δ���w�"$e��1��<g�4��%�~P��n���ޕ�W�� ��/�=��˖_����
<�n٪�{]�τ�TaZ��Z<��LWzn%�;?19`�s:5!C�ꄁa��#�Ew��������(��d�NNڅ�Q��/oKEJd�
���׻><�qe��<�MP��a�����͘�h�6�-4�EM}؆�g�=��Ӄ	OΤF��M+�G��&Dk����N��g�p	�Qg�"�.Z�.��7����&����n?�T�.ְQ#�Dmݶ[�2Nem��S�uU�Vhbܹ_��39�9����s��>8RDgHj��O\*������9sxP���I$��;x��2�ދ|sی��U�r=��(i�=�.;����_U���=���h����[�>��;X�ap%��+<7
o�9W5�2ߞ���e6y�,�����mq$n�h��݃ftY�#�KPq���vDMM�sY��H�a��HwV �z�|�)e�I��_h��a9.3_������i�17y�g���R�]�f�΅ K�}V}X�&s,mYǡ���c�4��G@N�gd��E,������d����EgI��P8H珳ā�C��@j�I /�\���X�3&��;���;z���Pgr�0��e��w���X�'�Ҏ���t�������r$Id,��Nw�%^0���	o��fL��r�tAPƴ�K�Q��,\Wח'?�;NsGr!��Ă��;�&�H6R�@g�e|�#e��\�tܟQ��v����w$�3d=�/"�zL�KJ�b�[∳I��с ���X���	T^������*"-\�����+(Q�و+��Y�xj�����H+��t/^b+�1�(��^�C�"�e��JJn^)���Ac��W!fy����ˊ��>���<�,�^����,|��ܥh:(/hO�O	���>E���*d��8�$>� X����n:s�DA��4ɩ�ꁊ�M��.D��A��W�ʌ�f�+k�0��w1c��2ia߆5���RZ�$��O���N�i�`!]��� #p�_QYDcq�^p���0�v�\�e�f�a����1�Z�'�U"Üէߦ,@x�T���_{�7�x�J?#��N=���hc��SWPЌ%��qW;tgF�p��A!�B�T�ҹ}&,BX��]S��F@ic��|��\���Waď�&�p�A�N}��-�������K�xCW���$����.mi�R�=�ߢ���8����+��Cނ�鄦ȱ����q����� z�ˤ�!*��V�Ǐ�	VX�<ެz�N R�<��-���M��7EAk-��bh��o@�%|�o���r[?E1����),��GYdtf$��x��Z��D�^��S��O{38M�R� Q�^���!��p�d�*�Bs	���+�Q��<e׿ �b����B����w  �
��ɳ1���wH�gB�
-��"`��72��!��p�Bc2���f��U��c����[������_���e"a�=�]�Y!U��L�>N+��Y8�`��bu5���B�Ua7���Sk<a�	��?��-�#z5���\{dQٔ�?�3��s��_`�q�D�J�EQ.]C������H�o�����&�9��D���sZy4c��/lJ����9j�������2��6�)�+��{��*� 5�W�Wf:�Z������g����I�-y�Eh���0�^u��^�e��e`��F�|x.��#@2wA��x޴�N��H>>j͗R<N j�~|����1����{ӂ�Y����<�`��0=�-���Ak��nF��;a���4h�����6oP��pj�8����׳�Ea>vXm~����F5s$f	l�B�/����"�s���GI�s�B��3R�ڲ��m\l��N� +�l�5~:ҮʬR��c��=���&s��m�f����䣥�[3��f�K�L>O��R9J#m�e�JS�b�������*�w��~�}�$)!f������b���=~���d���Ia���*S�m�1i����nI%��/�l���*����$,�GIǔ:����7u�L��C����3-� cȍ��Y1(�/�?Ɲ^��xd��XBM5>���0���&�K& {ݑ[��@��� 3��^V��m��-7`w����lG�������j���@_�L�`���ֽ�~kQ�����5�>Qy@@�>��œ��Ds����-����*����V�+L��P�ih2S�zxs�[H���������,hU��@�غ���Q��]p,w��>OP��,��܍��X�,W�r�#&(����U G��-���|��Y�R#�5@� ��4K-͌|.c�Y;���9�mЯ�� �7`�+?`6N��P��}�Ū�vil�^�K��D�(�U 7v�c������Ņ��H>�U� �+�Z8�M=�1�e/�о=�B]tJgS��#1*I�g��k���n��hQ<e�}}YMh��c*;s��K���2���D�ıU\c��9lH��Z���w�_l�1H��\���jѡ�3�g���n�'Կ����T���VX%-`"��^ v�Qz1�-W���� �M*�l�2�n߁�=�>�<�ak��x�~��v'�Q[y?5�f�f��yky
��[�yи���Z�$|=��� a�kRM|%�mA
،�/��cZ�-d���)bb9#I�`�s<q�[���4�_hS ;9���A�tJ�0�~S��^�G���Q�����l�z�'�M����U����y���>hWh�������Z]we�^�i�N�������t_�ѫs�R��G'}e1��X���^��o��O�=���n͈T�j�H��,�1J�'�+���q�p�H-}�q�;Qh9���:��0�J$��w<qa4f˥�?��i]J�"���7�唯��^��{�J�J~Kzà��L�P��U�:�Bk�jk�����°�M�H
���E$1͙�T����ʫ��_�h������L=g����_�HyU�"��˜���ؑ�$`%�?�G�U�S흫��U�!O�ڒlv���
A�n����Z 7 W]娅�O錕�]��N�w�(����[��'�a��Aֽ���ij;d���ۀ|��u�GK��8)��j���ޒ���!��`n0�h]o�9~�%'46�72\�$F0�-:0��u��T�����KFQK��Z�%��j��si)��������1�8�����3����Fe���)��Y9p<�v�cKD��ޕ4���$�9��#����۸��	��*���jr������e��a�b����[ǀa�ܺ���O�j�D�=򜓂F�]��&Τ�郺d��f��y�(��II/�w7!y���t7��ş��|�&����͹r9��\%���H�z��,��=�f+�gU(�ϼ�3D���L�[0_�a'@����Ѝ���g� �����
zp0��U�n��SۤD�m\AL|][��!h��5�[��˲cq�(X�g�.�Iޑ3���C�(r��r�{@*���*):�:z&"������hp����vCq��Og����⠚�� *��M+G|�!ʜ.���n`@m�V0	y�<�`o��!�vg��󎙜�&A�a�����hWtP�{� 87���F�l��xaQi6L�� &���ɟ;��j��l�nZ�E�k�`_dX����:�t�eWPJ�o�bf��Ӹ���Ih�OR[�#Љ�O;�2�n�"��ٻ���B��t,� ͸7mn�Q��,޹���$��>b�lE[�����W����WGP���m&�;@���Q��41��^�o�����T Z�N3Ic��[��f��tK��G�߸��R���'�D-z�:��")�����w	���FV��[Z9rq3��A���?LЬC3�j��n�hv�X�&?VK���ȕM[34M��:��P�j���L����X�������^�^-���I�ina���e�g4��pg,�@UP� �jU9)���7~;��ߢ�SN̿���z�W��[��D�*	u��D���^FMVj]מ}�KnR=4��^L�#��"Xz��O����YjG�.���~��@?�g��4�w1��N��0SS!�?䀱>����#�
S��7����"e���."?E9�s���Z����\f�_-�s������H�d}<�`�[��h�:c��p�u�M���N�m�R���� � C��]��g(�Cb@f���@5|?�d2���C�e��S��ߌ?����V�������>��.x�'-a�N͛��wW-�����|�d��^��0VW��y�3K��P2$ET5(�"kB)������ �x�*�+�y^6�H�����2�y�nM�[���
�)?�s~�	E����4���E���bp�����iq?)H\��E���F^��E�X=���-3וӖ�d�9�N�BE:	Z\!�3!Y��2�15ص0+����XY�EU@~l���j�&���L����U��E��vүh�|�Ơ{�w�]Ș7��v�߷r��%֮�u�;���N؎ �Ax�/��<m;Xw�_�Tg�e.��My��B�r9��|7#83���'m��v���οq~�kkh�/O�b-�^� 硃A��b̄F@��v�Ȕ=��Sm�N�V��<���9����{H'���мs?�sB?��h�?���wR�8!��FW� ]��o�Mw�͐��l�yu5�����H����Gm�Xf�j��ze�|��Q���ɝ,8�e��������p�@
��Z����P\T��ƫ��Ц���L�P>��D�>�;�e����R4=���/8.�pLr����A�嘜���vN�xW�J�����������#��hMhP��t��}�z������W�/��'ǁ/��b�F2yC�3Sa���Mc��Nkg��(��+�R�����,qz�Mln�t ߈:��ťijT%P�!z�����6��>M0�/b���Rm�c8�2�>��j���*��sy~k��$G�,�|l�C�@��x80����!��&�g�%.� >-7�WpXR�5W:���	��*v���#�}�O�h������Մ.x�F���f�����@m�pJ)�wI�ɤ��!�!8��ת����;^{�l8�����H�]?pk�c�y���4�]6����z�ӌᲸ���b.��a>����
���P�n|a�Xqe(�;��+
W�U1c���$�Bm�A������G��V��w�0Vg]�ۥ���iX�n��TwQ�����m\=�R��I���q����,�</���'����MS8�{	x�P�?>0�r�Ĳ��JS������M�fu)���^���k=�nz_�b����u�ʂ�i��$����*	f�(u�=�EI̸dD����^Ʊ�ڜ6}�ʭM��l<q��[�KNF�|� ��$@7�I;��g8�I�Y,���6ٵ|0z���=qn:�I��ʗ@�F1uG��W�t����ӸȂ3��>�j���P�����&ffy��.e6G^�kҸ��Z^@�荼^�L�3��/���j�x�h�P7�$*�����O�|��v9��2U���l�=��F]v�F'�vM
��`3ŭ��sEymyS������$v� C�$5(-~�@y5!�l��@����%�~�U�!�k)^�'Г�����Q�|�"Q��=�� �t�������^竧�����d�&����V2����3�2��۰m�4�G���0�$'nn�W��fb�G�jb6:�X��+���!kT��0U*���vӸv�n�§1���Z�x�!��8��U*cM��KNhTk*'���>]��o��b�z�u�idX�ˋ{�����&|��m���-T��Ao�2�fָ���O�/�i���c��gN����DCg5=aܕ���[�s�ML�s���J����ǎUx�1�S�M�g��j���-��B��U?dOg���z�����>j�����i��k��Ւ؇f	�Oδ.>���<���ԫ3����g�����Yq����c���!خZ��k�#15�/�l$p��Ha?���w�gqf�Uz(�f�*��܏�2�����[+_���|��&�C��Q�MOˏ�WRd�*�3�F�g�������3�6�����"�L�b>NtM��)bϓ�/U�0�Z�Y=�Q��#>	z��<U�$Q�55��J�X���]�GM�5>�b����83��
��W�t=#�:���Q'��KD���	���a���������c�o�U�F	���<r�����L�O}'|�Gͮs��]i�n����T��ZA�`�=�'囩�~�-AAP�{ ٻmY��6��[�����(�|P��s���zi&#B
h*RkP�ݕ����A�a�)k��z�*ʣ��t1��a��7�E�Hݵ��г�5�HI��z�벂�bp�?R�X_�h���9��@&�#�:��,���� �_'�1ͥ+Y�ߋ	�`��7�)�S2�4���)N���G�R%�FJ�6>�.�cW��q.��]�8�^L��	æw�6E���a5���j����||@N����qÎL�Z�.�z�IG?s�;���EZ�_�I���no�}N�B�j�
2vC�++��ɂ �^V��'%� �Q���-4]�{̽��rO���s����Es��8-��S�m���_�]�k �q�}V ��xO�#�3�@["��Y��Ӛ�\��o��.*� ��Н��7�ftԚ��؞�bc=5K�&����\A����³��8�g3�B���18��F>h��*��_�����ō�\?���p����.���8�1d.j��Ⱦn�ԕf�g}�Yf� �'��DQ�1W�Q��4���M(��v[���Q9�`��Ґ���'%�<�N	�M�k,z��~�V��[�Q���<��%w����) ZN���5d�'�Fhw��?^���5��80%�(���4g>���g�/��I�6���e.P�=GD�n2��3.XB�u�"�S�����_�CQ"Hf'5�V��1��	��e�O>�%z�|��.��*�=���baoO	ؽ�����+<K�Q�(A��*��Hb�5��]�C誤�
���W-n;��/�aO�7�YB�k[��B��-1����+����[��ؗV�W�!�+�!'�_�o1G��	!p�Rs?�a�)8Q���ŀu/����`�� �!����,��v"��0�%Y�VK���uYn����^�!ڴ;7i٣����mcq�2ԧ/���cv�В�	De�J«�L���2'��|I���B?�Ȧ=�`�h�>N\�691a���~UL�p�G�[�"�c��*7gb�r�f"ik���a;WG*��&Nآ*�Q�@�`���*�V��Lϫ��q�ϐ�gU���^��D�V���s�����0����+m0��x�GINRn����^����i��=�ͱT�G�6�g���R��[��9���K/z8r�d��_y����9q��K��|bJ����y�'|��BP���I?԰L*��H���+���rRU��\��+/�'�)b@��U8fK>����Vm;Eә!��jr�[���m-���u�w��#ɩF�Xc�ZS�Y���EI��
P��c�_� �S�{���w]�������<���C��ϻ(]LR�4�U��Sm_��fx�՚���o�Ԃ1H4�����,��0��[.���O�t_�n�V�12�)��`>�}��Vګ}����'*�rp���0D�@��M>5����^�f�*@15�#O�g�^�I��Ç� 6R�y7X�?�}~�Oўk���[
)�:�
�;bS������s�����.��I����V;	PvQj���+�4Ka���Nd�ƈ����Ԭ�%<u@-߽�j$���o��ՐϜ���ٛ�!Z�J[���Ǽ6o_V����_0[��S�8��y3��I�ҙ�Xҗ�:���v��p�4\�ꬍ2f�2�2�R"��q֝�F&-���: ��O2cd���e �S[pKE7R�a���guK���ȕ=�����e�mo�ZN9�w��r����,�B�&�m=e��*��V�Ϻ[ҼD�p �E���F��TK�z�l6�W�@fKo<�@�u�wr������Z���yt���n0ST��`�y183���X �HD�x0w�ܝ�0��1�������p@/W8���;�E����P�ͻ�t��3��5&�A��A��� ����0D�s�����:W{��h��u9�j�K/Z��uC�%�S�-כ`���n�(UJ�n�nNS�v[�Fr#�����z��L���`���f������+�?�&\^/�g�Zj֧1reN��?C�`����IA���ܠJ�팢F�����t�e�Y�.��ɡ^F�G�&������ZV����Z����^�<p�a���'Yg��}U��B���Z��P�3D��g��5$>Ex�>����4tG��� G�����]zk��~U���]ʁXm��p�kV��ae�9�#�FM�V�Bؕ�F��T8���|LGC�L�F��!3<��{%�x���9%NMV1E\B����~V�FDũ�$��s1����B�%ɵ�z&1Gx1�L��ԑ9�)`�/��k�)�~�A^`:A�y!�xAڪ��͡eyZ9�K�X�w9Xl�o��ю��*ǕK�ʯ�'/#zz��R�H{	U@9�6�X�*�_��a�|�8{7��p�=H|}�I�p��X��4�,4���2��S]��@_}����%�ݴ�j�2Ua)�2�|l�#`�03�U�'�2*U��9?d�U�Zj'|]M׆�$��쥼���$�z���?f!���	�o����Wx��U ��� a���L��mr=�w>o-���������?�{��Sj�7	�샓��Ms��k,�p���X�+�L���Fb�}��'򷐙�<���BU��-�n*zE~�
���"P���٦�`c� fƪ��9)9��B���fzɥD��:��I-�O�2m��h�-�@�cn��Ĵ�z�g��s��ƿ�*:�A�I�5��1[���Ƙ��ܶ��e�j*i
Fa�$H 	1$!
����pC\�0�;�{L7���MG��H/�k�ө2ѧ�}i�����0�,`��Agڣ��&�!~�NIk!���.#��ҋdI#�)���SC%e��r�h$�|SX�c�BT}Qn	�衤U�[ pV�P"P<�+�w���Nfݖ�_�Ux�q�������uKZ������;sv�.������E��[&d	]�t�
P�B�E�綀�A�j@���p��"퓍��ÃX���ǜ�V4R�p^���m_2ƴA;T�G��F�.�'޹�=Hk��Ix���p�4�������1�L��wiƜ�Q�����p�r&�m�}��)֡���w4���U��^E���\-�xG��Ğ+�D�qӪ�p�|}�j[�K�w4�4Qc����]����f?&v�Na;!��pd�I^�E���l�&W3���x���kU�{�fZ�8M�߿�L��(΢B�x"!3�y���@{U��{�a!K�1{��&��:�@�Α�1bK2x��;<�&s ;�6���	����;1�i$\�EI������n]�1b�����k�b��L�����Y>1)F?R#D���xط�O$�a��+�QF�i�B��=ts��8��Q�K�-��l��e���|**(�M����Yn��GH��U��\8EBӞ����K���JF�����
f���+�Z��s��B��['̑n��7��s"�
b�4��O �F��f0*��R��j�Wg�p	Y��!�I�6��'|�k�dޱ���=�SCV��Ğ�B�ݥw�������u��Ӥۧڎ�Q�^����P涞s��>��;F�㛥5�n�֜L��/��~���oU��z�y���q�f��O��C�q�6(%���^����-�3�n�n�IE%���>/A! a]E�PU�tc>�n�
���M�yA�9�,�Ϋx�$�|o@�i%�H��Ek]�P�&�Y���z0�È�[Χ��b��7�R��ï�-����a��@��3Jy���#�>�"*\)+\�-G@���氀��e\��%��g(53�!W��g�r�ӓ��H������I4�+5��UF,�i��lЭ$��'��W-���jx_�� z-G{�-����kM����n�4�X+S�u�P���j��|�R�PO$!���ֶ��Zu�C��T� #�0A8AȢ��\�]��a�'[�.����s�fD����)-=m��3�m�z��G��`y��	�~c4[P�YzuZ�3[��)F"��_I��y)�~o���uzhK�5�Le������_mv�Ev� �[ʏ�$��s>�H�A�S;����O��������;&��+��ؐ0�^�Of��of�B� �Ƀ��
{rS_`���(?#��7�w�_`�MH# 7��i8_޸k0�;0�\5۝&`.6�o(��R˱���땰'����j��6d��z�6U�><<�ACr'#��rm\X�@�U����K(�7[�$�*�߰�T����z��0��x��챀i��)���^?~�ń-eʥ�G�t6c���-awߧ5��T:�0�8��}O��#V�Px�P��*k��
�y��R���(��ȥ�WV�+�Ͽ�2����Q��x0H���Q�yay]�B�$�룔��;j���Bڟ� ���aRϢ1�?�Ux�%^���l��*���m&Î"���l���sL��s23m�)Js0Ěy�t�Nw$���e]�]�hIڠ��FV5υ�03܂�Z�GTȕ<N#����a�/8P�^�t��Y���]�}x�d�-	�$?!@j�1�P'�/z��^���n��v�s"Ϫ,-SK؏ə�	[�#>Ki�f�IC�)M�+�;�ѴeL�v�;@��1D����YdWC��1rJ��<d�؆�B����;nF��=��hX�o�8|�C��D�E��J�-,av\�t��_|Y�F�H�*�����;�r��{� K���N';w�l+���$��cqN�_��o��:�VpP�t4v0*���x-	;�@B<I�#�� ƜC3QLA�a��-����T��F�� ���2{K�M���ޔ�$s�9|��c�~|1o�t�%�k؛�0-v�NW����DzȠՎ�u~x�������@��4���
Kr�V��ҙ���U\��r�U�͟���Ǭ�x$!L�q��=�;8��(4���#��$z"Ф��'�*��ޕ����m��������X�s�*<>�֓�,�x�����/TKM�R�#��k��������?(�3D��i:�O[F3�Ɠ��H����
Ǻ���7]��pЏ�����2]۔݉���t4a�0s}��OD��R_�=�����E,A}�4��T��/P�^q�K��a��/��R`D����iMyo��.W���i]�k���������I��A��Tg5��G�(��r�s�;�܀v�J�Ϩ���o�+o����&*9�����ǯZL_��dh��������o���;���*�=���Y�DN����\�I�"eM1���d��ذ�E�K�-�����bk+�&~��]�_k��w-����쫆��n����ab��LbSp�Y�W2� -��o�>�j�%*X�Б�6_J�
r~��78��3aF� 
�<�����d�3�*��
��e�kA�0R�&�F�Ԥ��d�[������<9��,�v|B��l��l��l!ŏ�
CA�� �5���~����<�tn�G	6q�G���[�b�6-��\�l:+���}w�#xً�(U_
J_~�0����:p��k%,��.؏�TWWl�v��<7I�Ćd�.����Q��E���	�U�h����l�Ωn��)%���<�����'8ڲ�;� a�x��� \����C�>g��p��@ʨ�>:d�A)]

�Z!gB��<���A6.���R��޲e� ��_\���t�ն�x��TA�>��y����!��w����%Ω���<]�  ��\y�Ê��>��$�_(q��Q������%����T�����
�e�1oR֮
	��U�H;��8~݌&x8qY���~��o��;�1��衬C�n�?Z�e4��*�6̹�2�qݕY���v���M�.����y�̃pA��7�,��G�A @��k��v]x�E��f�����%���\ փ��=�㭩�5���P���s��
u���1��}�����$�f;�u�`�����>[�f9{YR<`�.�=.Q��a�os&��nWl�W��K�m�jF���A����-�M�b���@Fٌ�k�Nm.&����hV��uâ�@w��)^ �=j�\X ^���Uy3if�i|O������T#�K�z�����z�e+�ɧR�_eHs3G�u�:�}��[D�����GU{H�p��⨱
��Jw�^�4��G:)�H��N�,�V(RL?~lڝ�-�O�7��)��T����ާ�����gV�N]��}G%Q������}�ǜ�7{�ø�A��Czq��w	��[4��_�[+�1M�Mt�c:�4=\zoJ�s��U7�g"ўQ�"VI��\u͆8&^,�O�6RUoZ6�C?�ܐ��˄F�@������/�.���r�����)�����ݯݴm��{�I�mC%�Ue���t/E|�,=�48�r/wK�����J�}h�%�2�VԸO,�j�r�K�mM����.-&x��P�a�u��92�eaM�*6��U2�~@�:���c�3�b�-��$�FA�vBB�f���]D*�|�4�n13�%5MW���ډ�"�Y��^x��a:���1�����J`�bZ?5��	�ȇ'�,�4,��y�N���Je�_:֍�N��l�5��M{#���݄JO�� ���x"�CJs��s ���}��H@�.��Zԧ#�#I�c����$��>��@�%�X.JD2��r::�����F{=ZW�s��ߓ\SQ6��J��T+��Qx�F�+�+��|
�XB��	�f���4�Gp�UVk�S.��}r�B1}��t����O��ȉ��b]�Jx�6$���{���}|Bw�̄|��U
T�m�C3{�9d�������V�ʏ��*�ʉ���x�h��y�)�o����Q��I�?��݄u��;�6|;��l�T<+_�n\�(n�9���x(��#~�����`��vȭ� }�6e�;�4e�e$\"7�vG�6L��f�3��n <jT�G�U��C�7
��M�ۻ�z��UBm�ǘ2`T{ς�D�Aڤ�.�o�!�F�Lh��4h�@����?Hǋ�u6��lq+�Mvg�$�¨T���zl�%*6����
V�-J��J&]`t�F��W�u;}9ĨB������2x�ʥs�H��i��qVu>�Ƀ`{�Z+�a�aƇ\�Ne��/�0��v���'h���3�"6L�X*�}+�l�4p�܋�{����w�u�8"y���5���>��Sb��n�i��7\��F�pd��;�[w�*���4;��u��'���t";�>���l���r����,r7:��y�d�/9"����aY(�@"�C�6<�	��mk"Y��]�����&�*�o���Z�宬K4+��Ir/e�Ǻ� t,�L� ni���r�?�ZR$�*jdŞ��;E!�[�5��fW�(�V�`V�9�:Uϣ9+����t u����_1!�p\U�l'����B��h���a�N�R�n�1f�)�Y��9[Cgc���gX�>]��۹�9Y2ו��������Ar�u˥��z�*-/S�?J�:i���T�c�G���y�ET�y�4v�et��iQ��:ٙ����Xͅ� �H,�P��r�m9��-��c�a+۪v�s͌G�T'iqZ���aKj��6>;���q$���/�ʗ"?�@BG;��s�����``��0�N���P�%����bw�n��S��1��T�
5u&i�$9c�U�.�Z����>���.:2�+Д�ߑ:Hb�q��҆�i�9�JG��.��S�!��c�/S�qϛ�.,Fq�z�,��6���a�$�Jun(�	���y�}��o�b w�?_�k,��KM�Qs�"7��ԟN�"K_ҹ=VO�AdT��ؖr��'X�������`;g�3 ��v��;Q�9q��:H�,����ݣ@F#g��L¬�:A��4иw�?b��s[�௝9E�U���6�L�F�KH\j�������v��S&a%�g�$[���Qc�P�'��U2,�)jS��U��lu��>ݫm3M�н�b�8�3��	�Zs�F9��{hE_,9�g��C��"_���yǯ�gQ�6|��:Ԣ�rTOWg��X^�Ѹ�����ɥs�D3(1�4,�(��GK���G**5�W^ZJ����N�}D�h���F!l�]��TEL��x�:�V��-d?3c�8��w83�_�������pC�7�n6�YO5� pR�=K��F�" Pb�Q��<>���/`���q�)�z����q|�?m��&���ȩ���9[F���\�6ý�c���|Ǧ�p���%� we���s�����e�����	�;����2y��d_:���#	�-�I#�C�v,�#0�r���%�tߔ�՝o �BԆ��Fw��~5('Z����S�kK���$�E�ӛV��/d򫟩��N�Y;�T3j�F�U.�}����v���M
JJ�+Ҁ-��M�s[�5����.�>�D~3HD�C���&:7�j�s�y��ϛ59gD�7e��+� ��)���EG�c�6q��EDLG��6f�"�����㧕�4׮'����9Y�j�.��J7�Cs1䂪�K��)��nK��G&�2?8R��Rp�J9���7�ӷ#�K��q�k|�a��X\V�����t���T��Y�egX�C�|�`O �\�$z5~M�_�H���NZP �(���F�jq��	�؇7Չx ��� K@ʊ��~ L;#BD��0[p@ʍz?VL��L�Z�md^�'���~
&��F	٫�[���N�1©�/�
ᝋ@!��Z����D�����=�hy��l�))�j��Q�CT���Y޾ۂBRF��r�_�n#X떸�M,3�X��s�@&['2�QB�{ ���"R����/��"/�tW�R�ӈ�y���P:Z��"�`�D�x��Y��Q��<ԉHm��eL�M`��>#dT��ծ3��xw�b�����IB��@`l��)��L�F=r�4�~�c%���t.�����qBϣ/pfy���Iȏʰ�oɖS�&�O�	v��҈j��ߗ�J�������e�^�M�Pz�7�D�:�6X��^�Ju^�P��r������-��v7W�]=���N�eV�i�&�����z�z��@U��R.�@�|��>�h��wTJ=�!6�M��$��N��$�31?�3f�Z���n�.ѝd�*.�`�T�_Q��Iwu��U��k4��Y�v�����礪������O���gl��=27O,m��U4}�t�z�Ѝ-��e�wlȵ�]��[q�!}�kz�7���KPX<����]���Z��ԈG�/���e]�-�b�Ԧ�R$�0{$~�MI`�uBw�=�=!�<׻w�r����H˷��ªan�<�����P+�M���w	f̵yRt=A�Y�{LSf�
5����32��iU&5KG<����F����D�����h�H�e6�B��e+Jt �N�z�0�,��(�S�y�RK��c����jQ���]�%E;k�|R���T[t&*	Em.�����^B�<��F�dՑE��R�����I;飹U��1WR�S� �N6�Z��Y��c��E���:�N�~�Q�lwA"�x&�&��pw����\Z�ܟ7zS���F�PJ�WBm��,�l�1�!��/�V���,���R�fo�K�]D����
��	���)�t�6m��v��6A}��+Lm�F�`�����V!`e��a-�a^(J e�Q��|������l�oW���lJN�1�Nؽ+ `�N��c�7;�y�t�6A9O�{Ӳd��~U<�'2 7!�i|7�4h*j���Ga����d������1��|M��\�~I�pʵ��4���E}k�����;��F��j�λ#��$��mE�F�9'AA��5b�G�_���71��L#��M,�H�E�jC�w1!�S9�y^�=,Ą�G���t���(	���Dux��S�\�ד|Y��$�Z8ޘR�/����04�d 5�]e�*0{V�a�&2��D*ǋ����o��s��!�r�"-����x�����V�J���X}wu��Ժw�����z�/?{(j�/j�}��÷T�����K�ύ*��P�޹^��N�m��@E-�ѡ�S�A�n�$���]>��{R�n0�2/���3iuk����F����i����q#�⛬�j�&Ni(z_g������J�>���B�;2��Ԍ|o����R�,��o^$�r�4X^)�=X����+��*2cI�B`�1�m��k����`�����s����*����~J>�;�D�������^�������O65{��0@�P�j�kh촸�����A
�@�Ei��8����\F�:V�޿X�)���N�UfNm��1P����L�D�a4���uE#��B �$ɋ�#ȫ��d�0}]~��-�����u��s���k�i�MC���ѭX�Q�_T=/���/l���(\�E��4�{�<�t^���Mz���H�G��
}i�eF.��Dn�B�1>��[�U�4#��݃��|Wb�)J1hOL�R��T�{
/�'�t�S.�?{4�����2s�u̝�1/�Mk.��-b��k�8B	B��i��(;�F�C��Tڿ)����Π�X�s�ռ_z�@	z�0/!�}�*x�?LI�<쪭��$�i�u�ܠS�'�*GR!�A������Unr�F�g�n���}� ��)&��M�?@^8�H��,;$�㑟�39}Q�&~��)|���]"xX�0���y{i!��TF���X�
mj^m�zW0~,3ȣ�XB�!u^A,.���5�����Ex{TX���g���Ә��n�kk��۶�M(�����?hH��W�
��7'����sr��y��D�9���sB쾜�FfH������<I�ω�l�ޡ���z��M�~ϲc�A��ij��?�.�,�+�ҧ�A���E:�m�%�b�U�+0<�F��kT���#��d��u���q��X��W�� Q־�4@�oA{^cBp��M8*z��$�������v�/����� ������g䤓����M�S@%w�YGg<�4�ywP�y��3G��Y&��:L>
$�5��UYx��T���_��>K��[�D8b�0 ���Qs���E_�J0��P�u��&7e,k똛�j������ˊk�*
UicՄ�a��(,�c˅���SJ8����)��l&��`1�OȀ7ɳ��Ҁ�� (1�5\�p���{�ڡ�lZ��T||'9+����2L�rʌ=�F_�:�=b������q�G�_���F���/���D����@��I9���z�a���N�$EG~�?�o�')L6	�����1�h�,�k���V�-�I�V��9{LGN�P	��c�+#��rF_�*��Fʴ�&��u�6�#���r���Z N��X��:=�\GF��N�k̽ �MJ���g�ak��jX����j��Ò���S��#!��ϠӀ���`
(�
�#w�]���)�����ʄ��I�:V뗅�$]G���4��.(Gp�kB���2��m��6�m��-�*�܏����:����g#�'�2��4��g��g 7���0'�8j�gp���%�Tj�pf?�sMw�mlnLd�v���:s�c&1�dq�z}�?yF������r��m|��*�4r��ߺ�z�_��IK�õ�g�� �&N�B}�k�8��1�I�U�;ӎ���g�b5K����^��S���}Ղ�@�%J������u9!asjkTe�׋���8�D�ծ\��?�H�Z���A;��1�|RWw���k��&�ġ# XD4�ι�aY���C�]�G�H��+�z���c睟9�XX]b�� � @!p<Ĉ5U�F6*%?gQp���΅:��A���.  ({��)H��)E�b��,WB�n �G�C��o:�X�����'��٪�S*q�,��N����IF����q��@�B���=��qA�N��,uk��2U�����&�ƻFT53����M���R0b��-�8�.������a�f��].��/�x��!'�c�vZsX���3�ۡ+��Q�n��&���w�����d���G!h���(���d�u9>�Tkl�j�_�X+�by�*r�9+%�Ċ�s��p��yѠ!"׃1l���jT�W��2`鮡#�P���'IӇq��1����> �;�>��V���euŮ��F��&�X8�h�*Y�#q(<}�v�5�?�Tni�}�ؠ�����ط�@k�J?��f�^:n �1�v
��d�nS�4u���$f�{�i���3;�L����FVc6����v!��uoP-A����/� ��*:�T�cOȨ�=�cھ���ߪ�:B$ƢTB���Fںjt���$��b���F���w������L���V���ZJz�b�,��}�榸NrV��
 ��9;oI��0���Q15G���6ԾZy\��� ���F��ꗽ�<V�|Ic!�ewC�S�{�j&����}��G��;�]+N3y��̭��*�%�K������@y�[w�Q7��h Z�Us�QkM����G,��8gm�Et����2U45~��������Tad�5Z���� y�\8c���f�m��MИ�j	i���'��?H�4K~(`Ϸ�Q�%j/�w^]~��M��iG @���A����p�]�~:�&I��N��nL��������\ܑ��# AH4���!�XR�TC+�f�0p�I<},�lE�$i"ɖJ�r�i���2�jΠ�o�Uq[��0���3ÓO����|��zQɂ��(��d��TT��Ҥ@������3�3r�zA]����*s-vnDa�s���g��p����0��2��o��*c�~R.C3�l֨#��$n��	j�x�?c�m(?: ��%0g<,�݃�b�7�cz칉�_7Q�J|`����E�|l��Z[¶��n��Y�q�n��߰Ye����F_NY��߭��b�G��;�2x/و��� �U�J��kz��~��_���n���y�K�W��6,�k�Af7�Ґ���m5�Ŝ<ܥŤ+�|�Y��|�ӔJ�ר&���w���>C�g�C;�ss0~�u*� �1B�SO&�ԯ���(�\
�wR���������\��#�P?R�9�F(
ξNq�c)� gN_,����60��Mgv����GIev+#������t��Fl�19�1��6���㥌E���"<+S�s�d��(X�/I��߮hP�M��
��6[�c�dV�d������	]q�ےM�Q���� -�s�#)�r�ܦO=?��TJ:�S/��(�g?E�'��˱��J��y�Iix�\_�2%jtyb����aɛ��z&�'�����/�Z��9M���u?��~�7�_����� �Va���㟡NEO�#<T���R�/kd!�\�����D�l��%'|�Q@�����wYx~ꊹeu<B��Ι�U���j}������ԋ��K�q994�J/��*p+��s�Qdp��kc�(��/�'	���;�b��1����kh%�9���2�
�kό|��t�wPm��-ʕD���ϯ���t���ؼ�1T����"��o}�N����_/�K�O�!�=�X�����2���8�p�O~���
~�M�����AXc[�l9�b�	ɶ̭��W��%�>������e���\�S�(��A��b�O��"��<���5k�y����^j�'����x���3;�a-7��F�nU� �M�u�36��~��k�Mf�"���|�Y_�A�����#��r�P*ؕ��M���T1B')=-	p.��%˘[���>�i�����?�MکQ�{u��v+� ���qܝ�eht�37�����$�Z�T�U0Y��!�7(�Z2c���d�SVlf����R�EU:y/8o�7I��+[c�d	tգd�~�7Zq�8�n.Ҵ�������_{�BFpꢿ̝��]�%�?jO�q"�r�@���7RfK��p�3���'>9j��{�fd{b��0j���]��]!eM7μ��l=,J%�r^����SN�K �&�sb7W%��h{����kU��ކ���S*k�ϑ�a\3��\��z?Q~�Z� r���iz�/���K�����o	�'����)�,�M�J���j��
b�U���F���h�2uh���s����h[e|�j�~U�{�E�>[}ìw�F\�8z�"p�TBK�"�6c$W�I	�����I	T��Cਗ_#Y��T�3K>�^�V�R�� �7�Um95�QK�.lV�.���i��eƐo�Wg��Ɇx�{���=��� v* ���e�Ng�F�"��5h3�D�XkN�V��׻���<�ڪ�)�,<��ϕT��'��g�&h�}+˥����]�u�+ /g�^�6yT+'J))Qø�<��<�yG$7���:ȷ�g�!I =���%�\�\+�]͂UU��� �*���?��E��n�)����^��i��v�'��������X�K��*@ZF$�v���lL/���I��2oЖ�9MC�8�;�5�����2����f���y�Jfx��5�ιvxI�! `�ܦ�:��2� �diRʨ��rv�z���?nD�_�`"��T��ubJ_��цU�J���0��Y�yY4�S���I�,��4Ve�E�0w'�
��׮A�n�S:2� Q:B�d�s������̽�`-E�qΌ��,�uЖ��~�����y�&�e��5r���Ő��.M��:C�B(,`~~T���?�� ��9�PK��AU��hol�q���r��Wy�h�oR��b�dr,�U��`��{����f���5����B�ܓ����7����(���f�#�	�i*�5�m2��vV�y'v����S�F9��a������Ehbp���(�;w��#�M�GR�p�(vz�0���q\�#��qzo�qU�p+��{�D�\���A]3Z$�����:ǆ~(7ԑ9�g�0�Mp���-U=����ťCI����ӺlL�ݰr�~;�w7Q��:���C6=�.X�%9����kz��'oGA�TdQ���|������oìNu��i���#���%|0������R��Uؓrg�q{��H���%Y�
�l$̢F��۷75G����uN�T$��DkL�xj���h��N��*\�7-1u+&X@s�|��J�2�B��n�8J����z$%�X��rDO',Ȍ���6V6�EK���x-~�*�$����&����[��k�{K�W�|�J@p��衴�.�ǒ#=�*kNiz�����;��,C�B��<�m�Y��E�d��Fs]����v�h�X$Ȉݦ3{���q��Ò(��o�ĵ	Q�c2�ŵ]�>�W�$�gq�i�Qʌ��'0L�g`���8"m�(}����t��]G�H��}]f�Ų��o\P���{\9-� �i)�?�����>���*�	*�O|6�}YQ�7���|��+��_���#S"fΦa�N���Q�;׿vg�ڇH��W�S�,�AJ~�Fd�ѯqrٕ�wDN�xWp'H���	�7��-�lC������%x�y]L-�u�O��L�����EvY��ǭIk@ bZ(�����	�n�ղ࿣�("�-M�+uR��"�Aݺ2.�2M�������l��Q91��kǽ�_�x^��>�y*��z�Qج���-�дZ�Z1���R=���#��}�NQ���k��;U��ң�o�d	����O�������vM$J=���)8��!9��I>� �@�| �fZL��J����(�Se��I��y�e�t,���~��8^w�7���T�k�R�Lz� �P��b��S�L��y$�g�.�8��1���[����	�Y�O��^kf�:��R8�����u@��j���/�����}	a��
��"�<��L�����b�]a��)�VZR���<}�k�?!\��pk��ZC-paT��Z� 
��l(�~���� ���@2>��l?�gpЂt,NYE�:����?�fm��=�%.���Y\�F��&�`�
#�t �B���qWJqs���G|=�ֱ�)m1k���\������'$��Y�.�\eEX�
k�;��/�i�g$�T_.q{9�"#�����)�o �F��uWcl̼ݠ�UW��~�8�����0`ܹFSK`eI��!���V�
X���1� ��1Ȃk�!�d.��&y$�,<�>T����y��"Y`���uf��Oy/xb����D��~Gh�ނ�*4�*�CyL�V< e*UP:5�Z<�"��&�*�]	��h�Z�d����$�̘~$\�eC�d�v��p�&��Rf$��j�u�����)�L���H`%5�[��j�:��`��:<�h�D���<��E��G/�߀"�N�Ԭ?g�����?��fU�j�łm\��h��F�T�y��Wyb������P�y8�N��Eq��>zH�ҍP�t�/[� ���٧[`2�H[�071�RqR"�5kdv��Hv Y׎�	Q�ɏ͇{+	�ng6�Zp����57APn��0p���$�J`�e�+���?�'/��`!e?a��
{�R��G��Ms����
|�}Ү�m��f�J,�9�f�Mz ��჏��WR<�̴k�����a.�L)+ �lަ���̗�I�%�����Z�H�%|�<��E1���py|x�g�hv;u5O�����u�	����D1��	�����zt�����c�@���@�����	��z	��8�|�?y���ٙ���ҩ�癗x��&��rP 0���˰NJ_	bFvp=�:f�M^�[�c�-'C'
4$��G�R;׊Ķ�1,�A���U�]h�JM0�ԋ�+�94�^b�[bd������@G������&���	��P���va������>���:�9,���pa/�\d�O��$㍃�% ���8�3W����-���EBMWʜ�8������#�\Q��Л�l!<T�q{H\ۢ���@��D<�yO��C�7���JЀCS�uJ�2�>�	���I��BT���2�v��!��O�k��y�r�s�_�c31�����9�g�j��ë�Wf��G'랕W�vPkp#u�C6Rզ ~�[��B��p�H�6<��9Ӎ��s��1S�e�1�7@i�C�)���^�r.'\���q�+�X���c���?T爪�w/���ّ�A�6�Q�!�Q�t�Q{Gi���V�i�����bN�G���H�a�y�kS�Ͼ�b�Yo��/����r���$Ϥ�@s�i_��f�?v�jo�f��U�O4�<�?�{S�A��>IC�۸�k@����`�� Ǵv=��#_M��
���0e�JՑ��r�e[;c0��т��n�1���E3n�4�U��?�mt�G'�	�BJ�K���-C�c�5$q U��_QC�q/=��������� &�v���*�Tu�zk�E�C� ��V$���l�s�4��ܩ�3H��f9�U��1�W��XșlPN]�Z��������\��M
���0h�H^�Y�`�u�"�'V��s^��h����m&\��7Ȗ��-�;�����v�kA��� 1���[
g��p-�y��n��k�{_{�D3,�Kۤ6:���m�����:ΫuD0ҵ�,����o�7� "�	5őG��5�O|C�H���
V��\��Ә��3���`(��=�U;~<J &K�)BWr���%�7�A��>5��h�F9D�����(�˙b�/Ld�7'G������_O%6��|!�0�ۭ᪳�L�A�FU4�HU ����C��9QD�ÿ�BAW6B�����g��B3ؠ�v�/<�,˟�"}5}@�B����e�L��;�4p�DQ�2yeT���ҚGt5cj*�#;H�R?���7L��o�gl��lE�n��Ѡܯ��CO��2��X�5s?	iJ����7aU@[�<�ժ�tl1�z�cN��R��u��휼�}�;Zs�e����mfZ��E{�v����k�H%Ae�^H��J�3?~$lo�{F���v�Lt�<�DJE��-� l0Ӫa�J���	�g��|l���-��Cޯ��7N�l��蠍Z�3b���^R�H8��n���h��:�vz*:�y�*�C]޿��{���S��Z���=b��� �g��
2�&���� \J�&��p��e~@�����7:\*��4��b@�� �E�w��C"�ĪP�n��LWL�h*�\��x`A̲R��Obj��Oj�sX��m���T\ `~�EU��8�P���k�5"��U���&����:�еMR\��D��Z4y�Y�Z���N�b>���4	O�=r*�I��Jtٚpx(�D!R�H����C�l����d�:���]�9~\��Y<-�Eӵ�	��,R��9�����r�+vR�S��H%'oʓ����1޺��i&��&���w��_0�BGo�^1~���9�������t��oz�]y�"�ݺh��[Ol�e��l�!ky:و�-��	�2�BX)ȏ}k�jk��b"�f ���ǌQ��0�����n~� Ju����X��H�nؽ��{��-�]DY��x�{D���RG�i�Y6��F�^/8���0��B���p�g���X_uƦ��۞�kn��ŕ��f�4��A ����B��-�"m�C��Θob�8f������(d������ֺ̭���Ak�|����eiz��X�|�]Fي�t&N[�
p�%��a��eq�8���&�< @���(�3;�f�WRH,� �(�nX�~�y��l@�c(��'R��&�ߣ�Ag�c_0K#ʏ��(�p�'���¹�$6�8s�|[��{n�U�uy�JJH��1�8N�3���~�qכF��+<�U�5>�����t����D]�⤼�W'�P��{2��z'�>8s���"^�@�q�?�YDm�_m�r�/���4|�s�z_ ���7�u�^E��n�Ec��݃RϷs��{2iL|3wwnR�^HY�>ѯ�Zrd�4���>�qáC�9Y�jP���z��$
��Ѯ"{��/��h��5�E��Y�L�b��v'D˿���?�ۯC��r�V��$�p��wzt.�����OƧWj$6v���q<L�x���hK��,I��>7"�{���Yϣ�eeLI�꥙gʆ�9`I�U��������O����WʑN��ҵ ,��g�q1�Waw�ٶ���k����cK��,47Ħ�S�U/�L����������2~h���N�v�!��MZ I�V�C�<@K�@����>��@�_�> ������8J@P������m��J\IٸtU�{�׽Zr�?M��A7ϵ���.m֑�"�A���ш��`b��QC�W����t�s[?BwD����K�b�2-�����A�Z�@�ty�~qթ�=){�ya�A���O���~|60�}��mt@�'�y��]��X�����Ѝ��&��k{=R�H%a�Vxˀ�g���#�TT����|_i6�CN��'�=�{���"H��a�E��b�.ǖ���1D~p�(a���Ow!|䙨S��Ho�����N�Jۿ��CKٵ�D����f u�[7��4�j�@x�)]�O����z���=ڰ�h�����砬P����H���\ʴTo�:����}�B����IuԜ+�LT��l���d�6mZ1����os1s�;�'������xP�f��E��lH%Z�cR)�b��7����S�L]X�d^b�g�ko=��37C��L����*H�T��5���v�!Uh&�&�2���
��y�/j�&�r/u�~��	�	�v	�A>1~� �� Ԣ���5�X&�0ߵ�I��>z�ӱs�N�L��1��,0��Ǆ��e�5|��X�菭|"W�{��2LT���O��	��4�m�ޓ�wz	��D���� u4��`�|j��<�>���)�}�L7��a豩l�Y�c�ԧ{G�ψ��J�Q�O�F>��fs�"q��P�`��A��G:��6��|!=Ó��yH-PPǜ�Ka­�d~�g�g�ş?����������`��jJ�bx��"Ӄ7�9���֜���Xsw�:�%�K�\;y�`	L�^��X����_�a꒗����{}Uޤ������0��Tr�n��)��L����W1[���`�TwuaZ�K��̊�^i��JX��[������/կ��̹��H,�0Z����M�����4a��Go�O0=��]����s�
1���{�KT����Yp�{��l��$��f��9�4����|#����YA�`ɴ�t�zZ˯��Ѥt�0-��zM�I ���u/�ࣈ�Ih����ەO��)��!�9`���#��&��܄��'e���<�J ��Q�� q��g����F���{en��/~���?9��џ��������	��f;36*�bۦ�H,]���C��{�S��Ǥj���*��U�Ӷ�/H�t��5�I�{,hY�x�Rr��V�����������,�kn&��1�)�?�KFU��q"�'�͉>����X��]��$��7NK�J�#��[���QZψ0~ގ���>d�� ���%\;��YCIp��}Z���?��E�(<4���\��o9
1�KN�<mǻ:.��j�6�T�@)��SBQ)�L�'ӹ�ϓ>�����6m�%7���[$B�+�r �c��=$wv��I�vjn�8�Ò�.��<�Zǁ��B'-�J�����ܶ*��X�������4G��ă�x
��X�t���"y�J��w�[�����%9�v>w����=������+퉜�܀�u$itrol-���^xyn���˾��9���:;�*nQ���4�i�f��y:��aW�<�]�n�!��E��a�3B�����ڌh˲#����7�����L�5.����N�4�p��.S�x������oLN�3<�ݬ��v�(�R��A7A��>�򇗴���h�i�E�2QB@���c���2)���ŧC�'eӴ��ڳ�Kx,���JB�����P�rq
GݻA>+>q.%��jKsٙ]7tq�{�fQUb�z�K��`�r��M�3y	Vp�w�gG�.�Qr�7ő��w5�_{��5w{�䜬�R����0zJ��tN�(ң��5� z����IY}��Ԗ��k��y�|��LML����(~��j�~����䏗@I%�Uh���b	�U���4���b�A��ŗ�Ј�|����4S�����M�[��D���W�ِ�����ji���@���9��(X�;��G:U�f圅#�(⫥�8�i
�@P@+�䇛d�԰T��ϴ$�j1(
5-5� b�y��h��g��sp�$V�Zݘ!"P��o�xE�R.F�H��h���r�����.9�Ґ'���}*���_��Ƙ���ey�GMj�t��4 �tls	�G&���R<%��ip�Ayu�l�·x͢.����14`�'~˖��;�`F�2���J���@����b��DB)��?s8I:�Y�:q�5 Q����>����-O�U�!}�x��g�	�v��KS;l|�>z��Ը^]A�f�8�c���z}���|������Q�O���O�jl��7� ��.4��+�2�����w?���-3��7@�7<,����&ӻ�_��I��/�!�6��@�~�4�Њ:��Cn� ���`�ˉ��x�d��o���џ2&��\wݓ�K
�=��U3�_@x�%��o�x]څĀ�[~jD��&Wug�����6@N(>�G�S���?J��y�߰	��� N�܈� �~~���]�@�,�>����ɟ&ۢ�<����-�w�:�|�&��ꞛ�<��4�Tc�?<}�t3�s)7V^ܯQ�0��6�Y��!N��[���FQ���?�����8 ����RH8���`��D�B�\WߎV�9����}�
4vd{����t��L���zz�@�Ȭ�"u9QL�xaH�=����@Zb�x4Nk�c+��1��q��P`6`��X�@v%��ڟ��җ���w�!k�b�>d��.�^�P�vfU��C�7X��<W5�ɮy�S�j�J��d���3�޴�'9$��W�ck�^�j�o��#Bs�J���|�����&٣�ms̞оDo��Z��C-^�-Zz W΋8��ғoA�@�KF��NK��M>��i�a%hQE�/�������/�T�ܳ7�́g��z��y�G@���0_]�Bq�:��p�.I�(P5B1B�*^?7j�qw�o���%2�>����@�4/3i�z��?�'�P��IP+
_|ȁ}����'r��)�	���n�W�F���F�w~4������&����2J���mS�q�،�+4�Q|(�$�8��q��.-�O�� ��/5A�ed
�0�o��(*N�F��X��a�臀�_��!����4w4����~�}��$�.�6�1��u`0����YȣM\Uz�����!���}(����)�S�?#&`xX�CHn�
)���A>mE!�ڝe�Gg ��(�/Ōٙ>��	aw��"�A���5��Yh��V�n)I�Ig�_Ϣ���䝏��Uw+}A}�����{'�8�M�'�����[��0?�Q3��0p9]R&��L����!���5�OXzK�
]�si������c��5�(�����z�^:�����Fr�cu��^πS�Bܠ�s��#p�9�{*�ht^J��%S��͈ʫ����u���
y���҃�w��@��+7n��(�dߘ�v�hn��n��'�E���)_�/T�a�}��,!A�G�?�-Q�T�a�߭j�|�z6v]�X����,��Q�T�o7hȈ����h��G�|�Ȝ����	�RO�>�2{>�9��A��V��ƽ'Ǫ���5���$����Hya	Gc��2���`yqrp?�_v�ա0ܦ��A�[��-���r�9�tb��Q����'�m6��K�L��	ɷ���q��H�UV���c�<[���8����E�k0���M1��q�	��J�j;���M�7({�弫�3E�u���n���)�nνZ1�\-��n��U�3)�0mLj��Wz��ҹ3�	q��d���զ��t+���j�u�p���7>�!.U��u���)T��r�3��/��M�K��n�y�Q�y9��_f6�"j���*����T�Y>,,�ݢ�E�xz��ո�D3���u:
Ȇ�t\���{)��`q�+2���>����u.�߽�����9Q�%��KT^p����k�v����A��i*�\cZ,�)Do���$(�j�|9���ʄ����9\D�-�Q�u�łL��\�D7�2d�5s��?@n������A������cg�d�z*�C<%\���1-���у��a���cDc�~�R5Q�� ��Cqs�"[�lh��ȌER�����MR���| ��>��
�U9S�����zӸ����G��
9���!��/W�2���z��H��畨�&��戒����WTt�4�s_�l��D��|3������ 	��-)X��R�~��"�l t�B�@��=��\2,��D��V��#�Q <
�'Q-�@�Q`�=�-X�A0�)>���2��K�7��0�b�-�b���UM��~��z,������:�w�aCK�H�B�a��x�g�F�7U~��z����F┴ğ�zgeZjA�hs��X�;�c�$
�����^Ό_Mxa��8ޘ����'�g2�d�q��D �@������v��c>��oTә].�K�6��9� g�W�����%^C�Gt���Fi�wN�8!���?6G����im������Hc����;�#�&L�Y֤+9UW$蕲[�R��޸���L������SS�y�Ё��?%	%{����$6��l�E���U�"���[�<�����.P�}�^O�h�$IiR
�
f��a,�M�ܑ^�!�P������p�B�� 7�K�G=���%��[\k���h-B~�-�7��GXr�kR�(�J������l��M.	��W.��8Jk���e�D�i�t	��[��
�����#ymy]ߕ>ӱC{0�i_��F �#�S+K"!�Y�N`>���k}FV�'yH���\O�H��7�� �?���{�񲙳{y�:���u��� ?�g`���!�QM(��?Cv�j����9Ϫ������~+IL�<m��ۉ,n&��;�isQ�"������^)H���Eq��5����%�qV��6�"/sOS�������P��1?_'���C�8�s��c�4}��2"ɑdo$'���F���=��Z�.~��*SC6�YX�1^h�	��B!�݅��kE0G��:�p�>��;�Ǎt'ր�{k8�)�[���G��9�~��%|�1o����.�[��l��$�q�[h��́�ב����nJ�S��#�s1�C9��+ZT&�{[�+ı��OFv&���s��Yt8\bo�TR)�ªWai�N9�U�'!�bd�a)�n��u�4p��*��nDR��1=C��B:��ޒG����9��r�D�@�ʹ��*�7�Ǻ�,M��WQ���{8v��Tv�qDݲz@hYm�6�0�(v�J��j��Ey�P[;xV��ڡ{�<EVR�9i5��5Pt:�o��_��i狢`m�<ȈgL�H��J�$Bl|��	rm�U�QR\ʁ�����>������45��y�f:kxbt��#��V�ߗ	0Sd�V� ��SB���^���r�΅M2^�U�M����hN�<E�'#���n^x�L@��o��9e�f3�{�se|a��mv�'�m��аaB_?B?óO`�Bh?����n#�;yH�
y�6}��y>�b%�M���� ��3�4(q'�yhq�)���#�o�;�= �nCD�a\ݑ�ڍ�U:��=�֛Z���2 ��S�1��4���i�=�aܥp-���}�k��c�`B4����y�8����k��/�DR"������ч�OZ�6D�p3�%��Fx_0�2�!�s���L���^"�}���1%��T��f��}`��chֻ��!����/��֠��U�NBS�i����y@�|@ѢS���BU1�>*���	#���U�x�����]S)��G��L�IY�sȸ����;�;�~�=�c�Jk50�4��b�{9v��Щ��� ��m�,GWkFi�!v@�P�E��(���sGGBB�x����!�68�|(�F�8��6���*L��`"�X4�M��γ�M:�<��T��&�q����UX+�߃�D`"��}G�rD�n�)�^��K��"�|jw�kr5�/x�B�K"p@��7�"��g�����Ee�}[}8O�a.k��ɔj�x���	��C*���1[����huT�w��Ц �Ό��C���:E��c̰����ꪒ�e����C+lB}M�p|
�S�(j�R���r�o����µ�&�kD�x�7-�͗����qOz�쁎���kim�G�^uչ}�+�9�0��[����(!5ZAW+�pSm�21q�5\�N0��NR�~�+1b�o�t��Ow:��%��Dl�e��^�J�ɜnŚ�|,��r����P@�ڙ�V�Y��ML~��QE��^V��b��%��B�n���etn�!�U��g��`��0�Yhq_n��[CY�Y�Wy.s�!)i��E�M��i����䬙T�O$a4�$���Q5��x���-7>	�� E��d֨��p�_��[��xК������$�"@2Cm-�ܰ��J�'_$��e�$�{�Q�h�*�TY�/�KQBr�!��@�\�cǴ�ʹ�;���lb����s8z�y�9��1��Li���1Ѿke�z4�F U�o0sji�I����/�!�����'��ݝ���r	���|����~!�si����7ͅ��V��R@� �Fu���^�.\�FX����;��4��\�o뷥#m���L;f1i��nIa����5��ҭ<ABW|�����$�k9��6o��ќP���5�kq���MB��[[&Q�˦P�y�#��?��A�޶2t�&����	���$Խ6Kn���������P23.B�r^D�J o���ɸ�2{��U
#ˬ�����:N.�'���)-K����hP���Ńߪޠ�j�1���h��6v��� �^dɆ�{��Y(D����}�z�ӫ��_Y9�"$��dC~)�L�^3x~�2�|ߣI@'��P2 22ˋ/v+�T�:Xq��N�W�G6�%r��e�n�����*�x�"<	2��o.��4��,����LI�*Õ����cT�@���0KNV�B/a���ª9�#�P��ɴX}W���wP�V���s)5�Hn�׉��y��Φ��Y$�ҋ�:�Oy3���}d�$�kJ��攪׻n��2��
(K���`&�}ZFά����-��FT��b���A�D3�J8����z�>԰��Z�]�53�_�]in]D�i[�*�K�ޔ���kB?|��c_�d�B�@k�s	�m_E�L}&������+7��#�*��@�Z�8j�^�@<L���2��X����(m}/��xLZ���v��L���� ��f�v�@1��]�<-��X}���-A@�B�в�;�M,��ţٻ0e��A˜ �dH���[S�g�J��Vݧt7���2�V��>	�dI7V��ߍ\VWkD�TU��$�֭�\������*}
3��9/R�� qд����θ�1�o�|��oK5fH%��>�Pܒ�C�=���*9��Gsi�xX�D�6W�'���ƙ��n��m�ȳ��(�ulۏ-#�u�j�����߉��%�%�>a;��ĭ��yY>x�i.�1nFK�ӎkOT�kT��wSz��<�d;��p!} HX�X��u*��%�!�X�� :����Z��`�B��I5Y��6l����;��!'rO_\��(}��(�lWц�j�$���zKj��zb�I ҏ1���'�m���sLF���T$%�_�Q�Ű�����V�ȓ��|���9OJ(�����E��h�o��Kf�]U{�9c��%�s�� ,c�>�3��˦Q$U�؃5_�6� ;[?�e>��-CF֣v��<��U��_11�#\��R��>S��U�mD`n��o�hzW/ĥ1B�ĉ�r�Š��z�� �r�����C%����S���t�ot�>b��,ߔ ���ꅋ玮o����O�X@
���AO�*5��!��rC@P��Hb�w�VN��*�r�ۜ��}���Z셛B��n������[C�	��Zg�J"���z#�K�?��<N��˓��朵�ף���X�=n�Ӈ�1����CHЋ���F/��\�3t��0�=���đL����.6�rx��n(Pt������r|c�*��8�]��I(�lF]�;ƶ1��B����d=�ls�2�XndL�P��-
gi��4�lo�}/Á��W����A\�����)Nq�����/��8p�eb��;<#Uת��)��'r��'����,�C���(Qŝ<�t�W	k��D��h�H���e��1c������j/�tM����4j��-=�n�t�NvtŬc���Ӵ�gW�Wm��@9�;�1��i���*e���R�*}��왁$y	y
�.|l�P��L���`����,�Z8�z��`bb�|ʉq�����{*o"`��*��'3il?x���$�~#=y��J����	?�t�i.4���W�-[�: 3H;K>7Y�-ٷ�~����*4z�lBT�\vH!�0��J*���Pp�"��l�ݶ7=o�������rpBX�i�P����|sa��3˲Fi	�kkf��f�0�5���v+Nz��l}�MI7�5�~4�Y�<^qR�!2I����`�~õ;N�g�FI�Y��odo�r��2���0<gtj���fC�ʌ��
@(0ֻ�� X��l>]1��)
�[��C6��]r��@مӰs�����������������Qv	�-u���Q�g�V؜��ǒ]��r�"�V�I%w��9N�}�i�Up�#�Q/��eaI����` t�Y�y��Iשr&�r��g۱S�7HϞ7��p��vE�;/ma_Hw&WX,���u��@Ǣ�}�U�<�R�4���}���h��}e�6�?N�?}]%V\ ��3��������S
Y/������_6+���Ʌf�~Qr����R���̣���\z�aL������Z5�K�0 ��� ���*M@u�g��#�m[��}*n�'�vԛ�nfz��r����B|U��wuBQ��m/�a�Gw���uJ�sK���y'&`�̞cO���o�{��%i':�ƭ��� �F��U�%ǹl5t_vǯ�0<�����Ğ�����3��LČ�`�w5֭���JV����L�3*� �RY1"�C5� �}A�����,g�w�j��?S��FӋ�5".3���=���]!DSg>t`�YnL^�{L͞�A������t̋2�cW;n5�GQ�i����Z��ί��wx������ř�D���3ԛ�]�O�0�I�u00�l�L��t��+@WC̤hJ���m�Q�6��:lkt��ђ�@�X��&4cS��o�$���t���sn��(e��CkqSJP�9�%�d�K�H�"�;�~��A͵��@�u��4hm\���f�t�8�E@d
�\ ��,������W�Š���v�{6;H��P�!���d�p�ae��C>�S(��k�����uo�mCpO����k�0�a���I(�&n�]�	����Ih��U���\��� 8��l�e����G���2�0V��,�r�w�	��0���QX��EF/�?�\6�zГP�*8���CD����jlAQ��`�6�2���^m��[&l�%�)��
��]�֌eoT]226�[O��d(������m��l�nD�';ԀP��;�\2t.�M���%���T>"���f�m2�KQ���-#��q�<���g��TOuuj��B�.;Q|$I /P��ï�yf7!jq���0z����ҧ�T���+#����V" ��EA#����d��vO���x�	�(�����e�V��u#�����w�NZ%�����m�ef���`�G�~���A	��1ͭ��[Z������Y�x;ћG=�,�5��Y�~~?�/&�w�����R��65������4?�?��J5I�)Y|�:��P-�D���po��� �n��m�U�<F26�^aLw�����t��zo�a������K��k�������ۯ��8LBqI� �S���.i������h	���yd[D.Xɖ�Xc�g��Q�6�OR;�WzJ�c��ki�vK����Z�T];kd����-�G�UC�ķ��D�[�>�Z"^���F�,X���~K�\+��}Z��$���C_��W��t���vL��;|K��ҝ��5މ'n3v ��=B%�6�E�	�e�p4�u=y�6e���J�u�{�`��W��PF�L�6�rC��R�1Dd;�]��3uSL�k����@���\8l�\<,�?b�0]�g�e��r�"k�$썄���3\���UYg?xڼpG(NAH]�U��=q~}���$V)�.{s��i����j6��t݃Rb�o���5�Qj��M�Vy�,��}e.0Z�?ۖ��[������d��\br9���n,�V����}O��O6hbī���h�V�.��q'���{�
u��k����n{�-����R�2#*��~=�n��l�����ϛ(:
Rә��1S��EZ:4R��W�'�5�
��;�T���>��ߥ!��M:�kg�G� ��A3c� [Tn�ߨ@���{J�-.j�a��̻�����	���°w!�^'���/��>.���6x�2�AN��t�$|f�S�����f���z��H���z��5���Ȟ��Od��nM�mN/�]���[�A��d����0��z�>$�Y#�D�n�Ɨ<�h�CKFu���ojvZ$[�� %��{���Y���(Ta���������߁����S�K[+�v+��4���҉!���l_(-����Q�C���xoʁ��<y�j8������=��Ț�>���3or9f���Q�phA+�Q)��GA���l���G�2ղ���?I�Ve��)(���a �)��b�D��D�.�?���D����w$i���Ž�<�"N�:��bY@�����b�����Y���2W	��ߴVHE�my���1��Yޱ��.�������GuI#�[<��W���
-;Ue���QS�.�����z8��4ܬ�G�1�WQd��Q�n���] S6U����D����)���y�\��	}}s|=����K${���N|C��\M<ꩆr���_�E}��}Yĝ�f8�,A��"A�Ux=f��ޝ�9ϽFc�Ǡ�5z��d}�ԯ�hn:� f�C*�!?�ը�UqrJ��!rf�b�?�C8���$1����&J���3.�&x�2�;�
0n��W{*��s�����%z���}��s^��c
��T�����[_����b�BP���q�}�+���͉X����sk�L3�P������Q��bᆧ�z�Kck��H�[	�=}��VBf��S�{�-�ї:���4�0'#^߾z�xkt��<�����JR+�=��u9������.�pEa��T;iW��/�h:��ye��տ�}	ԡ7c�S��I��!E�r�!��7��(���DͰ�g�06לƺ*���W�b q[QE������T�`�n1Uh�o�3��T��D�T�,�N�EC��C5i����J�Z�D��Wl�����Z���Ǡph����X�cZ�%#����[�h�u��P����
H1�'�n"�4D.�˥��n+���0y:���t�-���������^P��J�4�	��9��mA��1*�
m�\&�9�u<��	V󅦔��!�үN�+�2
`���vx�����GD\�\W-C%@��J�Kwbߕ����p"m��&��`�h�<��Xi?�cR��r�yl	� �~{��Z�L$5��X��_T@�S���3�$aj�NVTO%e����sg]����~V�Z8����:x|�d�5u�t��Vc��5��*�w����b��+��k�^b�sȪ�' 2�L�K� � J�s���e'c��ɭ ����.ڣ-<(nk�)��R��c<?��qJ��X/꓆�%Z(R�-=��<$` ��F�1Z����[X?7ք�g׶?zΡ���8o�&�!���M a�
xzԱ}�
5Vقek�.h_�������Z�kC_sN�S��:�HO�e[�h9�e�.E`!ȇ̝\���X��3�a�-�-2C`��F�t��k6%Nf+�ן�I��3cX���D��>;9����%M��f��(�/uR�����AA)J��q9����^*�
OԱpOjH:�˶nUW'�J<4��n+oR1��̶������C��� ��=K}"��f�����;U��>��6X��Zj��I�A�����c&�܉Y|����|j���-�"$^ʃ��^��р�z�\��jKsH�ptZ�Ck�S^xW�q6bn��WL|P~��@�����j�gY;�s�*�~���n��g|	m2�(Wۅ����Ua��ٌ�km4���iHMGԹ���A�M1��*��ڕ��lj7�\��#�6eܝX��0�҉.�~-�r�=��53J�S�izB�axL�z�a���P���հ���~�0xZ��7�l��)��W��%�Q'}�2hu��p-z���<�\�G�_�X](�8��s�o͓�*��P^O�o�;���PCS�@���B.���c�(�B~.�W�ԉN8���S~u8�[V,��*�nH+w�d�����u�H?�5@yJ>*GyI[֑!��ݢ��7��;�����Ԝ���m�je�|(�5����e���:�K΃^�,�&��e�K�����7Tl@����(r=�_H���X�@�^��p]Յ����q1������ޘ��*��Um>�)�[Q�./\UI�_�(�k�hZA��r�K��k�{�S[h������B�0�yI�P�ܭ��sK�a�Ǥ�uM�ᥜ[-o)h�&�����(X���Y=1��9���+8�pR5�o��S@=1�_�2�weM�٢�W��j�蕮.��<`�)��s�-M���_���ov@+�T(���|?��Il��K��fs������
j��g��!�U{]`���5:��	�~���	�5ΠaM����и�D瓮����0��� ;�nA �p�����z�2"s��V�S5��ը08c�u2�Kl�t�74�Nx[�̏�ux�^s	Q^����?m�rcdPS����I6��1�>�R)|�J�c�+FT��@�zzz�����k��QWM�z�4�Y��Ľ���d��dS�g�K����ܸ�^�li,�Η�?��]_�B=s���z��FE �tz�G�;=�+O�8��Lc�9�ČzPغ���h�깓��,����9�!0�I�_���T���t9��/���0Z )��˽o��6�Yϑ��v�At�2?��㝐ο�����a�F����=��rP$�A�b�j�%�I��9�o����	�V֭���{&r0�a7ٝ�W��}}���c��!��e��P�\��m +R`8-�	�)' �����q���F�o�X��9"����s�<y��0�5�Zy,��Co���+�xmO7=!V�!B8ֈ�6}�����e�g��Ԡ*����=��Am`ɘݻ]�Ǚ{A�c�
|gj�?���7=�o��^�;~+?}���x2 /� :�
�.?�հ�(P6$�;��n17�krd��O�57ދBQ��v�������20�( �7���g�߸a��m�m�qe��	���HL���]%��E[�
%�ܾM^��cLt�	ϟ�ܱ���
J� A�5��f�K��/��ub>&��˅`�f��:��h[�=뷏�Jc��Ee<hl����o���Y�<���ߛ�՞� _S��FS���I�Iq_��W�s�ّ�e^ۆ�qVE�͞�M*\<r��@b�v��LI5����HǢ�$%�usb\�Q�����o~�x�Mms�$���~��U�x%���|��*�4��Z�<����v���?\��7b�֡�y�|�f@����X�����l�8��������$���s��m ��-�ڱڻw5k`/m��7�$?�"�*)��P�M���`��9n2x���Z�8L�U�>�����8C��]����z�٢A9j�f$��wf21���E�%d��w��s�'a�PVL	�F�@�'E��@ܟܰ!j�=tRZ!c�5�c*���8���(`�cvB/q��00��0�H���;��#-Վ�R�t�1��l�L��C�u���|����X�Ԙցsx���q<�d����ˌ�)J'�V�Wq���Q���:���s��riH�Y�
Y�̙��Nr���n�p�a�?e\U1�ː8ׇ\Ioz�/�++ܩ߬���M�e9b�@���%d¬I�jʇ��F�;��&���x�6zmw��)�+�q��)V�VoK�g��f������^�3��W*�Msq��BO���ab{M!C�Tj��-�
�M�|[�<��.�H{�[N����gMQ�o`�\q 2k_�F1��b���{m���ī�d��ɇ#O��p�t<�t��Ѱ��� }�f/�r̟m�V���X'�P̫���H�U��=�B6Y*��Ms>y�$��S�D��1m��O;�F��Ǡe*D#��T$�Vۤ�q�aRP�ڎ<���S��������C_؄��޵2a�˺F6���<�\���D���r�q�(J��K�Uf3����t���[ё����K4�6$��:�(1��醝�8�~K�F(~��fX�.S��B���*�m�)��x��aW����d�\����˩&��#�⻗�L[�˿-i���0�L��,����a��e������`M�o5O���&��m�)���+�Q_����.L)%��;������O>TM�ʂ`xl�+�~�-,9��F��S5la�#��m��0%�&I�����:5���("�n�'��ۍ,���������/��8�"yu�����֜��N�ߏ���G�q�P��''r�����GJ���s�-���D���e��gU0gi��2�t�jٰh��!$�1z=:�D�`z׌9�5FYQ���Tk3pD�� fU��Ul��aֶ��h5p���l�?���^�p��n�\�Kh�K��GS�^v����B��$��|,���A*.L�l`�s?�tf�|��J�R��D����{>b �ub�H<����A��_�f7����L'������T�$�#{	5��
K��%��e@��+�w}�����\�_rvO���l�u*�Ȕ)T?�v���D�|=y.�i�uTLɘ�)��J�L�5�o�TX(+��z��bC�PދҖ-��m���L�R>����.IJ�E��y.����n�����VT�?�!8�ךP���׺���*5�~��8���jI�;���#jY��Zd����K�oBZ�X����~�|Zo���F�#0��l��H��'1g
м���Z��w^�.�/�T�t��UD#$%1Z��B?��P�7>m��T� }Z�0ɞ�#���2q�*�>>^E�kր�Z�m�m�QJ6^5����X�&��ys�XE3�܇��N4�ED��nѫo����!v^Lڣ8^�%tV�l�H��$3��n���'*�07�d|p��H;�$���o��\��:5���~��rG.%4�i��\/3�.������/�0�����ϸY��$Eh\mҹ�KC&�@mu0h�r?��8��Av�+���8S@2E��#�1)���šG�����e��G^!��bc����bǿY:5�k�d8&~��\LE܁��̌��)'M���K����X�rX���۔�NgL�oWY_�ߵd�|�8[k��R|���rĒNM�d���F!���ia���J��J������Z����r`��*r��#-13�V�y_����>�VE���V	+��V���:q�l,�~C�"<sU1xV` 7��xQ�1�ދ'��E1�͔�/]�^�Ҥ����Xbp���PX�F�x�&��hM��iA���!�O)��Wb%j	������o�h�xe�#E"�h�tYY�ӜՐ������9�~B��0g��Xx��Z_��#!�jȶ�Tpܫ@�w�+�>�BO9�r���?o|�������ꁞ����C���)�ޡ
Q�����(`f���~�+0�1�TI��·��rL�N͢ԅ9e�dw&F_�fv��pօ�8�2�Q�C��)eqg?ա쿦�a+��_{@k3@	�c�,�=U��?}�*^��oo�f�f=4w�!�v��>���5����=����(5���d��8�.q�m@�Z������5�s�]�,뒰wP�hݘ��D}PV�X�؊/$�S;��A^k`�/�� ��9�iن� _耢��/��0���������$��}L��"g�����1��I�~��5�]cN�}�Fś��H��1Џ�*/���6ʬV�� ��:Ms�>@H�e5�+�D&C���H��� �u��0�/�����Ѳ=xC2]S:����~�=�d!�C�W ~ju�z)���Q�7A��B���q��Q��Wx��o&��Wp�� &��+n?Ez�9����������V=
�Cx�B6���L�l��126�<&D�=�: �OW@�u�sLu1���k�=|�1'�ˊj�C�F�kQ��<���;�=��� ������GlM5�Ofn��w6�xw�b��"\���\\�������~31�<H1���I$� {�s7jꤓ,�ӗ�6Z�r�*�c�(&��UrLh�D ���Dբ���5�_��,V6k�1���#�W�Է�qEg#Ԫ���AA�d��������H� �3�V���� ���P�L,�jz��J5��"2�:�K�5=T�<�G��re�:�����߭����� df0c�x���@& �޼I���j��nYYj�#c�ƥYcR}��g.�p5���GTG�9�����/�~�.�(��5� P�h�����Hy�څv�q�	VfbV/5�f�C����#���~�'Z+� �J5�Y�~��u�\���&��2��A����.�ʹo��QƆ&�	�M��~�,i��B��O��{P�Hj��1t¦��-0�P3�v��s��mY���S�,���L�2�қ=v�9�Y�O)*FS �j�n���e����^v�i����a�<dFC�[r2B�c^a[zz'P)���N]�g�6�$?�G|q/�9�F:[� ���۷��7=������G*R�2�J����?O���������6� �}2qPq2��&/<%>�k6�%_u��22[0ֺ��F�Ml?���g�9�&�?�iY�j��v����f2�N���$u��P��h�כV���\��L��ah�Ǌ������
`*���m�ݡ}�'{�Iyf� pe=<�Ԛ2���!n���	������<�"�C�M����⋍<,��D��P�
T�C���˲x(�n�.=��3F�Jg�:F��ɤ�?E1���'+nT�䢇�L�s�eV�l����.�Lb�O�8#-n�MZ�-	�eM[�\���4G���l��&�!^h�^��tQ&�{<^R���_��i:�G�ؼl	e'gkX�^��A@q�?zq+J[�^��1��!���!,���!�cKI�Ƞn��ZĈ�c4e�-��F��p��i$�|�����1�+�uA���q���e�zK��Rh� �r
���2i�H9���e1a�^��NT�*�L�����D�2U�'	)�_?�i'X�	OP}q*ˉ��ը��e3֫��z~(�����,�}{�͔�|
�]�ے>��Emq���7��h���sH��.l%b���������������_�09�jAԭ��b"��<(���J��G+�� �#�۬e�z�������m~�1��&T�z���ڮgc���Hk�}���P�� G�6�\�7�J�(�k*���s3�������D�Thy� To������ ��ݤ];��+��X;!��~�X�]�h���:7ٌ��~(}�3jO���yM?�.޼�QUU	"l��wc��!LU9�CI��r8m*|�,JA|��
.K��C�$�Պ$��AR,VK�l�C5�Xd� Zꡂ��Ԣ�d���S�L�~��>��p�r �;�!�82n�e$�*j�!c�6�2r.b~z��?!��S����v�\��!�s�j(c˱ܲ!\7��p?��A"���Q�[^ �:���\���,�|�Q�OL�8t��=Bp~�U�<mh�$�=�+g>h�Y�J� �kD�#-�
=��I
wP�z)9�r��{K�b��hvns���S��o�;��hz���}A�U}�����<S&�K�7 �(���ҏ�O�¿� ��h������_���5iI��֌���W�>��9󀄒}	��Zú����˲LN�%r�����;%u�{��$��;���e���=�P�T��{�%��5B�����sD���*�h�΁�7Mh���Lr�neyo��=��%��K��+o
��T?�r�ڱ9��K�h/��aճN�p�y�"�p|��"jZ�[k����{��:�(���79��x� 9�=��
���9��Q��1s=��`�F��R��~ϳ7��,����d�pYl�}K��E�l~�q��P�3��	P�ٓ�6��,ܷI��Z@�s9��������⭊�m-q��S�oa{m{������'p�^[��VO�~9�2<�Ӳ�٤\>��߲>ԑ�[��RF�����������;��9�XH/��a�C�h)8�򻬪��$L�t���H���قg(Q��A$]�F����'
��l�[��\�'Z%~I�ҵ�"��[3��G�Do.�:8Wi���8��R���=q�b8s���}�th�a���!�p�Z���w����t�$�Ђ,ÛNr�W�BQ�;�L��?�b5�`ҝ�"
���{���EC��q�8�3���	� ��GuGᎢ���y�y@d���]���_L�=�//q�Y��{�K?Y�w�B
	y�*�4`�ِɈ��������@���z��dƪBV����j�u��k����V4TM�

y���#T���ݡS�{]-�En�vh��%l�����z�!QJ_�°��"�J��B�՝�"54T[Ud���;ɍ��HW ��~�q�n��]8��"�-���~� �G��:2����`-o�f���užv�M��|g��-�E�ӊ�dbuެM�1H3��eH��: ���=x�H��**��)ہi_ X.�p
�W���R��*k�'n�Q^�NM�K5&��C�U%�p����\wK�T�l�pp�q�S���7�{�Ήuclw '�'cp��IE�ڤ�gHʟ���"R�F�Y��=�����r���}&f����)y@��Y{&�ı�M�9��(���]�1���<�\Z�R[G4ל5�ѫC�H��L6��u����vL�����j���n��J������s[7)��`���T}�n=E���Mvn��̙���d\e��{�
QgG�ϖy�����~M+�V���w����V<�_�B�MI�϶ӎ�+�b��|�U�BF�̖|������8{�\f�Lt*r��4��D�����cgY(��ڭ��+�N�92Ok��y�u%��ԏG?�~rT�i�3|C?�K8��A��ޠ t
PC���Լ#gڼ��6�Z�3��qe(�}{0��@�Ye��U?���j3��fF������������x4�6�����z��-�΀g���Ze��� \���)H/��mQ;|�/(�3�`�OU�K�����I*�.�R,7������\E��u=?Q�H㚃�2��)�]�E[�u��LA�f|Ҫ�'<�) nB�ɏƀ�J�.Z�����s>�����auzFZ��	�+�C�P9��7�L8�5K<=B���|&�Z� �`,6�U�dr����PYJ��!������3K�E���]�:�@�
b!�w��4�;?37��28Fq��"��s ��������(k��mX9��\Z�����^��ĄZ��s���I)�?�;Kf6Ť_5 ��p%|d�}~�_:��^�R4�O�L�!�Ox�����j\Q�{���_Yp�w_��ot����K0�S��^�w�?��./����*Z�q���+ �gÇ�M	-�X-�/�{��n,��R]w1{��ֶ��Bx-?�_塊�g	؋1	��VYE��0㺑�!�CL.��i��!Osy"=������f���s�؏� �:��5)�{�+��3���Η�>f�.+�|p��wm:I�I�n�Tֻ�1^�M��%�]́#ܝ/���.?p%t����!� 6Z/�T
����0�ZI�A"6
i.�H+���"-�YH���@��}
��ʂcS>�^���9�3�^W�pL��ч�Çk�<�$@jmiw�ҲS���:�`����zN��	?KE����:(?OLL��4�쮈v]-�#���1x f͒M���e�;<`�Ve�&�<יTA�a�&��./��$:g<b�]	��.;}�w���i�'�L�&�����Vn-T~j�~D�>w烢�|B�~Tw�u�s�M5-���"PĮ�Q���Y�����2	"&�+�B�B�K6�?kQݺ����������wCi�y��e�RO0nk_��>�>]/�j��#h3���9"^Cx T��z����;Ś�\e����R�+�KȚ��s����a �����5}�®��Z�
���}��]�Jl�MlH�8���4���jYK�L*{"΁s����"p6�9~>�?�)�E�֢m�ը;߭^��)'�ڏ���5������m�dIo�I��?�����8r�7x��xU�i�Mb�y�BŌT��"T�j�f+�_Gm霪Ihl�uQ����:$�J�@�0ʀ�y�:��.F����-�hՉ����AG�7�K�8�Ϯ�l��*N�$���i���)�
��%W<Yq#"��]�}��"X7�%6���ʟ�+�Ɇ?޹�L	��I�]2Zc6iO�8Oy�����."��h��B��L`;�t(/(��-�l�Z��a���`��4qDW��m���$YR݊���	��f�Z=\dA�L*�([^��S{U:�Ո�ѳ�6?ի���0x�	����� �oX:�"^�ZSA����4�c���=zF���c�d�)����3h�ڌl��A��㈢��䦘4�+��@�$��O~�6�U��>(yCMֳ������~��_��hfj�����Z ��%3`�/�\;���u��d3�-�ӏ��c�$�M�!?f~�α^�T���� ���?}���\�em����������l��~m���R�?�q��HM���螷�X�dCd��fӢ,��x0�~�7�<g�\T������_U�X7u#d���Zy��kU��U�ﴵ�9����*ɹ�B_�o���9Oi�Z�[���X�Xz�?]tq��H; ��ciy�����2�2�S�=cy��_��G�M��N[WS�c�^�Q!�vx��K���C}�8��fg1���F�a����^�E?O��=��q L��R�P
�6S$gy�1�[g�vl�,'D�.���o��G�-�ZDJ#��o����N��]v��jG|��f��_Z�CXRWDB-�{:� {���CwX��d����AI�}!���nF����(UT�E\�5\{z)���5���2�-�!T0�� ����]�Js/�B�e󖵵�~A!)�KB��_���	��뾄���i�wm�Ty���# 8?�u�ם��<
으�l.xj1gj�l(���
���l�l�P�ȴ�<��P�;߄bFK�� N��/���+)����5*�
Q�AEs�5��׫�E��v��V��A�mq�͚�j�ڞ#
O�'R����o&od�@>0��P\x	$�Q���~�B�����~��Q���!� ��Q��#E?��R���]&�W�L����	��(�_>m���fa��5���w����E?��������U�#K�ӗ,����A�|Rɶ���S2!�g�hE����Mc���@|�#��<m���L�_3�郡�z����J���ֹ�y�U���zV�.��G\9���_ø��μc�hy����`,�d1_�3�s��~��S�,�X_��0x��㖧dfi��B��Ae�HT&u)0TW~�j�u=Ώ@&�ڏ�2W���A]A�����Cq.�r���A Ruw��e_Np�i����g�SS��:��(��ͽr���?C`�rcE(	�֚��)av��&��V7E� �
���}PNIѿVsYr��z丑?!��
��&��l�-X�����]�O��M,��d6	Ѭ���ԉQ��$�� �u�-�Y7홢+|�T~s���1ϚW2����%พ� J��ϡ�v�PO��+�Z�|R��u�kJ致����7����2Ӏ<��3M�?
��$�LN*k��.	�����`���~�v�o�<s��������C���1��,
$P�������t������!���X4f�����VL{�ӽ�����&����89��p�[u ���z������9ݡ�������ǡ��}��y�#,��Kf+"�*��`��"5x �{��S��X���L/�Yľ��s,2���r��1�rD֍;�i��E�����[��u8���#2�$J���6Oqpr��K{�"��ܻ^�sز���g���Cvyt�>�1W��o�n*�I�c�B�AT��c/��!&"�� 	�f!������q��6�d�٠�����!#bm���p��I;���0pPN��CM��n�H^.^���Y!'� 8:����%��>�G�鶢3 ���3ׅ�L0�S�/x��D�Q�}�k���)aċ6�9�K��Y��x8�T-㹲B'��\���t~�ff{;&)�f?}n[�7�y�S&
�p�l�nl����J��*���`�~[{��&�򀹅��oc�Z���W�9)X����Ҝ&XPx�|�s��[�.�H��N<J36.���Z����Eb�FE��L�JI��LP�y�67,YZ��/d}4��sO�$��(5=�j $%��%�?��13@8�%m���uoE�@.�Oy;�l�-W���Q��(�7;k������e�7�̞
w�rː]h?�+��0��Y� ��:E9�K�1�}fIF���)h�KCWb5_�?s8����|����^^�Q-�8�G�9O~e�|��]|�d���i)�����T}uaPv�\J�u��ϯSl}r�!Q-����$�V��3(��E��Ab&*�@)`�?�M��=��ՠI��{M��Ξ��a���r�J|�K�TM�y/,|�|�y�hs�$D���������6�"��]X;��ZhX�n��C��8���ց�N~�1�A5Eo&<v��|�������D�ٷ�љ��,W[A2*��؃~Te�łua��p�~�XT\5�Gִs<�%�>�T5w�.=9GqB��n���?x�x��Gbb�.
�����u��霅��6�ioDP#wR� m�i�b�w���㸴�fb�;���i��o��6�҂��ұ �%��>�Hv<�䟆�|2�c}o�LB,5��2`g��B/�i���Ҳf�����{Z~-3�U51�|�0A{j�O�և1)y�e�j��ӎ��E������y�Y�?^ȇ��9j�Ц#�K�ƍ��H�ɻB� '���b��)�r��q"�8��_?(�k�/p�h��+#9�Jǔ�[��Wb���q�G�ߞ���uw!]�Ae�{b)1|X�	�d[���ۼ-��F��Γ��$�n�VLE��Yl�>j}�%�~)&d"� ���@J��{�Ƽ"��Zn�A�<�b'_���%���)N�>�ͽe��(�(�r��Պ%h��9��Q���&��MM��-3a>!}���4�cx)R*�|�:i�,f{��Dhr����ƨ�jlX��ghܚ�gD��|�n� Жꥨi�6H�뚺G&�r\4�3L�mɹCUE���}V�)���Ȯ��$�d#��t}��r�y�D��ƞ�L����s�����Q2�9�${�g���Y��Rz�/Z�2�1�$����t�+��S����tr��� =�Ό��GH�s]�����Z��<�S>�dP�����7��y<}@�_��Z�-�"��va�F�-��st����PN�ZI��}���߇1�����Ac�P������h�y����%�cnG���"��S�y!�:�y��UĎ+@���~��T4�磋 %��g[k�-:8!l�ӧٖR ���eP�ΜUd-)��L9�fq��A[�x����cjw����Ĭ�DV8ލ�9\�O,-�x.9����="�j��'Eg���aB�y��Y595D���^l\�l��޵3��v�'�p:�
^ k>�����i��Jo�u�Ӥm��v4�*b�ȗPV��.�~gf�����|j$rl����/L����0`�ζ<��
��9���U�-�����6���&D3c�cD����ģZ����wa
ON%���r9�=�Ĳk�4�n���(<N���Q��tCBE#�L�Zhg��������e^�X��%h��o}��o8����D�|�H,�t�E[�m�A�����C�)�*B6A ��#�W�/�@���B�y�0ǣ9��5vP�� c~��:�R�&����"�R&������I���2]��Dʱ�F��E��?͸���ׅ�_�~����Lyk���%��)D�M��\X]����3��!h���Bؔ��������$�a}ND)�R�Vc�qJ��k�����W�Hϖ>�����F��k�V���}҃��i 7���@2��@8�lC��d��d�f=���n@�2� �{�YS�}SW�,\A�n��4r.�v�����^k�̈́�E5�����T�2�a�X?���KpuҮ }P����d-1\���k&��r|[-	����8Z�mO���5��Y�£l��^<nk�e����-����[H�;��V������(kX�]*�� ����b�	���A��"�_���#�zb������Lp�U;ӛ?��0�`߆By���%p��V���-g�)Rە;Y`Gě:��k��&l�EC ��z��
�4�eV�A.���ˌ|�~��3���w���_�Z�1�i��;ݓֈ���֨[���s��֗S����K�1r��8��麦+��*[43nL����<����g����i?T�|DR2�ف�8��؆W+�?ܜ�����ZP�t�l�ꟄDL��k������K�t5��s��nd;�r����ɵ,_�&�y������D��_�����:���#
1ըJ�Hg�]���-���H��s��_�~�N �Ms�N�`4)�nu��)�] ��o�K\����`�9n?�����/6{J�?�.��W�@�Hp�_Y1�)�M�c��z����������ƺT|����<`�rpe�0*'�a��l�eU8�'p� 07=U0��b� ��-������JA+� F�K��;ڳ�dV��@dx�.#��Z�@��,�?�܅_DT�b�#m�7GMZ���Tj�6�_0gQAZ��)E�C�Y�ޘ����g��^����|d���{ �%�����]8^�����9��L�쯚lS��f�zS�v
ڦuE����"�ה�3���@��L���'8�0u��Y��a[*V4���D'_ƭ���������	rR5�<\�њ�L%o�`��_��ռ�\�Dr���yʤMI;�<
��u-L�H����!���t��@����/���"��v�#���+v� V�*����˰�i�f���l4�/І�<uTG�`�O«/IDRyY��D��'��	�^�]~�.�pl�խ�3������+�%OF0��ؠn	���%>B����`w�w0M�r�I���m� �nX  ȭ$db���O��9���V����5�1m��i���H�	�[�*��'d�O��6��p�Og���N=����$;�)W9�D�Õ,�Kd)��)�Fi����4΍��WJP���4�-��tLI�2����Z��������l��,�d�ؽ��ЪϨ���dGw��a���aY������(�����f��5�d����S��k4���R�	ے��j嗐�a����1��}��m'�N���1�7��Nzmrr�ܥ��_&���7q�O!S���42���p��ևvɯ�c�˶�*Èk��-�|���ɢq�pu�kpx釠?"+-?���L6N���j��Y��2�[ �<��n�.���t��m~0lN@h��B�z���:݃�e�X����8]M�p��8O���������z��\�����x�{��h���<G���s��3�PkY[u|�"!�3�H��+D`��M	��
l��P5˴ߜ��!t��T���"M��mE��Ϥ��v#�	�RȖL*mq���,�5�	�1����8�'?�evs׵��>��O6Uv�ղ|�2~y����f�7�@���8
�z(B=��Ǧ2.{ˀ�a%e��h�\Q��h�9��1���~��'�V��뢁��2
Oʇ��Җ�P�)qߝ�̰^s�kIP�D�31`@�P�m�^)NG!�prMw��ס}��WZe�N��
EF�>&ٮiA���\5U�v���w���LNߠ��Ct�׿m{_�S
��a$ۀ܂�R��'��坕�{�6�����a����/9�[N��� D�W���Ԇ���0�bt=��^A0��k_Rr��a��E��HlT�N�@NA~?��2�̖C�h�ǿ����FH�[�tD���u���ZU;���U�:Ky���?��P"M�)��X�اؠ�{���+u����{U�}�}�X�׊�ބwG�ʌ�m�Q�z����>w�T��T�%#{_�8�"+�M�W�F��b�a�9U�/��.�3��/o��]ѓUY0�x$W�m�l�jpK�f����h�J���,�t�\Ȑ�L�&�Ƃ�D�Hw�>�o`/�E��VE��iq2��d�eꭇ8R�)Z�d�����qjOR�
	�ɻzN^/"9y��݃�'Ʊ|�zy�|�'�YM'��o(�L���YuA� ���E�ю�:�s����ĝ���>�����ǘ;|,��F�W}�{��6�O�?�Ѿ
�Q����i/��	�x,�y�xf|����>�U�I 6�_P��X��@��2-<�>�knL���
~M�.|��N��#8��X\��.?�x��Q��42�����c����D�x_�2)�H0�$�D/�D4�8���{�e��v��$p�~��R�NԂИ�ψl�B.�� �����(ͮo����V	cS~�3~�P��<���sxU4�|��0��~/�O��P���j�ٝI�1ue���K�d|L�'��M��7_#x��-i���$�~�b(�}�i�+���2�gv���S��9���(J]�x�榉�e	�Q��21J�����MX�����kQ���H�l�%���sn%��������J����c�)C�x�\���@��WZ��~�Q�3
�8�,ݪ�ܺ��9E&ߠc`��o��H��,%k���ܨ���Q &��>����Xj�GH��`�o@.��A
`^��݁6��~L��`��@�M��R�|�n5���ߍK�|8�1�g��$ځ�(�U��
:UT	2h����W?`J��/Z��u�S,��'s:�̼����V r������6ɯ/�[�`�B?�z v^��a�J�����Wz���Kp6��&(��`���1D���\嫟`5S�6M�{��{�+K3��䁃$x�"�=� 5��gr�oz~�Ӥ9\]D����uv.�X�v�0�,߸߭F��tG\�qTK�r��Ə:vu��<JR�A������uT��e��`	�E蛨�`Vq�K\�kG8���.����7�+
(��F����vY�������f�)���N�pU>[�ŝ��3�)~�� �	��Wq0D\��
L���u����y>�?�[d��'����1�^k\�P�ݵ�{D��%Ys���2�@AW�ĶJ�\c<�o�kEe;x��cc�uU�j-J~�;�@��K��`	��UDՈQ��G���k�֫�D���f�͑W�;;�ֿ闽��j����zI����ȯ@���}w�K~��l��;r,�9yAXa���F�t;=�跙��A<�S6(�D�}��#t	h�wxR����b�=� V����͙sp������&���F2M��ݎ&;I�������ǀ�G�-ҫ	��1̈�h/z%�����xk!
�68�(!��QFY�X���y8�
��u5sZ)gp؍�4�q���m)Q���T�1��T��P�g[�6X���s��h���da��I�c�R<����fk> i�"�xC�e��e����#��6")��7�Yߕs��9���O8�6H�k�����5n�*B��Cf���n�h�����.��eP��z��2A���y}����[X�0�0T||�D��q��إ	�('r��+�;@�F!p0�JJh�/R�S;_�N�h/p���F�%޼4�*�k�������t��o�tR?���U��w�+םX^/��Ι��t㬉|����&)��H��#%-��Š�n�_��f�P�Xu���^n��*��n;g��K�A��S_�>U.�7�a��KF+�r�G���9��-#�5Ď�ռ����4E:2�B���r��G��K����IH�\o4y��lQ��H2���W�����c��|���z;����~�r��=�I�崇x:kF�b�]un��g�N2K��m:>��_����>	�sFyj������
�21@���@�s��:_��*R��W��>ݥ?�a�ɬ��Sô,��	$�~�W�Qg�wi�ϛF� ޙ>˓�ڌ�ԥL&��i�z�u,�� ��s����}ȃ횴VB8���]$b�j�'�*�@J�z);7�uR��?���*]���_`�4����`�8�tȁO�`ne��; �I�5�����<�,B���,�:���$Y|X��{JJء ?z�P�0���soұ��!9E0���SҊ���4?ƲmH���<_j��Z��L��K�E7{*���`^[�з��iy�������eA�O��Y4n����V9�e��M$�w
���<�Y8���a�D��Qn]��o.�D�;Wb:�8j��?LÛRC�%��at��Ug�ʱ�dg����Ϛ)���G'�m>�.�wX�ۆk$r0�d����7��'�H��9[�{뻴ػ4�	3��wB��7� ���Gx��C����VM�V4�i쌬�m⭒{�3�/F�� T���-��.�㌷�ނ���^ʌ�Wn�r��57y|�����]8ZJd�����;�l2��#g�W@7gS�6��"H��\_j�k�M���3a>:���4���j��>3
��`z"4H3m�f �@H���9�d�1~�Aa����0]�������F7��J`"��������4*Es�J��e
�h��w��z.hW���.B�t��te��mml$���$�1V��}���pK�u፲X�/�c5�/�!�-�J�Rg��,M��Y�]��M΢s� �dGS�fdR��\�@���_����Dv��:�p�l�r+u0uzճ.��bަˡO��9a:/�@���y!(���$���9>U)�}�E��yE���Ɠ���ް�N��˾�+�� I�H"/0z[�c�q�ԠǙ�H� Ք��|1�����_�����/�%�z���Ts�ߋ��k�cj�co���=R�=N�K�VL��}f��d�kn0	��*dD�/����v9y�'�-���`�Y��z��Ȝ��GM��Ҕ��<���x��h(x���o�=(��T{�������i����8x0��0XK!�_[��	E�_\pgڎ�Z�thk�e��'��c  ӿ����Z"�=�-�6-�֑Tpb<��ب/�>�ό:�;�B�� �R����T-�Qes�߿D&F��'؛��hu{�)�-M�f��#r�u6��1
iB���b_5�A��.�%V�4^ʹD�l�����(�2��<c��I�y�@M+�^M=��:'(��T��@�{ʨmpe�|N�Q��+@v��}���]Y8�C��]�h)��9��ѥ���d�E�I�ɍqbk5����h���p�َo�Rm�ޢ;�#gt����$|1�?O����p���o��C���A��	�犵��� *q����N&�;�W�5�bbzY� ��S�����w4�M�'��i��գ��Ҥ7�Ȼ�n��Pd���L�)8f���a��{����K?��7��Z+���X�A�{��Uڊۘ��o���y(h��YW��l�����2�
�/¾�a��3��*�.��
}CV��q.���È�X��L�$2�C*�N�ֆ�2����2A�j3/["̙Pl��Y��Sͧ�҂�6��lJf�d[���02��~�����?e쟽�K꼻j�G���hzVHц˗cg��2r��l̦R#�E��'x�����}�jO4��A[��֟�,)��j�*p*��Z�����κX�dR���%�HR�=�k�`j�$��߀[b����ǰ��3��t��8^Ӊ�(�j\��/"�d'	E��)o���9���hH�5+O�E#�%:���͉�i�>�g�Oi�8��|L�u�D{�TiנK�̤{�l��~Μ;�����<�����b�+�:�v�p�AY������lw��&��!�p^���)�>Dk�_t5��/�!�=D��,A��0���1 �td�ы��}���'!&��� {�1�"���.[�v�O״��t�u��'>;�o[T0�t\���7���K�n_{*�20�bӔIC�[_��Sc}��k{5���sS��ă��[SP/!>�^�h�&��a@k�(�H0�m:� ,&+��
�U�
g<�����Bׁ ��X�����%�r�r;
#�U~b:/��93�V�˼
�w�_�P���qf������	n+�_�!���%���K���H�!���uK����,y�ʹ��2"��D�����M�|�K�F�����
)~��Y��E���h��@�Ê?�?��_?���n�!9����Z&��fF/��Q=q�S�U=�9wL7P��7+ 6&��͖��(�+�a���z�7�TV�eee/�I��)���D1el��l����+��3,�ŕ)ui��lLd+,?)��H������euY0�s
�\�Bx7�cf$���)���� ��"���Q���<��=���$��NH�mPE���d���؂[�U���Q0�A# ?E{i��A߇�=���$�ŀl0�#�k�.4/{>�Q����8ow�4^�R胟��T��jaЌ<����-+��W��&���it���ΡxvK���dd|$�~G߃=��#^��?q�+������)�X�1�?�>��d���ՖP*�)e`�Z*�2��������)�<f+~
�U��wv�|G��
L�=���� j���n���e������όu�;�2
�����=��f��.��L�B�-%�-����3U�ǃ�`�C��z]��Z�ye
�kp�$G *:�Qև�go,�������H��ȧ�/z�~&�%�:�	���&KA�Z����t�L;yyyJ�����̈́G6���~�2O��s��F�܅S�(��)s^]������3N^��)rY�'��O��{�Zi��K�߻��}~՞s�����?t^ë]�6c���M�w�8�[%0��`��w��;�lr�������wϛ,ܣ�J�v�0D��6��W��sO"M�EEzC�aߕ�IKG-��8��A^�����*���/��ܒ�s�L"��Jr`��jb�3" �g4t
}�̥�$�3kL_.��!? �����Y�ڞԣ�$di��N�Y�ʏޅ�ܑ�Cۍ5a�7�����(*�ޝ�~��/���o
4�}bC2���]V���K&i�=VB�#������N��8�t�T��ʹ�z��ց%'�� $l���ոј�}����dL>�Ң'�g���e��e�$1�U�SX�km��޽hn��uP|����Ϥ���1�I1�����
��L�Q7�J.�V4!����k���3�J��p���:�Ĉ�W9se�����Yq�n�Lf�ǜi�ն�H��݌�[b&ͷ��Gn�n�r*Ou:����FU[$1f-�G���@��A=z���y���4��i�t����g0wUg�x���H#��0��)����FZ^�aw!}Y����/O�Y�dS5�<OwӰ�i����ھh s�XP���>�f�?�xE){�sP1����r�T󽎔-q9}�\i�Ԇg��0ͪ�э�]���1Z{߿_)��U�t����ۿ�%t�x��٥�DT
�ܞk�>���x��K�,��g�>�_؀8DRu�j8h�^jBw޶ O�"m%�Q�+)����0��6>μ��{�=�{�tf�$���E�;ىS*������L����c��Lrv$��cV����g?�iU�&��D��S��j��:B�P�Q�.�E�]4�ΓV<����Ǩ��e\��f@��`cp��(��;#��j���������K�H�U�l剜3�5H�70�K�[���>��t�LxY��$^���K�ٴ�����&����^��zFf�1���l��V�h`�E�)f'�Gk����ׯ�O[8�8.��S���z��?
�fn��gO��֛$H*�`��6Yd��E@����Zբ�fӏ���kzg\��	����b" cq�B�'���MW�L���]M�TF6�h؛�9xЦ�w_$�|��B��$ ���;ft�P0�(heG�� �-�[+!��^���ɜ�L�����Q@Hΰ2��aAb-���)0��V�5�L��F�^I&[d`a�TBZ��@���a����3�g��������ڂz�@��\,���U��y���ߴ`�,�7�{ Iw�3���I?��7�a�������`,ϖ1TQ��l,�;Z1@��}���P9�]���B��NR8+�e��9�@���)����PW��A
o���ױ���e��W7�Uh ��]��m̅'��G��� P��MŽ񷼠��-@x=Q�J�^n{�Gx?�\auԇ�N�B�a�T������k�&R�l���X�7S1!qZ'�b&��F���8⸣�}X���*�_0ky���98�?K����J��(i�9�;'���!�KLb7�e�İ�*d0�t�\����L?�4��84�{����#��c<ؓ���G��V����ו��Ygp;��=n�H�� ���>ѼQ����l$*��À�H�@)%�n�;����xYD��Ӥ��`�;��ގi�{v9}�;�ni�;�3��^��5>Rq4;�_��e���/�*��:�T���q�n���{��ǹo�'��l�Pf���I�E�Ƀd�[��cr������._&��gQ� A)��1R�� �� ��>�x�}C�=�o��"�x��/Qx���R��ﺹ�o�f��I�!@�߄wz$G����DuQ�IG�ǌVl��,�_���[ڙƶ�j~��D7���pژ��^�n̷��E�v�|�:O��|a\Mcm�֔�1���-p��� ķ1�[j���6T2����	��"t��#W9
+yM�x�D^#���E���8H�y:m�&$��$A�pW�����
����-��+�b|;�1�$"��[�V�nÐj��.�K��nLa��!N�Ͳ�9ޞ���'�i����R� �푻�	",Q����Rj�� 6*D�N�i0�tU���c�3
�.�4���!�������dv�����]���R�ӛ�<�:.k� �tf�4S̚|������ﻵ�-L���X|ë�a��Y�A���r���NV��qt+�pd�RG�� ����m�8�]p����@�8�_��Y��d�h�J Z��dG=�?�|�p��a�g���;U�|�-K�y��6���O&S�O ���t<�I�R��������?J\^	F@���.�k�ܭ���D(�kI/2r�?&3�rh}�)W/D��&�1�y���{��X?�V&��0����*�a��MUc$��$�t�y2�r=�^D��cl�9�D8� ��T��٘���h̜�b%�w,Ny���R;���;2�,d������VY6A��/d���B!��t+f�~�U��H�	Ѥ4.�$��q�~C4bF��n�}�&$O�X�[2Rt]�=��(��e�c$CBx��#������� �8t��5�gF ��3j��.M{�q�3BA�tLs�2�%���|����~h���{� DW���w�L����3�@{3�Ns�Y!��=���Q�����޵,[��a1����%��8th�03i(���O5ͳy��
+ 4x�?�&V�Ŝ5���Q�\�o��78~��� �#�ji���Ъe�,��O�:?�II��+9���]�o�(�g�'7�h(1�w1����s)�&�� �OzE	6G�al"�עB�˜CQ����_i_�8x�M�tכ��W��/T/�Y2����7&�w<L�.x�:\�9�
��+ze��;��S����0l4�2(��~�sX��Qbq|��Ϧ�yo㷈-�Ï^%n�^�*y���T
ZC�P�.#!X�Yv�hcS�ɬomb�ב1��6��Rf����l-^S<f��x����.��~]�F��-�;�֖��(����5��O�GAK�2N4���~��.
�e���m�ɪ���w����e����E,?�Y&�N	��U;r{$��dv�r8�f,��<�>P�!0�m��(�!������pe�.O���JW�<NE��,��HC| �3����V2蔗���J�j�� vI�rD�9��um������s��Y��bg�����6%��,͇7���o?Q�ds��^�7��>hY�G��hG��0��!����c�7�ƮS-fR�dH��/��8~��,� �p�>F@2�닿^hc[!"1�J�F��Q���ͪ*pb���}A��9Z{�-��D�mM��o�;ov��̅�����50���iP�1������,��W�����:�ZpP+�I^���UD{�Un�<!+���?�J�{U��t�%��T-��q5H�!v�.t�U)�ET�T�*n��GP�\I�htu%��lם]o��~�a�Q�SU��~ �yp]լJ���j�:��U�W�%�� ��M�Y�-��A��W��\��^�?�y���+���<��Ͼ�7�]]�e%fKp��Q�aK�: 1�I�HT�3���뵋߶����e�Z���r�D=����a�w-n�o+ ��x��#H0��@��܃�d�aPO�~��9����2���Y����g�FY�s���P�R��V����C뉷�y�]���y=��ؗ1pZbMk"�Jh[t#1+��ō�Gr��s���H��KN�翽�_�\��m�IX��bD�����
�QX���������GW/�x�_b��ĕu���~|%f�(Z�
Ð�K�,�9-���N�Ņ�@�Koo��*]�f��ac7__������G{�D`i��,}�NnY��j������+��U��"�Ml����Da�ϧ�)$XkO�O��p���FG���v�W1���6��ۑQ/�jx�y"uR����z3�d�]�h��cJ/�&��
u��g��j��#��r69#�J�|eK�N�������EM_�D�_�+	qq@��I嬊��U��	큈����Ƿ��� ��\k��;J#L�sQ�W~B����AY�Fs/�8�h#fixf��w�ȧ�,��m����,N�ts����������4���%��|���
�yj~V�|G�h��pL���$�{O�[�V�'�����A���S����9*�7dײa\X�8$_��>��xg4!� �v�en!s��
��N{�ן��"ZG�/�5�:~~G���cA�R瓸C��������r<�� ������>�߃�^���q���c-۞��������~��7u��:�����Gun�er�Бҿh�|:~@���)[���Fg:S2����Q��\L4�]��.�G��|h.�)�S������o!�)�+${oA=�����=�i���B�WV�{_#��=���!�����#�G�э9/�R\fd�0�o$�.�Ϗ�7Oe�g�Z��M�v�_4���Z�����t$�2A2���5���"�3� Oe-��yZM6gQ#9<�P�3"ø;��n؞���m��JI)����$���`�x#'�Wϡ�ku�F�p�E2H��D�E���
��f���[�T+Hy� �Y�j� �CL����֜��-� �bhPGigg)�U��~	�zV�W]3H��
k�6b�{��6�չ �q�C����xU孔�W=_$"2�Jf��iPL�yz���rv��]_L>D�aP\	p;9xu�n">�uP7�5B�|��>n�1pG�#�}��f�KR>F�mX�t�G" ��&�+�%��Y���F�?bM�t��s�]���a�&ub��kb̻-y��<��Y�I��[��%}��WN"��?�}Ҏ�0� ��:}pkw[���-�����R&��Ƀ�Fu���y�&B�ʁ`cO*�]��}�7���w%���ʄ| �,��kp��zW��n�|ha�&)^�SYby���u���<Oݬ��>d�9	�-C.�K�^uZ�Z�QV]"���c��(޲c�P����7�e\}\�.�q��I���&+f��2�����V���h�ϭ"-��l��L	B^඙�6�,�AYe��Z��ıכ��$�F�i�e�FK-j.�f+�]SZk�|7�>
��eKp�!'�ѱ�Q�AHE�����Ju�b��g�]�S��}�oH�U��U�:^�zmd8����Z�Y٠s��m=,i �q������dk(���lظw8��������L��5�D��ɒxh9s�A@�S���n�HD�?h4�qJxF��ц�y�a`�>６Dd����W̆E�O���F���輆[�c��'�O����*ؿ��8�))V��G�o#!��h�[�I�gf�P��0��ç-�>��T>a�*Mo8�%����uĐ�86���X��y��c�T�_{�	�}��h�]�N�?�T׺�ӖW�e�$
�M�������%���(_�+i?��@�;��XHqE���D�$lX�t�G��E��Ǵ'����Nw30D"2D#��g���Քܱ���b�[k���#�d��(�k|,��q�]�3��o���a���w���O���q�e�p�0��<��:r�7��4�-�u��wF��8��+�kef�Y���q�hv�Ũ��F-�����EZ2�ۊ�>�V�U<����:������X��3��.Cj�5�zRK�@�qVYp�S�@�(~[���]�J'Z�ѵ@��⊢{/4���n�^��OTr��F߲��	�X�=�g<��j��	,�@��æ�>{�;�Go�j�<w��� O����d����h�pK<���g�X�j�-��D��bVZ[m�.6�� B�3�y����*����f�P���re�ZQ��y��u�-��abY�)�Q����Vʑ9�kN�~�^�I4���ay�4�uj���)�3�K$��g|-��c�Y���(H�-ӋЄ���8?� 6�J":�lU�{Pd�`cQ��#%5$�|���l���*c�
�ce����l���z6�x��\��$R���Z|y3��G�CR�+w�ۉ��hu<�ɦ�dq���u&�q[@*��ը�p�/ęˏA׸�'�c:�n����a�[�RO#�Aq�'G�9�g�����$Q'D2�� ����p�S�@uͺp4�TZ�>SR�m
ck�QxG�;��=U���T)E?Y�.a���X��Չ'D�Z}��Y�������[�8=j�얿��y]���()W��Rn�8���5`	ʚ�XNV�(4W�i1��b0�u�����.�DL/���s!v5�k���' A0���>��g�q=\R}R�����n�m��7ߧ��r�2�vӖt��\� R�l��d�p���u^���,i�h�������o��c�V�~�&Zu:����K�A?ajQ���.����K?�嬂��[�8���K��7��x���C-R���Vle�Y@�Q C'�����VVZN�I\s*���;��5��Ш�ZQxb,-+�滙��L����S��
��'�k�:���������E�~C`��4\З�:1q}$���,1�~�˫����PMѣ���V��%Ե���pf��"�O�S{��TJ�J��[�9��J�7-�[w��1Xlg ���N�Ep��)NY���3?����Q
[�:���*���� ��#�����K�SO�Ӓ[�+�fn�,tW<E�P|l7�<��Qym��J��]��J�C����m(5���,U n�C�FU쎢�U�gI�x�9�*�s#��i����p�N.�*ZOU��3Ka��Kɐ�°]�\uh���!Q�ݡί]e-���d���(�����R;@hJ��\�1r=�]�I��Gl:bB��RE{� b����N�ю�	��ÿ�m��#Hʎ�v�ۙ�>�^�Q��
��)���9S#)(Ζ���hJJ�0�P�u�B���[wÏ����+>�"=��c�7r�!$���QB�e\"K�R�2�a�N�/�j���ئ(I��}������hK4<m(Q7V�pǳ��ǫ���}j��/x����#����і.ąC��<IbU-I%��LP��t1t��Y�MX�(�q�R�����	����������pA[gy�Ɗ�*��\�û%v��O�UR��|,&5�d֏���<��]L���T[۹H��<�-���=�[G�.��a���g{�\0�&k�������ȃ�`�:�'an�H�I��G�G���0S�1k8�5���P�x�S���
���rG��V��O�?�}f��� �
{��zCs�0)P��j$o�(wUƜl��� }���{��tTal�A&��m�F���#���`+C��־��ݗ���.i��E� �s����C +ч4��A��\�(�vnI8��,Df�pn4��@A����,�ř��5-�����aϓx�M��{�CED����7�}�����܁��5��7�+�Ē\��F�:R7ԗ���"O�y@e��3d��g7�!����� _Yy�!����/�^��í�D�,ir���y#WQ���p�T�k�~��~���bIF��n5��+������:2���"C��j
�Zj��S�ZP���PHY���5�F"�- �΀�
x�_E|!#j�x�Ld��.T8�:c�\6��!�rD�>Y!ꘈ��w��^.%��뀴�'N:�p�x�9�R.���(�_��wD�d��r`���r����^����<��5>|Lzo��Ż�K��2{+o�
u�燾5�񞿈L��.;��,�J(��f �������j�3>�՝����^����U��~�u����ҙ��1�C��c��I��*�0 ���]����y������[�>�)�-hY��0��Z��J '=$�Q�E]Q��xp���&�bP�\�����'UL�s�ᅸ���0c֫O~�!�1��8%���SUf�xf݈�-G9���u�L�S�Ņ )*3�_�r�T�㚉;�\ٜ��;�A+�fS9�~��N�ю�P)HЪ6}��7�?��s�ñ� ~���/�>M
%$����Fn�/wV�v8�v��R��P�U�J�ӽU{SKpcz_���#��=]��a�f�����d�[�lg�V�C�Y�섩N�gr�դ��'eL^@��fh\^���a��(�+�Xt�V��4M�e<�z�O
x"����QO��w�B�S�)���r������f���2�;9h���. bٌ�M;oOm=tZ���H+�<ܨI4�Z�ܜOjp��H�w���Db��?���K	30m��' LsU��<]�n�א�d��LL�B�@�r>BAtވt�x�X���A?�&��gtJF�������H�棦c�~�x~���g-�PCX�����c�]�t.snN�u�כ�4$�S�eq6k^@�i�H($8�s����eU�o����!��������_(��0|ye.�[x�a�%�Z*��:���Pn���m�U�>�E�'�<�3�����f�J��x_����c�����k�S�V�~�4;�%z�e���O�Q�F��[>�KJ�~J"fˢ2��aZ >8�5g7�m�#��7��S*񙶀��D0e�U5VG4�q�r~�=00��@�j�#�lf���i�n��S��������������2���'�R4H͂�����,VU�u_j�R>f���ϜA�24k���A���_dʥ�-�v�qǗ���j���O�� J��$&52�6�qB�fȧ&Њ*첸���wM�Z�!�&�J���֨����g�9�^�b�%�|�]���ʝXV��/3�{{��UxB?�W9j�j�ё��J���I�U6d �7�Ys[�z4����8��0�Q��칆��QNw��ء���ω�]� �����u!��5��B�Жל��
���9j���~�x���嘁�<��B���u˝N�5xL�{"��S3!�`#���G�:@�9���jV��zM���.k(��X���J� ���q�a�+��]����<��7'�7*-~�3_=Dlg��PӰ�iZ˞b��s��ַ0/����B�g-�wu��G�\���'��oA��z�y��:I��j���
�ޞ�D���)3K�d|��p"�lZt��8%]�09��sR�/��6w���Ip4&YaKGl��>#�.Ͽ
����Wv�S�#��.�B6u��sԀ�Pc���J<�+n���!F'S�;��J�8৓���f0a�ƘTRܟ�lW=���ue���'-{�U;�Q=�,J*�ۜ�*���?�x���vTKN۱ޕ6�����pP>�t���˺�u.��v�L4����_X̹���lYq��f]�#�J)�؅��K8D�M�5gA;�
��R q��6�:��m�J���v�L�t;�"��ε�N �Ó�s�D{�Ԉ�8�/5J����	��!WQ�_D��L���i���(Q�(����4�k���hÉ=�2��q�� ���pjyο"�ɭ���X����%�rݑI��$��`�����#Ԏ�!<K�`D����d�y�;,�+p�	�/�_�Ν]	�v~;Adb8�d�N�I��|Y~$��-2�<���� �uQ��3�tc���'b�De,�=�J�������eο�"��a�Ւ������-	�����㇦P�(�+�a�G�;�<���P�B�{�L����XH,U7_|=�� #o�:���8����We�g��(m��`/N"/=J�YbDXE�&����c���x�V���-��ގ�%��{�^R�C<���������k����>̕��V���k-M��4��wFG��{�H�����su\����T~3���@��s�-Gi�:�+z��h�$ V�����DR�>�u}�������u2;�P�a�ܣghn
����p��t3��~�!4F�uGj���3/� Q�V"z��j|���<Jvq�{�D��S��/HC`8�%�\j֜����VM�T�'G��/���KpU_�k����e�� ';�j��1['4�Q������dJ3>�ϐh�φmn�hh�|/����	|:��P��>�>��u�JC�>-5����O�Hfy5���42��fWly�h<�apx�aΠ����q�QsG�W%�!6'	 B ����t."@=��͘��A��J���`��=X�o�w�}�J��=$��ރ������#���-X�)�%O��e0�2ubL �V�r���'q�9X��А�S�.P�2�Pp���O=��O�C�	�a�y�w����S&���s�<T�_7�.8��1��#$N�D4��X��-�M���m?A�/��(�BHoq�*1a�8���Ռ��C,3X����ՊĚ��	��0�b:<�xz�	��j�7�Qd%����]*J
���Ǽ}�
���.��[f����L�c�r_�e"6�|�ai�g5<�=|���A�)P*����WϷ#T7��pgC=��F̺ʡA��0�O��(�r`��D�p��D���F>\L3m�Q�+�9���E�=X8�"�(�g��x�M1A�Al�y�ct�{�tHq������q�J��EΥU�$(�J�#��C�
s�v�N��-p[a~�oh"$�S?�����Ec ��=K^}�C���j��s�t�����A�qiy1ڶ���L, /a���w�
�k|�H�a�`7�ơ��~ x���&��D)����*|x��Q����r|֠�A"�E�Ls��ʞ�=����T�.�ṉ�Dh��c�,Z��Q}+�0Je��֥g�gfM���$4����I�	|h��=Z��1���n�G65����8?��1Z��^TD(��5P���/�/�3�Ps	�^4�&�prhs˧L*�:`�c�΢���\���a�f��DId��(!���q{|;�e;�����e�ʃ�=��>}���+�-�)лCK� �c�'#��K�	e��D[B"�����O��*�$5ڦ�Q��,
����x�Q����+����������5
*@�,���h5z�Om�%�������ok�b���LQ �����!�ɶ6�U�=b���9��&�����*�ps��E/���IHiw��_�I��tO�>���;�X�Dו��n����Xn�S5)���Pړ2S�m]���� �㯅W�����7:t�F!+��u7��X�,�)er"{�1B�*W�DayP?����S�铇�A�=�9�f
`B���S��
�W��Z���_�
�0>S<|C�W����/��\|%��_ف���Z�����F�L� E,2w`$�؇Q	�XWu�~���>�wh�[�J��
��T��&�#�s�D�����u鼪��o
�3a��d
�c�]0;'Xi���1Fk��s��o���vo*�G*Y���(4l��u����w��<3�T�g��)�Rn��`�"ܽ1��Ұ��T_N�0*����������B�*�=Q���ՙ��Y>z]P���Ee���[�����]�S��0i�R�Ű'n����^����E�TX��U��Q�]�^ x1Z/wy�j\`��aMw�����$��µTj��8���ՍLl:����R���Ӄq�~�q5r2����j��[���J�]X]����4
�!�{Kղ�mw���C�m���j�e�DS�6��°�r�9 _[�<f]1��S.C�pO40��TrC��T����'��wW`��`�-2�g��U�+�?K5g�~��Ia퍸���,�Ü߽@�� ��P������&^G�����YA?M�Q��&���\��_/0������������h��q4u"8��:�)�d���=iT�4#�~3j{��;�_�W{���s�:�!�U�����q�І��%Cl	p��lµ���_!�?Rt7�t#҉7�H�E l��;�Y�|�&V�C�����8T|�J>��.9��8��K��!T6��+��4�^珺���*2-�m8�&���������:�6^(�~�hl�LA�5h�{86� ��+c��}!cg�_EXSO��p����3q����%����i6V�g,tI��I{��dճ�zᥞtI���.t�2
���x�#�cߣ�)�({5���3%ç$j�W`B��X&��o ��Q�?�$���)r[�һl�4�'*�(�)Ҫ�+g:��=# uÌP�/��n���0��o��@{��r3%8�����\����ܪ��A,VA+�#{�Hu�i�t&�䙀akə��U��"Ůe�F����iR��|��m�t�j�X*>'8O륈4B;\�/�Xk^e˱b]��*�t��+_��ʤ}�t����39�T��L����ƙ��ZJ׿��N�
$k�'���a�n���r�o�:�~ ��2Ս�eW`�ysf�[d+�;LkS��+S*�ʈ��Ls����BBWlɮ0�@�x�Ojq�'>�2�Q�́��L���Ku;R!:�����gZ)�n/�kJ���ӧ�X�����CV8U�}���2��٧�7OǠhN�Y��S�s�����B4�����̬��gq#Ȟ���r
W��f9,Xl��S��K���R�z\���-��<7.eBvI�ޭw�����	�%)��"�J�m��������+e��2��+�����������ol>��p��"�Y�$}�8	<��v�
 �i�p��xH�^&�'�d�z��4)�'�\Y"S'���txnGJ]�A@�2S��]�a
n$�ޠ�c7��et���b
�Z�G3�7gȧ�*_N�UQ�@i����׭��-r��325�:l�I�e�^�P�ob_Ȳj �߄`i͇����w��C�g����2��B.*y
�^ښ����l�*��{��.� ��� ^��s�*����=�n<{!�>	�����μ�~��A@y
Ҽ�U��Y���B)!�J�<����d"���i�wM��@�t�7���	�|z��(��#X��W��J����J�LW�џ[��Eg�]\�>�^ 2d��7j�jQ$S�%��,�s�2!KNrl�Aġl:�@�fp�f��c�ي�X7�h��i��gA��b��^�x!�ofD)�1u菫	dڠ[�l�K骘<^�TL�I��vn]��sT�YI2�0i{�ј�S����O�98��V�_J�v����vБPj�u���5~�H���u*�w���%;����]*����H�q?�Y�w'�+�0P�.W��o�p=M:@m��e` C�=]��?�ZHl�A�(����ԏt|�8E>㿕e7��Ip�9<�]���5���B�Y��v�*U�{ݟ�a��z�f�WU��?���t��fp7l�M%�ߪ�d�kC]	�wX�>ئ�Zጝ9'V�@zq��i��j�)��k��*���U�3K�x���*�AX�Uz�(o8z��ш���*f���h���bՋ�R�Z&��d�<����M�盢H���w��oZ��7믒�1`I�߫@��l7&~|�c���?4����f5,�J+�`�Ϡ����+n��*�}������
U��
����0�,9�v�8�=[Т�ܤt�2�?Q#>g�� ���Q=��n�4��[<�Pb|��8���oRA�%�ZyCnЛ�n)ߺv]�f��M����{FN�ya?�r�r'ADI�#x�g�8(�V��P�������u/�^����
j��D�m���_Įՙ��6��<�~���/P7*d[ME�e$��K$
w7�]�q�niNη��L��w�E�F�4�EBw�4�����?�w��=?|T���\������]��9��$�E����C"�^wM�4$_���e��J����
fǭ���Y�/h���Pd�yM���a|<���4Z"��º?���^1�Z��T��7f@�j6���¯n���x�`mdD{���Y���4}� �*���KOZ��=���f}U��+E9�ճ�j�&Eϑ��ޓ�4�	t=?Ӽ�WX��ڙe�	1��Om��\<ޏ��BC �L �E���;?%"��F�g����X�L��ɍ(�������
��ꂘH*<$^o'2I���(H���5<$�8��o6����c�h�K|�q��[�Î�,c������b�d2�s,��l�F,x���*��Ri��1��m�yA�f�.����	b��?��I�������K��v	��$���B�T!U�V��$3ά���ɲdbV!�{S�c|��6����Oe��\յA����l��
ŦB�B,.YPb�$�Z�=q��;�@e�)��eg} �w2sZqw�x�[��\z�`� $��,��1���;]-��y�D
r@�[����F�cZn5���X��n"�I�_F�G�uu}�4�v�r(�1+��Y�o����Cn��35���yQ����v����={���DI|`u�M�n����^�N����zF4l��̖.6H���i?J�f��}�a�-�\n+���� �S�[�C����w9aW��P�x�*)������t����e�R�݌߀�(�䷗�O�u�]���6�����v:���"~E,?�&�I�.r��6w����g��z����{j�̥h���b�+˯k�z<��gt3Q����U�+�Z 4����b�VPN��^�+�a%�3j5�@����;��p�cg)�$��Ty���"Ƽ���c�Ƒ�=�a��9��0�`�|�� �޲�Y|G���٨y�>��V@�MP������*��u��~z��/�(�:7&��Y
����Z���`�f�j]潷�[u� ���v� �s�)��$���m��<
H?�����K.��^i���q����.A��σ�ƶ;~{�B1���F��:��#�6�J�Q&ӯ#���(�`|B�����?_�k�j��Ρںх���>,�d��k��pu_n��q�������&�����#���1�TU�q��#M	-R�uijK�T/�u���t��b��>I�h�l�~(0t��4>2�!sor�zv,�����J���]��M�}��Q����Y�7��mu�wA���t
T��:
- �iΏ�����d�'J%���`\��9�[�����R8g���P&�:�ူ/VT��U0��xUߠ�0W�ӽ��GUL��~�_2:a)*J��Ժ��{i�Mq��bYS�Ϡ_�:?^��u7S����"#{ڣN1�,^%����'Y'��I��I�
^�D�jƊ��CC
��%��R�q`8
%�:�$͇��.�o���%�<�AT��m<�4��'K����e�4��<�T>��}�2��6 acݥ4���m�0�*3��'�Vt\��U���0��k���u���z���9����XS�ϭj*I������vz�1]�&��{_ŭc!��aM���ID�e�;T���*�k�W�����0�1T���a,��>�AnO�� �,,�8pID��'	.��	A�hRX�a�j���Cp��kY�/V�/�I�˂����b΄u�H�����,n����}���~�Ls��ؑ��O��/v��2_j��M\�q�憅�,�յ��w�Յ�w����վ�̾u�1�^�ʸ��(Z ����@ɭU���F%,�.�*�"�^i]�y�ٻ��}H�"�(�|��V�9ª,�r���Xp0r��:I!��PN�N	��[]�H��g?F�Abҗ���� A9q�+��] �ڙ$9w/����y\�%�o+M�h�#	�f�Q�� Fh��Y&qq��l"S�uF�FI r(���m��^�hI���&����dz�Bׂ�s�C�@�¼PbYf~��qW���D٣$̌��D���Gt��w Y��0K�Ni�Vj���M�6��xR����-�p7�zWx�"R��J>vƉC��85}�9Q-��(����Wx��͑���a|����l�?QҨb`�C5���A��x��dY��l�{~96B6ʖM�;���F0�ߧl��>'j�w3*�����Eݰ{�&}ԛ����7��ʀ�I̾���<�����^z���T;a����ƒ|���� ��0"��:Y����^��ۣ�h�[9��B����*��lUe���f��[kI�u�7,�$��V��雿��p�?s�b�H"�����,��?Pl�w
si�����q(���ȑ�ɤ����G[��/��E(TzD��d#�V�/pbI��t '�I#S�l���[azO?܇^�|"�X<�F�"r��N�cg|��B�.�ˀ�����N��	J̔-ׄ� U�6�Ρ�^D��tj�	�PM�t?d�
�8��$�����:0�W��*(q߳EMC.yq���u������Md�����N�c�^�K�G� S�ʂW�N���nD�5f�{S~�;R^�0M6�a�E�ɟr?��{_�*��	|��pSG�ulx�k�oT~�_������r	����g �s�ǹ>2�UsY�Qk�Úz�a�j&�������W����uQm�U��p�Ia�i{𥳐Ǟ�H�ö�l6�$�xm��\vT�;�_�B!�Q�-�k���\�e�����(g��A��� ����w���W�ծ�U�@�$c͞��c�x�e>�UD@u���@`8j��C�,�l���A�D��W��1�M�7�w��9�OkQ��k��= f��M����f�i��_�I��tU?�)!��fRv�P;���R��FH��z���qS�K�.C$��$كAͼ>Ę�W>��7��fW��gtq8��2P��5G���\�v�_j��܋L<JuMF���v�wQ͌WphIbi;Aޏ�q֡�h��C���g�x!�.���7�Np\h��R(v��!��g��$���|��mW���ʊ�6��sP̅t��԰9�dH6�>���-&$:9��O��r�K�W;�ؾR7`�W
�b�E����i�*Q-�]��e��?	eFJ�0��B��?/���f��4�rP��I�L�C"Ｗ$w9�88
�U*޶܇ʷz��1n��1ڞRUz8��ͬ�QWS�ܽ�lx"N����[[�F����Ē�oA�Em�Zj�s�3FOWE�Î�w��t���y�I������Hw�<M����
�g��6V�*E��;�b�m`��z8�f�p<Ҡ��C��o{S�߈F5ŵǁSs��d2�
*�q��K�7{7�����=[<WԘ�+��0M�u��HUA��_��9;ǏкF7�ϛ�����ٓ��MU 0��}שG%a-�L�vtQ������|w(�\��k���}۰7�2-3X���=�x�z;(� �����F9�%�`����� }2CmɻZ�!Y� c�S��,���b�L�i��4��ǉ�S��NS��RگK/�I����&����H�!�0����9�1	D	�� ��{�¸8"_�D�64cvO��{M��j����{����T��J�;ʙZ }~{g8L�jSr{].|Ƕ �v;��_`��&|���
@ܹ.Ȝ
��8�O�ol�n��S�[]Ԯ�o����e���N��(���c�	m���Nf���F�
1-�t	FX�}��c��8T��PH��>�j��܁(�;�!�~D#w�#rG�$�o�(%�  5c`���'p���eݦ���+5;� ov��}������s}��Ie�������:��I]6��#�]��Ȅ
F���tb�5����`�����h�?��3H��i�4�N�A`�<T�3#�k�@�x/)r��n|�m�]��8=�?94.���D��E��e�~n���ұ����Rd���+����<Z�>�|�ע��l��>^��s78�}�AS�T�̚����3ޖ�r��3a�z�3�<��P�22�S� ���4�{� Y�pT���c�]/��zx�k��#�2�e!S7М/�R$QF_?�Ў��� ��P��~��B^/6�]�ʡ�}=P����1�����*G)q:|q�_bIq�s�Ʃ��qE��^��=���w��.�+*!P�+�d�@#�>�]d��T� 7�|0�$�&��ĥ-���C������pxZ��L&�퐿lU�������������TN��vwl�F�*�{�zSC���C�z��!r������	�R�c^FX�EopB� �_kKai(�ALP+J�[�Ie��!��%Va�>߁�y^���F��:~���{ˡ�Ҙ��1����.;H1�E��+@ ������3?C���X�7��2�e��5������KF\�`L���t�`�I���������3�a��#�ऑx�t�m� ��of����?�mܫ��1�O�7j�g�m�ۺ����{��J]�4�y�h��/�F��	�4$.����ū�^��(K���Hق � A y���K� ��b������k����~���Dj�����'��9
�3!�V�-��mq��VK���ud��j:��ޚ�TA�}���%s�JK���3��>�6s8�-�y�Y%�
��.��@�we2�M���8��RR�m��̕�yX�\[��ǌ�D��e�cdӹ��_�\�f/m#�R	�/�"��h��Q��������2��!*��(�7��ӓ��H�C�Gap�ʁT�t�O���j�.�58����w��c��+D3NK���O�ҘY=�2�tQ8�ӯ�?�������:��l������$�h��	Ϫ�`1;��7�/�o�kX��0��P�7}��B��S�qm�ѱ!�8��e^Ո	n��-��m�(շ:i~�ܣ��Lr�%�E=#�z�J�F7a
ǲ 'C���7v'$�U�gn���e�/	�0�c|*��K�7����ڸ{)�	�����+;[
�'kH���|��`��!;\OT�%?�*���إ �V����ŧ�iL����X"6�D7�:�?'5'(>�l��T ��w�^x)3uI����M8��+��6 ��Eq�LR�a������^����Q��9�Ѩ�ޘG3��c�D���iAIr!��t4�])�J)�sYg�FRH�f�Sф��vԼ l��1ƞ޵	T�EW�qXy3>��O-�D`tr�=,hIld-�Ӄ��E����8Q��8lQ�L�m,�����jچ%HMe�Kƙ)=t�$*8����9h����l���(x*�w�i����*m���WdїI\QW����Y�$�b%Q���o�/����kM30���H6[m�ːΘZ��v�Cq�{�&3{�>H!s\W���N������]�iE�>L��wH$'b�Ԫ?��ʭ��tᴻ$�b�.�;M��>��n���4�)�pD�SA������h�����z����t����"�����@1�ť���n�������'Ao#��[��E��kRV��űm�T�T��O����Rއ�Y}�w�� ��I��c!�A�<bL�kP\]g4�������?M8�T����:�HYy3� 0y�	*�5�B2�U�1ۓ��=d�����0�Lʺ�����z�>��B�V��l�}�YhO�:�=j�x
>�UB[
>൝�-ܶ�;�;YE�p�~�.�-��k�b�������¢��$k����x�w��O��i�xKh����d:2|�vF#>�Zؗv4�)�뒈/��R3��9�W�I~��N��w�|I� |�����d_	��[���8���l�K��eoq'�b6(y�h!��KL�F_�ԥ�:༗�Yt�{���+�������4H�G���	��w�	��<��K2!��[̚��q/��^B���:�6/�N���/��y�2d,C)(S	!����.��\�/П��v�VV��M>5>� ���fի�(K`c�Q��X� i��h��)^�%5�~Vw{x�\�!�c6����]�sӪz�r�k�r |�:s�u�S���J��U���z\L�E�+p����"}LF+!ڠ�9�c1���p�EK&+�BL�M�w�=�8	��tAê��Ub8���^�#w����*Zd�4�s�S) '�W�_���4{h՜9�������Xj����^VF]�g�W��C�vՆ��M�{��f�[��o���I��8]�5�Ѡ�@u�f_f���v�j�b~�y���m�Z ���
�!��t�!cሖ���GR�L��e0�Ul�T�"���1gxm�,��*�����R/"�(���^LV�Q>J5���Ǉ�;T3�OO:L7�F$ё����ݐ����jhH/�Ve�hݘ�Cz��m<�Z�L�e[�4|z�ޡF�*ut.f�#"���%��͎T饪L�!ޙ�K��3�O��Ee{�<y%y&m(��7֮��1{wPt�kM.�tKs��!����l�D�-\�W�E��:�g���1�I���d�k8��#��F��o@�2�d5�Ԭs��O7��;i�)N����,Zb}�ՅDR��Ha�N�k6�A����
�(f5bjc��� Y�W�n(0c������49��	ʻ�����{CކUڒy���%Y~�9��لwj��A6�_�S�'�/���F ����P���� �/��{� �f��*��{�܍P�k�S_&�B�I2ٳ��E�H����[�mf���b���J���VկR~�5'd����'�����ęWH�e�J��є9XF>?>�����N��#'��-��jұ��Ȣ����|�wmLjk��i.2r���Q����9�}*�+rٌ���c�;��>��ax��z%�K�����h�g0[[��2EN�EKJ-��	0�0\��g�	t(��	���3��2�ЅJ��������M�ɣ�`rD�<_?x�=f�&4��ִj�1s��#<�jI^'�11��reb�����7��Û����1tVp�ل����z�cC3�j�+�Dܦ�U���<)���wHF�p�1f�&�����Hl���n��3�[�P����x+j�݉%�h�ƛg�,�^��^�_�~�\]�$T�T����JP�F��!  �B4�]��u���s��z]Ч�4`g��	���.��� =$���1zFR�B�����˞��΂C��0���Q8�"rɹ��Hf��{�J�t��L���1�H���*i=+��ތ�t�>'��m�Gi e[�a���i��!��,�&'��>m�-7��Y���ь��K�)�I\ì�) ]D|�/	�����I��9t�T�X���t��h���MC�V|�D��*�����4�l|��HtO�#q[���9c�L�_%j?x���6��H�J`�z
F_fK��_��M(.���
R0f%�X��9��!�2�t\�5ˏ�dk�������9Fe��'��0BBDe�HwH�;~�J~�)Z�K�$���8�����[������Y�ۏIh�n���jrX�鸞�-RK���V;~���})��զ������Y.�]���}<�n'�rt=S�Sq/�=��cd�����z�uR�c��0055k��h����s�����1��-���˽�f�����w�35�2a"�@F�lE�훢ZJ���v���>o�>kQ红�?	�	�eh+�ք����d¦���|���`]6���r8�XΓr�3ڎT'��Q0I�����믭,�d3`8�ƛ=.ma�H�K�D8�TS��ni�<%6`0���J�}�l�du56����� ҥϧhԭ�d�h?v����/_#Ձ���wi'���e�i:��OF,	#I��E�oE��w9�$���JKS���o�T
2a ��Hׁￊ����:��DP?v��:Х�ucn��eX��S#	�}��
��<���͵h4�,�&����\�����nպ��q�ː��ԺM�<�c2?9�2ɍ@�N��4�Zv+
r,gc�ά����5��g.�h�~�Z���MNg��PcUWƧSY@&á��$w��X2�����O�S�3�U���-/�"3Kb�{1�M�����Ѷ�P}�cϛ:�擁�ƌ��D�nw����ޤX��GV�H�b����KS�2�_�:坎��� �XI5O�2; �6��
�B�Q��✾���>���`E+12�.�)�[��*n���o�,aLi���\H(l�i|P��Ӫ�T˾���,��$�z��<vS�}�m� �Ћ�j!�L�+z�D�7"KaZkQJ %�t����jz�Φ.���;�aApъ�����w������>���K�$R���&z���ց�d�]�q�����>���Q��6m�`��
	�fm��:pӀb����X�?��R�Gj0nMw���N���>�E[.&�������A��c�8K+�F�男�w���̙W��xL+#�s�z���\iRY������ډ%%�i8����v��r�*��;�@�30�I{y�ľX�s�О^��"�d�s�o�B��(k�9%f�=`_
d%��fG�Q�ǎ����?�Џ�Z�<�����~Ԓ��}ڭ�;e>A9�0T��'@�������aa�G����t����2�gC$��H��M�&JI�f:E���$o0��3�_V���63kTfzi���UR�f�(���b��F�>�P������ku���*�����I)Z��I[��2������U4����;�b_4\L�f��	L�|���R�t^l�ػ������`�۲_-�Cx�w��&�J^�l��}5�*`��	d���\�W�AX$Z�������ȱ�	ssH
�/V�rA����σ}�����2łRёk2��
���f�YO�q]Ti6|,�d��;?h��,��]�U��叒�#���Oj���~�T�����K&Í<h-��B_�Z�,�r�-�J~� ��yͳ��\���c��׏,n]��7��?��G��Ď�z���㿭m��r���X�6�{JnJ����t��]�:��mt�Z���Ċ�3�!�פA��P�1l���oz��b@��|�9�ز�g�|�%L)�E�i�ܴ��7�yos��@B&�A�+s��u[�{�2>߲7��(�O^1DCvu�'���V���*e����L�R�F1 V�.�p��}���׋��*�978�/��i�`5���*/a�@���6-	}�c�\������A�К@@rl�Tr֝�1�ehF��K�ǣ�b��ِp�	HȼCe%�ȭa}b���@<�������v����Ќ�'%H�]ƽ>a�癍rs���k�G��n�.��8���2�oy�s���1G��U������İ��̔��p������@�\2w��|�5S����r*��y֩F�޿��V��1|���8<۳��;��Zn)f1嘑{���	�^=ǉ0�eVE���xc��3����f3�m�����o�7{�9X���Ur�'܍�"�Q�����r�I��*�е ��o�N��65 ��Wx��������w���$�ڜ�Rc��ͪÌ�3+8�'����CV#�3is!Lr>=`)�|m!��u�∡O�J��)n�q����X�X�wV�~b�����f�	<A_���m-&��R��K^� hFT���돔�[�x���� U�1��t���� B�r����VkPѺ�,�6�	���f�c����C
d�e�E�`�m�˄��m��Ԅ\|��i(O�t�}o�9P$/�r8�e-F蟨��K�C�_�}y'��9m\O+B>�R�N�Á��)�J^��6�'�1'�V�ʕ`m(f��j�_w㸮@+>%��s�,S87i^m����15�zn�U��l�+�X�"�c�gkC�n���9XG�Ǧ�}Y�W���"�
X�h�+]{�K���Vݺ �A���7B(O���nH�D+*e[�0"Ua1�?���#,D�爨8��#8jN./�
쯦����|�G`�'�+�U�G�t��F����6bg���W���%�l��'�����>�i��ϱ������:�n���p�xYdEr�oiU�?(�]���+E˓�[(�Vz<���@j4P;(�`���QO�
��U0����`E�X��_��� f>;���9�GT���ԃ��')[�F����=R~�i}�)1�Ҫ�5 \E@�u��Lr���//��CY�����I��Q"�?���s��<��9�ce6����m�w�rz�q򲤲Շ�%b����k�O���4����u��֜�y��<Ym�qD�YQ�uU&�)��,�����r�\��[�/�oϐ%�u�v�N_<�-A����{.�4�;�77#h5��Xb��p��u�PC&���it� �g�w���"CZs��k>�O���c������f7mh���y+�_��VÀ��$�]?���F��)��F3ڧ��k��5@
7�;�f�[�n߇�0���;��o,�e-RS�+���a�9sx|�c`H����EF`O���ݼqZU$�TC߳w�T(Ҿ9j2�7<�Ӫ�A%3�i,�ȉmdbZ���0��hے.2jH%CuL�rAփ paA�����[c��*-0������ބ�P��Ȱ~V�]�K����]����#���b%ᔫ���+gHQ��s*�(����E�?zL�V�xl��0���~ 5^��Q�ݘ�U��
cv>W�'��(��!��L!Çﯻ�$�e�ES�;<���|��Z�Bݾ�� �~C�V$]���J�A"=W���Rs�3�B�[��x���̹�/��V�1e瞈�a�.ݪW|�z�����jT�r��r�M_��@�Az��4�a#�(�8q�yZ�f��e�̸hk���p�w��������pc �q�,�Dԣ��g찔�4�:���oEoΩ5;R�ʝ������A�o��VG�I��p�uǔ�}2�2hl��÷�B$E:
��Ns�8��G�_,�Ki���\{�1�GӾ0v�)dD��z�X1����bD�#a-�=oۖ�M�iJ�]^��3�ZZ�wT�k��c�р�X{5�VZ���<.	ϓn�5�����Rr��̔b�����H��:�^�8C�>P��)-�̍
�]�s���)Ӯn����/�`���3ӗ�{�-�(X�ې����H�ճ���3��ƒ��FP��u�!e�,��\E�ܶ��U˧+�_�<���F�m$ �接����T����Z�/���I ��A'��S���d&�ܵh�񰯔��[
W��8H��p�'��nЗv��G�YBU�5��*@m�gE=�#p���YQ��t�'UY���ĉ��S��uTuSC���=� ��-�sC��@[}�`��4���v4h����n��sc���g� wad�%̛yZX� Xy���k�^��C,�������:���,���'�>��7�q�L!������=�t5mfGX "���mP�����6N�H�Җp`�[�T�t圄����0,��<+0w����)��yE��$j�b(4֭�U�,W6~�g]��q7���J(�ZIT�A��>����<;7 n=��텳�2߇ąR�E4� ��lO~���?ڝU��6��i���X��I`�ٌF�Y���m�L�#����4"AO���B%& �R��(�g�W?< �dO��Ҿ�,�H�x@'W�8�&2��"ߤ���� �5��eٚD"}�}���B�g��Ss)m�,��L�����U�Y��B����K�b�|�������k��ӐE1�lRN��
z�6g���F[�t�ҵ�[��4T�	�/��^�p�.�X�TK_�V��	��'�\זpi�3m,bf�����#0�s����u�^p;�F��u>cQs��i���^�^��6��q�<KS����C���J
rb�B�d���[��֌?OPQ������O;8��fW�3��:��:Ԕ����^����f#��iӮ &\2I�lA/��K4�,�y���`�~O*�d�D

$ط�S�����~�O�.2��<��/����oΑb���D��z�X0<wF�Ty���JL]����62���l���j�Y�/�:�>���)�c���cE+8|�2?�N��Ќ@p����g�Wk�<�`�R	͕/GQD�Q�1���wd�W�kc�%����Oo9�����k�|��Kt:6l��N�S��*A.�1�����92�#�`"�[���"A�����*cg̣�0�IG�^puL𥼌ӑ��\<3�t�(��XWSf��D8�xI���*�*��20N<�p��d�W*�C�y)��>c1�?��+*��zk:lS�.)4�N%p����"\�u9��cWg�C�Egޙr`l+������{�D0���y�,�*�Q�1{�DbCK��c��b�N��q!��xφ�o<�K�ϓ�6󓆽p�,��8<�Du�%�7;�	�w�a"��5���ħ ��K,���z��ە_-�{�B�G�\�%��t��,�ѕ���O���y;���(�|z����|���bD��j6���pj�S��o�ݧ9K�]�/gշ��B�W5��:�-�*���{13��@�,>�{�]=��`�5��)
hqkY�'ӡC��3��--A@0���3;q8����"X�ݫ��?�6|��g]�V##��m�=J���Kɷ�c��63(�pn��;$�4�����d���������-�-�p�Bv��_�pm�u*a/QKm��
��w���:����ssf-/���\�<����J��f��Y��t�Bny]jlD���}��(��-�xZ�T�S'��5���B�@���m�~#P"���܇@��1��}���A��Y���VC�]H���:�Ш�%@m|Q�R�Ě|��#����s.�T@)�o<m+���Bk+ESw�����Uir��0������?�c�	���z���wNR���֘T��D�`��H�E���M��=Z�4�xr�YD){�%�^���?������2�H�9�\��������b��FE�(���E��Y�3~nh-<���u�P@j`�N��MŞjيR*q�X�4�tQ��,� ?F��	���<�&NZZ��)yF�:����Ѓ��ӿq �H�B4x����C��^F�t�#�)�Q:ơN���c���.FT�x�|�%J�I�����-k��p4�Ql[�|>��|ZO��8@Tr���y��YuQ̪�?�)�����٩�R��V�p,Ԫ���1mC����{e��}%���ȼ�b�v��	��ݵ��˻����:�$���?`�����@�6��+�0�Y�(�xR{�q�k`)2��@~V�4�M�����y��r#(�ԁ���AvZ^��I(J���OW�D�?uZ�]~yr�SN��E���o²�� �����~�.$�~�.If�ԩ�M��1g)�pc��L-�Ep�.E:h��t[��j�<�8��TS{~#�#���7�3��gQع��ϐ�a�㆓��Ն�A&��I�������W��=�,9 ?���޴�U��N3�B��l�_���[�,�ND-Wv���� 
��Z�(F�`��G΁Ȼî�P�0�~���7�rT+�b'W�c:�񟇥Y�lkL=�[�y8��3nw��Q���Mu�_M��Q��<(_��v�A�����	�MXèڢ�5�j�ۖ���h���.�i,wQ�Asq�M-�re_��`�NM�g��L�!��L����a��`���4ԧWF(1Ԉ��oȤ)��dP׷�_����~���N\�фi�g G��Y������;��z��o	���0.�0�-r��W%E������0�����a�z�����:�Eݡ��7��	u��[|�s�� S/�Q!�M��h-�/&=m�R�dQǤB�}��n?,;�N�(�t�� L�׵B>_ ܨ&�� ��"�w�A�o�Ǆ�
�szN��mi�5JO!1�ל_���͊����e���M��� q&\˽���Y���	��驡��u�2T��\� &�Ý�ob��/2�6�H��.�D}��TY��2WU.=2��eTǠ$��R��$�|(,�̝�K@t������V��Z�<�X_'%u�z�2����6��zq}��Ӹg���~��������vO觀$�m��%(X*}��mw�	�u|p�PVc�173��;�鬤B�H9�d��{vJ�����{`�F��R�K2����K�=f��`\u����>����8�j��i���q�6��~�6>� x�'�������<�Ԟ"�d=C�)�U��O����B̙�t4ىy�ZC��GB���640���
��d����˻����<��#��w�c:Ĭ�V�6I��Qc<Wf���|��~P<��� ���=	g�9�̓��V&H���l+v��[8����7c$��CL��rk�`K	�� ���n��Cy�q
\��1 �JO<WЮL��S �ׁ����0�,�x�:>���Йl��T��e�=���[J�mB[��P:���v�WƁRv>%�h��.Wq~�:�d@@4�ȏ̏*��Z�~��u��U�uc
��u-(�fD�cX%W��)��A+?Eӡ��;)�5��>�� �UL?�	_Y�,��&.�@�Fu��V�[���3��`G�\�����O�3�#�!,a��Gv&I�a��X�ĴiOk�z,�:.�(B�ɋ.�q���.݉d@��i��x���iiNî	����L�;�y�7��?Ϫ��@���^5�P�N��	�� ֈ�Q����l�4Ce��7΋�!��ykYF��.�KpK�� �g��[죺���Zuß�B�� mlM�Y��rN��p�����N�+6[D13Xx�&�b_���}�e�g��	V�&��D]L�<����`R��+w�Nz���T�/��-�n+�Ld��$��8���ƹ% ����ŉ�'BJ�)]�-<9�����L�aOy��A���A��������Vʅž���;��q5�l˹;�Vf���+d�E��W��7j�ޤ� =���V�����a��*�2�銘�X�T�q��ɢ���Ƙh�,�IÈ���qvF���+�I���O՞C��28r7!y]s��ntg�@���"����.�wm#˴��ʨ���YS��|�'o
�c��z�N���j�r�T
���SPU~\��s� i��C������v�����]���1%n�����	+j1��d���#M��lF��ֱ��S�~�;HNAWI�r��y�fP�cI�_U
?w8�:i�����b�V�{�L���Ae�馍�t9�]�K3ct�lD7^�b���P� ����{ɛ��+z:e�'E�wF�鷮��\\`��5ݞxp��7>�<I�U!��i��2mwjƝ��v�Ã�*v�y"1�tҫ�~H���>柿��2�+qx��"e~^ot����J9E�<� �?����8�`TuV|!Zh �?BF��U��������@4A����a��%��k��.=��"�.	1�r������(p(�� Hl���s��H��f�䯘�w��\��5��`�����3�5}
複-0\T�[�ҋ���
p>J��&;�g�Lb����3��M��ǫv�Z�5��Z3����\�A�AmS�?>������}T5����*���F�a���beHj��s$r��GU�? �o���gc=�g���&ΡY��*���lK��~�VV���j�3� GIl�u�����:R��G��,��q��.!�0�7���ﭜA
�K��ɻ���h�C�����F��S�GOџ��8`����=�^7��&��<;g	��3b����ܥ�����2�bŵ�"��5�̦�=��H���eٸ���P�>���Ϟ�O�{������x��a_��0]��kI ��;r�j?H쨍^������ԛ`�C�4:���K2�%�f.ٺ4��yn����|�n�}�dwl��ʍ���%�X6+f]ul�cC��fB�7�k��=��Ȫ��߻�.ǅBt�?�=����`=������rY�D�<�Le�6�!x1� ����Di#$��l�w�����	ns/ɹ̒S
 1�L+�}o��		v��k<�%Hk���f�r=��k��q�%yx��@��q��L��"��ۨc@[�����*Ev�W�F�K�Nt��d��#4�,��F&g�+��Jw��3��zR�R��0���i�l�\���SY�6Es��W��8���]s�8�B����q�9�!�y�~������nK�Z!�E�m��PS0^��jN�����Z��v
���>l��y��������B,3q0��wS�^�J��JǤ3-� �"�O�jt�3�H��+�?ͷ��7��?����\�B{�e��N���k	{-����(̄p���	��MV��T諯ο_BcMl�KO>����%�2/����%8]a	S\��@��ugrp�F�r�1���	��֥�dx�D�Ѩ	nm�raI�f�И�Cڤ���0E���v��:�.��e�!*��<�2�s���-�>. ����:J�}M����e�=�9��!�B�Bap����%�7��7(�6���;ߘ������1�p�����#M��g|��xX����n����>O9�8R��P�^k�Rvy�a%jA���QGT���)%N#����jp,�\b���	�M�x��c|�����]C�^�,�h�z4���;2�Z�{w��!x`�>�an���_�x��h��2�Y��z���b2�M�!�}w:rǪlV�qHE��xG�o��,L�&�D�@Ѷ:7�����g㢽�+P5+Q%�h��;�/)�J��>{|���n��o��VZ�k����I��pU�H�uL@���K̷q�c�қ�����r�%l0�K5�}�ؽj���o�s��YgFK�ˀU�ONƴ��q���q���E�CLgP
B6�J1�:@H�U�
-6�t]���n8g(l3=���u`�$ �n�����+��`�Z�h'>¥�.�(��'�w��+nVvs\��Q{�-�]�s�H���`�/�Z]�z8)x�69
V��-���t$�=�(�v!MG!7Ia��V�u�t���zu��;����,��Q���R|~'��qg�D�s�s�]� u���G�P��*o���m1{�ʇ�sRM���d]��]#UK���S�fW,;�k�u���rWU���<��$���S�Ǹ!k��|������"I�)�d�m�\��O��`#˸�&��a�{O{)���献���L�҆�1��E�s���/E0sD���o%l�x�o��O�}U[{�O۠��ki%1����et�w��Jgr�2E��������w����ǋc�S������o3s�Bado����}S� ,+y�ǐ�K�#����rBo�9]2���������)���Mø���"Z��)�� B�*ׁ�0�ŔE<sRR�dj!-� �k-�Rk�jF�9%B������d@m�,�M�f�|Е��[�[�0��� �"Q>ٶNP+�}M'�栖%�z�K3n_�^�4��� ].����@��w�50��b�h���T��R��v�9[�Z(��|+��Hgf[�׻��5�S	 gBzX`�x% ��d5il�ӿ{�>�=�c�4�)W���cj�	��[p1<j�ʳ=���5�.n�dD-̩ݾ�L�3�ӆ�^x�uF�%�rc|���;�U��,i;J%�'u2*)A��p��N�z'��q��`m��W�=g�_���c�����; Da�;��e���G��D��\X�h��h���@��	���yp�+�Nл�iW8d�xpA!�yQd��i˄�룹�ש\�."KP�d�Ǽ�ʏ�����1�(��9��6�&���az0���{�s�D	�K�5`�D�8�Ǟ�\��I�!�ډx�Ɯ�P�x���4=�����;�Ӄ$DkE�����[�pQNi}_�~��/EC�S�4R�h�+sg@�����<APˊk����B����r&6.rS?�V���+��M܂+��l�g;#����0,u��fȳ*�\����
A5��c����f�z�(�b&N������ĬM!��FS:T.r��.M�������zdU���|��!�6�[�C_yÜ�lp�b�?�(q/;��[v�i���K�N"�}���D���w*tۢH�O�|�� ����%�c�d��el���|t��D��v�+`�K�t�%��~?�4-�