  --Example instantiation for system 'unnamed'
  unnamed_inst : unnamed
    port map(
      SRAM_ADDR_from_the_sram_0 => SRAM_ADDR_from_the_sram_0,
      SRAM_CE_N_from_the_sram_0 => SRAM_CE_N_from_the_sram_0,
      SRAM_DQ_to_and_from_the_sram_0 => SRAM_DQ_to_and_from_the_sram_0,
      SRAM_LB_N_from_the_sram_0 => SRAM_LB_N_from_the_sram_0,
      SRAM_OE_N_from_the_sram_0 => SRAM_OE_N_from_the_sram_0,
      SRAM_UB_N_from_the_sram_0 => SRAM_UB_N_from_the_sram_0,
      SRAM_WE_N_from_the_sram_0 => SRAM_WE_N_from_the_sram_0,
      VGA_BLANK_from_the_video_vga_controller_0 => VGA_BLANK_from_the_video_vga_controller_0,
      VGA_B_from_the_video_vga_controller_0 => VGA_B_from_the_video_vga_controller_0,
      VGA_CLK_from_the_video_vga_controller_0 => VGA_CLK_from_the_video_vga_controller_0,
      VGA_G_from_the_video_vga_controller_0 => VGA_G_from_the_video_vga_controller_0,
      VGA_HS_from_the_video_vga_controller_0 => VGA_HS_from_the_video_vga_controller_0,
      VGA_R_from_the_video_vga_controller_0 => VGA_R_from_the_video_vga_controller_0,
      VGA_SYNC_from_the_video_vga_controller_0 => VGA_SYNC_from_the_video_vga_controller_0,
      VGA_VS_from_the_video_vga_controller_0 => VGA_VS_from_the_video_vga_controller_0,
      b_SD_cmd_to_and_from_the_Altera_UP_SD_Card_Avalon_Interface_0 => b_SD_cmd_to_and_from_the_Altera_UP_SD_Card_Avalon_Interface_0,
      b_SD_dat3_to_and_from_the_Altera_UP_SD_Card_Avalon_Interface_0 => b_SD_dat3_to_and_from_the_Altera_UP_SD_Card_Avalon_Interface_0,
      b_SD_dat_to_and_from_the_Altera_UP_SD_Card_Avalon_Interface_0 => b_SD_dat_to_and_from_the_Altera_UP_SD_Card_Avalon_Interface_0,
      o_SD_clock_from_the_Altera_UP_SD_Card_Avalon_Interface_0 => o_SD_clock_from_the_Altera_UP_SD_Card_Avalon_Interface_0,
      zs_addr_from_the_sdram_0 => zs_addr_from_the_sdram_0,
      zs_ba_from_the_sdram_0 => zs_ba_from_the_sdram_0,
      zs_cas_n_from_the_sdram_0 => zs_cas_n_from_the_sdram_0,
      zs_cke_from_the_sdram_0 => zs_cke_from_the_sdram_0,
      zs_cs_n_from_the_sdram_0 => zs_cs_n_from_the_sdram_0,
      zs_dq_to_and_from_the_sdram_0 => zs_dq_to_and_from_the_sdram_0,
      zs_dqm_from_the_sdram_0 => zs_dqm_from_the_sdram_0,
      zs_ras_n_from_the_sdram_0 => zs_ras_n_from_the_sdram_0,
      zs_we_n_from_the_sdram_0 => zs_we_n_from_the_sdram_0,
      clk_0 => clk_0,
      clk_1 => clk_1,
      in_port_to_the_button_pio => in_port_to_the_button_pio,
      reset_n => reset_n
    );


