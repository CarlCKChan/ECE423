��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�+����Rq�����������+�nS�U�F7&���S����"�M ��U���@�˴�5��.� -;P�~�oa|
)k���BЖ�@�o�v�4ߘ<��4�l��D�4Ak���-.b���mC*��D�i�M%��%�k�~&ʳ��0!����nY�qe��3��ck����o��z"��,f�ը��%$���|�;+#�0f�UhOǃ��2刑�Lc�����|��|����Q��Ol�pf��\�4Y�
A�Y�a@��qnNAz�pד��ݮiF�?��'~&{�X�v����H�	���Gʲ���dӤ�>v�� ���K�B�x��X�[#s��W�V��.��f$�n���:Qn��24"M��<48�}[�� �(�5��t�L�6����ئe3Xa�|=�X$nD�H"ď�Vl��⼞=��5��n�Q���6;#٬"I�L���P����/P=�}�㟂���C���?�ZI�r�	5��]%���ē�2FTC�Sh��Ds]鉬�@�0:�?"ܮAۙ�>���?��i+c��$�vf�:��P����LX�Z��+�'��Y�}�G��)��q��ʋ�X�]���ۅЅ�aڴG��i����(ް?	�P9���y�
�����E==6�iS��=م�gU����!��8�د�§���g��d���B�Rx%��E}��8�!-�U��@=�R ��s�/�ǥ�;,'�f��|�<�\W�21u�a���{-��������k�����@b��G�9SK{[O��Y��7�vb���yS�����	�63ǲ�Sr�,B�/�t�(��� bc";W���"-�����?�1\�ؤ'

`�x��4Q.�H����E�l���5��S���kd1��{+Hڔ�խ8�|$�������؄+����)���gn��+砯y���>3T��Xw5ӗ<,�C���   ̰�78ys
7�s�m�MO���_���t�3���d���*�۱�)!܃�9��-�J���.��qkT�*)�
0�Fx����t�g#@p��s���(��ܐ�q��U)ײ�Zƚś�!����qp� }�̚ޒ��	�v4����l�a�+|Eۺ�m�%��~�K~�u/+Em����	����������O�����閐��q�p�4��H@n�� N}���dv��m?�:�>!���GK���7r�H�0O��ߙ�	�N,���;�XG�Hw���2�d�lD��
�ϻY>�R���`������R�i�[~�~�<0�|�8t!��l*�,p49Ọ�2Vj������N~EG8��!S�K���͙�}IjV���l���1��Cz&3���\'(��]AG�0Z}?���=�bLϛ�A��3%�$�[G�j�fuA'�ٰ0�q�,����\�I���w�%�7pc�/ ���'t|�M�-�X3U �������fܨ�ZI	�:�:͙(:��}$@Fۢ��q|Le)Q�>C���ӆ[�1���E=A�	��j��WQ��;9�L�S�V����X�,�`������DY,�m�?��!!vC�yu��Ȣ%������S!G=3��i �t�2h,q�&�"���'+t����L�G��_�/QNvsN�UK�@+���[#��yfK�+�2)��/� =�v>3�(>r�'�(Abz!8{��>�G��Y��ϕ���5�
aiY��%ZӰ^#�KJ�7�_����r�90�"Hf�T�F ĳ#4�˟��?��ف�2@�F���Ƃ����M�]>�6Sy3!����=,C Zʺ�}p���݂�<�\��	kI�O�>�~�?=�jXF[XX�� �\)�h�\�v�GE�hOZ��y��6*I�(�ϱJgٕ6� {�� �l``;ʟ�`F�%{Tѱ� ?I�K�^�?�G��V�}t"��V��oń\���V׿� ��{9q_�� �\���F���LJ�����tn
ǏK�񍱖��}c88+¾R�Yd�]���R�2���W�+�Pw`ބ�������%[E�J"+�����q��0� �Ȏ��vML�צ��g֒��3��|��`��&9} ������\t�y9��w�*���k�[��x����f�!��캩�G;�ǻ
VA'�XS�B�g��ҼG������~����Np�*�G��F��|zH�3��t����d�'��Lk�p���1�~'QB��A�v�ah�[����7a�yJ��ӻ�t%-�0ۘ*�
��>(�޹-�=yG�?KK��:K�~�� 2���j��Xv���d��=��|�8Z��F���약_��䋨��8E�;���I��|�j�+�����h.aC�i"��j�T�y�F�>��_qS�,�j�*9eG2ʺ}��-f]g殺���-�hGk�ViR��q���~�l�_��WX^��"����{f��h������ԁhQ���×���uC1���������������6���<q��L��TZ�r��|�&�ҫ���|}FJ��T~KȪԅ�_��H�-u�x_8Fg�<�2���Y �CW�tnO�HZc������}XD���u����M��r�!
��pi��R�����{Q���
����ک5;G�d�Ƽ�'Z�%�����\��5B�P5��*J�{�r���N��J�vlF?�/>�V	��Rf��)�2�RX-���}&�Ө�AH�t3�����Q�/iӢw	wۛs1N���#*_�U�A��ڂ�ہH�a6H�^�Ѐ�}����Q
FQ�2%�c�T�������xD���#H��H�}C��K�ܿ<�a���-�0K�#�����@PȖ���B&�����A
�@g��~�^���XR�E��Z�'�=�8�v{���Y�^���"(���2 ('�a�7�ƬR���r��9���s:��<�."��ʌyP�mE�ۃt�^�g����y~�H�ヤH(3)�k�9E�J^�l~O��'z�?��v�I���LJ���<��>�?�k���U�m���pцpbV �#���~hB�t#$etU�m��r5l�l�5U�v�(_D{���q�����7��˟=��2T�d�s�K/٪7ԓ�^��� ˠ�?v�jץ��)Q����,�ͽ������8��9��q��v���H�͖҃0��L�-Õ$7���()?����n��P���7Nn[igx����ȡ48xm�ɴFju,/RVu�0���{k��̙���?��И�}Q��ے+9��_t&�O?e���K�)Fa"lx��&����P*��e�����"�U/1���Q*j��0�Ö��"_�ֹ��goE1
l�P	�ދ�걽69�щ��	3
4����ﭙ)�U���T��H�dҽcͺh�C_�t����,�,����4��)A�f�=�d���\���x9	tWU����h%�p -<��˷�7C@�f������k7`ڋy}�!󃩊p��窅���V�LO�6e0���V� �*�Y���0ltδt��74�ϏM��j
*"8Xkr�e�)�W{5�#�+������M���Q0�mSZ��8�{�[��kܨ��h��N�/�;����h}Y�)_�f{p�o(@��������c88bUej�`o���|�,�#�P�&��9���|�Oe�;���4	�O�}�ẎB ��Ԫ]-.�Y���A��_A������2}rO=���R��&��g68l�6\�!�n��YJ�О5�q�t"�tܣp;�t�ctд����i�����ԏ�
0v��%C��	��!}��)��ͫ'L��q�ɿs�����d�6#�4lr-�}�m�뮭������B�{��ON9v2������׀W��c�����.hi��g[��i"�Ш	�q�b�Ct�
��s�|�A}(Hs��(��p�R@��ړ9BӠ˔�]�`$�-�K�C���;ɹ I�;P����x\\Ȣ��*,A����j'�(���N3�3֑�ǣ�jF���]H�&�聪�:B�I�
9��L��U5�.�F�%xD���1�Y��A�۶�U.#�I/p����D�ף���B�JQ�C�
<�/�y�����ܤ����|��r�:�~z�G��_�MO�K�m��i:� 8θ.�FUo��V�'^�ꇩC����9�UM;���^{�������˺�E�Jmh�5�]��}�{#(U�1\N�+�`~�1���~�:�SМ�B�>��HاHB�_�uЉ%�1�>�5]�w��rHD�V�c�egeI;�/��6&98E��b�e]q���H*�$ѱ���{I���\�dhI4���O |�ś�t�uӕ���	���u�Ղe��.�?�ڛ;�.	j��!$f ��0I����R���[�#519W�/��]�<	 H�[fhE4�Prs9"J���F�B�/��|᭒����an��L��
4NV�(m�ݗ�:s�xU�}�쁆��W KK � ���ޯ��['>��9��:��_�VV��/�Z_�EYd�M0e��]A!/�m_C�����z�m�ҽB��Z���q��(,L�ˉbj���H
�������B;��0�Ă�Y��p�=e��9�
乞1:���X��lj=��L�IR����q�q����=�����Rah�2I�k� %�h� ~9�)�������aQTn�)�P5n�~&�d�F�y�j�>�D����v3��،�W��C%��p��Kn�K��\�a�pY_G^�	݁;☽�{:���Ig���[�;2���St�jA~��ld�G�Gd3--z��Ii8�*�
�t�
��.Dؙ\[�"?�Y�#&M{�-�I��V�܁Y#����G7qDc`��{�l���e3��(��9�?���A�x�YD��� [\�8�à�k�ӂ���\ZAH�G���җ�?��3��4�HI�sy�c�P���aӟ���9���dx�%	0︣z'��zm (W�s�.���Y�a�B,6�,�3?9���`�PˊQ�V5R�B�w��#zs�YK�l��}A����*�'�=�Ǔ~) ��AJ��8����q�:O
_v�bK���<,?^�.	3CK�jQ�<�41U@㥑���"n�$��9]�,Zy9D��e��>�H7��J���te>��e���R�T������ٓ��ܪ�P��ɾ���v+�h|�@���Ѧ}���2rΞ�>�ͨ�Tk�h/G��,.���p M��>����8�K�}c�H��i�JuO�p��s8�x�f;�E�&�dj!1S���j�q�p\�Wd��F6�mjsq�&��B��{�������X�ڞ�<|������.OY����xL聙B���w�T�0y��37��ƚ�60M�Ӛ,ݢө�
����Ϗ�G���|�����;QX���}B� �[�z�љ�.7_A�03�e�ؽA歚������Ƒ`SQ{Ԝ��y����e��W�ˡ>X|��[b@M�qg(���FC�i�ϟ���v���@T
X�����K�-��{3���{�I�$NT n�,�qV�����X�QO2��LH>���+�&���k��n���`��~{Z"<�y]7�2v�p��مx��EDG�P	��G��1���x��ʷj���Ȣ����Sg}G�8̃����̪�����|�i�-�"�D�]�F�S1�F�Ư:�5Q��Ζ˫��R���a�aB;�{�aO?mF|��P�u516럧��}y����ނ���uv�o�E�h9��6�yt�[�2>���\��ug'*3�{�b�@���G�76�e��<�t)y4}Gg�~��8��IͰ|7���V\%�W�qЙ��q��M�~�A�1bKu�SoM���M���TWp�緥��7ƿ:�nˡ�Cjq�(bͨ'Q���J����5`����Â^��y���$yA�l�S��jc�Q�8�u����21��wQ|Bt�k��8<�K��
Ouj���IH�7��]<E�sȷ�6��S��_�[}�^�E��:.��tL��QD�]H۸n&,-����g۱�:��J����r0�4ohQ�u�?jO��Ҏ�޲'��I!�jE՞�r��ZZfsgc��aF���Y���n��E�8�0L\7V���]�����:E}�]�&ܨ: ���ǌI�x��Yi>��r����[SsRW�z���L!�9.zܒ�Z%,hFk����9�s?d���`��.�rSl�����O�ŕ���*]߁���I��8���i<��Ͼ�0̱�V�[�9�̹I�-�e�SՁ���]>��+G`(����Q։as	�I��_�L�Y�h}VV|�T��@�B��5�f�|���b�l�0,{�.뭺߰�c����?:T���UJ��i�ȑ�gĔ������*���d-�Hw.�e"Y6ng���p��.���j �iz��zwr���o"�N:�K��ɔխ����1��&�a��n�r���ױ�:y����fU��pU��`-��';�-
���2�.{@�a�kp��"ϡ���8�e����xP��(M�,Y�mH9k=�K�����<Z�b}#���j���t}����k~q��.= $�˧3�
���z��I�Z@��R�c�E��t���	�I���H�џ��e	����)\b���^<�/�dk=�
���:n�|�����b������o��K^?2�aaq)�~�`=�[�0b�>|���M��5%ǈ�����s��H��Q�j����c����[�C翷7�G�6�SJ��.f�c5��?FN*�D_7 �f�D�Qt,a*��.Oºi5�/�T�n��6"�d�38��J���5��/2٠"��Q�1-���y�c[��d@��öF��9C7���@��=��_��ޏ����J�I�c/��i;���>�.L��yT�15��ܴ-�.t
�%�������L*�>]�d1�H��?����!�z�x�no���|�SPL�=���I�],���Y
���?����/�C��J��Џ�(�`�5Gjg�>ʁ.�np�Hݨt;�^�A�9gQ��Qv%�D��Iwt�h�=h�UP�r�����ޯ.>���r�\m�H)��<�����UY��-�S�?iA�� ���@8�sL:�$0[����Y��[�o
f"B�5�=Jg�eC��A39���Օꠖ�ݘ��Rο�ag���q�8�F���Bu�	��j�Z�؅h*ܡJ�;�y�w��@�s�r�5���k �c�?�uW�R�v�|lG�xy�*��?�7��j-5�59dT"s�X���:)k�m��
�T6��Եj�J��  ��@V�o4��;�M	uZ�Xe�^k��R�$(�M=*������[A��(.���t#�;¼XYݧ��O5����'#ht\�n������:�����Rs�->��4�s#���M�(�y ��H�L�d��?�7�϶�����22"c`ؙr�HAg���R��P���w8Yz��<xW|tD��$T�A���w'l9��3�k0dyy�3N�1�A9nP������Y��8�rqrX�����-�G!C�ϝ��6��6Iu�X��~/�(���Bq���=��+XD�0�%[��b�Il����\J���5t����g�����K��b�����-)��d��<;�C�8���y}���s7c���C��0�Y|H���!2��w4�9���I]�U�Q����"yK�ڟݪi�"��KH�t�8)"Q��|t9V�A�)@�_�j]��3>���kISձ3��}6x��E�@�=���|����<l����[��H�U��.u%�;q�C��S���2�����5yo�#�M��p���{cV����+N�P����y�?�J�Fn�H����tj��T��1�O!�����>��`5!�r,E��!��E�oC �/��H�*TL����0��� �ϝ`���_��ck8O�c��Q����/�Dsw|$ҡ�&�T�/>t���b�U�����Da�u��;
B)�ձc�6��m˻O�m��#%.�T�8����Ww�͂ն>�[��icx58"ij;�??�y����.���p5ɲ�2J��L�e��ژ.:�(/�
������
��ذgiJ�g�'��Uǲ+�3<�ރ1�hϗº�-����:�y\�y������A�w��-�8X)A=߬`;�ҢԀ6���L-M�����=E�>��ݬ���>��(V|���C��l�����`���IZ�!^y��H;.\���̚:d�%ȟ��}�}L.�ƯY�e�y*��V��3�_~32��7k�/�ʾ�Zݼ��g�1���������'�n�Km}4�1}���Ê!y���xf3���^���Cm��B�=h(���R��).p9��]0�H�>�,������"���w�惻�pt#���"x�9TC˧�ۍQ�f'?;F�`�N����<|!�5�h���� ~�{��Ԕ��[�1�|
^��zɓ<�q��@��]�e���x�M�A[�`���1�Jq'I��3 �c�C�q[�V�k�:sō�\�z�}W�]�G�0k�G�YDUǌ��t�0/}!�:�����r8��1ú��� �&��}�!���G�L���}C�y_Ԍ'����x��&�Q��`DOI�c��3�#J�,��[	%�_��(�O�_w��X(-�/�r���2�]�/grB��~U[�M�&D�IW�c?uw�թ%u����1�\�������&Fi4oW����ۘlSI��)א�<��]�&;�P��`r��5����5�K��Ω�ԫ^��Tn�K���q�|���gԣ �n��="���)�״c6�dk��^�~��z��m��cJ֗�nM��
:W��ݺ��&�
F3r"�ʆ�qÐ�Y�
���:-���p��ƍ��	,A��1����3�^�0�����TRl�����'Ca1����Bh�'&n�*�mP����/1�C���O��7A����0�m9\�`���%���|�S\	(X��ewn����������j=��B����`ddW�$��ө�(�}&#�S�D�w��\��챺����I�پ'B�4��z���ԠX�K���@$�'����q6-5�DF����-�X��_bw-�=M6��>���֩ԓ"A�_W{YO_�/�ύ�-5��j�?�`t/r�Ȏ��2M��� �7sנ+�gt��{���F]J�� lb�� �Se(�u�3�� |�.������&�T=M���+�A�����V���~��`��+�sX�QXQ�v@5�/ν�G�)�|�C������6nܿ&�$	���j��``U����
��5��P�C �t�S��L�Ԗ�RIB����d^�� ��~��ྖt�}_TX�2bϵ���������vw#ѮE��*�d��Q��m��?;y��q8Ë��eD_8O�I���b�JW�Mj��='����r�GI^^	D�v�ɬih_���b�1"b���&#V���?	�����3l5��j��k�~�7�_(q^r:q0z�x��$����:"��[�� �:�i��v�椷�nL�/d����y�	�l��$��ם��-���k=�0+����0U�[��\z�Ȃ�ʏ_v2�y�)wَ�OƦVs��J'5'�x������|����5vL
�ޝ���#�ד@�;�FO�]@�"�Fo[����bPmͣ@�9����m�E���[�[{�+��J}#,!� �<'Yv�ߛqqH���o�kH�$c%����ߓd��\�4Pb�@C��h�������ȑ'9ׯ�lhQq�zj�-/��ԥ�^ղf_ͱ�r�.���qƮy�jG��D��6XH���vN �wLN�XR�������͢�E�%�E]�����N}��G�+�DSz(�NF|!EHR�zK�X
S./��솄�@v��)ݹ�Z�陵7���K[�w�yF�_z:%8ךX=�i�8w���=���;}ɛ}h�)�A���U�^�0Sw���&�=0WJ�1����_ ��K c�
��k�z��{"M����E/D�?���m�h��;ξ��Ӯ	N:�fG�Á!8�N����%#���9}���`�g�3��7�q�"���q7����ǧF��tV��[<4�J�>Z�Ȗ',��.�}9��!��w3�Y
��
�mC�v� Xy�$t���{��,�j\zx\��p��1O��Ê,k�x�TY:+����G?��z�K�1�����r 1�[:0Q�r�>��Κ���RC�xn<�w�������1��S����(����, ���p>ǠD�Ќ�y��[����(>� 6ZHv��-D=�P��������ݓ{VϚ!�+ �����8hŤl-wrKh��CNHA~f�c��][Bp���>������0�r��b��S �:��w��u�r�{E��l�@ �<mZS}x�����wi�|��^��Ut�v�~s��'��;/Á1kC�eS4Y
u���"��_V!���]w�koO�@�]�$��eF�ß�K���<�?�D���O|��%D���D92}x� ��60QٚNi��mX��ǜ�d%�o��ȋe��Z�ÝW�rc�zz��l�1c�͏ҧse���ժ���J� ��1A��r�w`l_*}L�ei�ak���j�0B�@}Yϳhg_�$�uH�sc�U�=����פ3�l��D1�be9]6s�7ơ�`5���q������䊘~k�
7'��w��wo>�G��x�P0͞y;�/�^X!��RY2v�e$��i,�WR��cN�ya^:�a{��%�s�́R��+T��>dN>�9#�����~u%�h�ϟ��4�-�||�ð�4�	C|DM"�wb��1F�@<)M�3��u ���#8�t��MĖ�"�'H�r0"Ė�ꮞ������)W�u�~��4T�p@j�dӅ�t�5}T݁w�Ĺu�꛾���H.���v�݈/6���eTX��~w�&��&�~���Y�e�
޺�}ں�_4��>�f�tf_� ��c�-�*$��zG�3)S��IE0�q���W��_<w�
U*�L���-��w?L��t��y��-R�h%C"\��m�c<ᵜ��7f�>����x����]���v�]u�u��ų�B�E��Ė�w�~�mt�W˥����`4�G��*��ދjށZl'���0A�ě�\S�r�-�3�Hg��`&�`)a��������-N�Q� 0؇�ST(�%n_CCv�� �UP�A��#���]Zg��'*�!��a�?i�U$��K"D�}����2��g~Q�+���&��J����L������杄�L>e�o����z]1���{�����9�l�po�v  Jx˗��$Q׷k��;H3���D~ ;bϪy�]��t�F�6��oBfI��%;պ�BH�M���\� �J���՜���;��^�����[i (S%	ne���߬�Ƅ5�����e��<Q)�F7�l�Ƣ��La:��oʩ�.���F����L,����!1��s�r�Nl=�*<8� ���j.��G�q3M�Y7G�������ldg�a�G��ی�>�3h�Ȉ�'⤰����K��c��m=N/�g������dzy/�pf��L?�:~��wr�����լ�R�L�䮌k�,�P�zK��!�Z��/k1u�IV��!�<��Q�R�4��3���`:�p'�FJK>3�\��FC�>\i����w7#����6�F۽�x
3��[e�C�Y�a��j�!�:\����j��\լU[oBʛ�U�@�Pj�������H�o尫��;��L��E �6Gɮ�F�)�KsW�!ev���4��݇���Fe��{Zuv��M���2梉�)��UI%���6ۙÅ?�Uy+����P����Y��0�$v}���ZF��<&�F�#&	!�1(b��IV�(�e���0��G���Ϣ�� y�&+n�N���p6J_�n�A$$������[N�IB���[!�j�54@��lɄ$�ƁB��P m�S�]"۳��;)�{�h<j�t���A������b<��,8��Jxq���cH5t�1˙
�xDD�������Y��Sr�����}A|b�����U��sv�<ӽ�#t�E��KU�7_��^l���c13~�@Z�V�2I��G`�L`V"��~Ǐ�Z���?t晸����_wO�d��;���6C�$����ڃcy��~��ZQ���2���M-''�ejˎh�h���s����r�����l��3��� ���
��w�b�d��H��O��<l�|�,��ջ+��O��N�,p�����р�uGb�6I ڍ����i�r�/�����[�0�!%�e���?<F�f; Cg�xU��Kdj�����*4�Γ�!�\P_~"�Q6���yr�p�|3�W)���7��4��y|�#20z�t�}��-��ۯcq���X�yL�*�&ddz�.��,e��l�8��H7}�"�n�o�%uN��\t�Wh�����4����`�r�9�4u��wz�kV?��s7��m��C���1O��A�Zq�m�J�	L3��󩓎y��a5΍���K��Bz ���_E9�I���$�$�%�yɦ5�4��}�kP�X�����t�����<ӸA!��Ԭ'�{fO��T��E�	��mc�(��)��X����Ruy�9��qYsD�"�0�N��	,-n<Jag ��(��C�p��k�H�\�	�AL$0F�^�d���}Y�$t�ES,lD��D�W��K��0C[r�xoY\\�p+F��q�Ȃ�n����<��a]�I��/�&`�k�di� 6�T|<פO�@u���k�U�a�;E&�,�)C�A��OO�XFf���������an�r�#�FwP����&(D�������%^H�ek1`������0#�z�l��1QD!%	���t���u>(�R������j��*� ��y�(�,S�0i�@d(4L&�כ��f������~,�u,��h �V!���ѺaR&�l����@O���}�a�t/��F技�Z
�n��h�.O�u���j!������CMdd5kܟ��������5��S�ˢE� 1 ?R&��M��g>ek�/�:2Ga�ǧ�C�Q�v�%�<9<uܡ)�߰��r��|�2ޑ��Ϣ(��:ޥo,���0����s~�C���j��[C9�c^�~��U]=�xƽ�Y6SX�1�%��G�)�pUg{~I7����T�u��T��ہ��%RaΞ��oz��Z��}?�W�PѦ,��nB3h5���K͏ ����5R�|��i*�?BQH�D'c�����o�aN��8��v�Ᵽ��7��W�C�H|[j�2-�9N�9�,��n�<�9N�1�:`{��ah�[�f�:oY�5F�F�Y*��蛓��=).�ө 1=�O[�`�b���en�j>��y�$�PՍߐ"�g�r �*�![�օ�����yVp�m�P��	j~�ֈu��5£��������E�۩JZ�5�qe��1z��j�%ǡq찡G�OS�]�`��I�4��Ш:�'�ҍ�[�'�Fu���>.�ҏRAISyhJU�Q�_Ug9�D���ER�BĈ��T��:=���3����&:�\ZC�6�m���vB���		�h�/�=���kw�c����r�B��Xj3ȗ�E^\a���<�����
xߦ�$w,��"�H�R��?s�x��n�C!� �r��T��DܸU]0)?yǐ���!����G�fJC�6qm�$| ��+8���_p�*w�}X�r�K�AD�����ٚ�@��`Q���:�6[���|`?��w�H<ce���I�L��i��H�m����M���R���M���Ң��N�P2ت�!`���>�X�']�fθ�*�A��x�&ibȬ�ZlS��!���� ���������s���2�lє��9�V�&�ε�7��Y���ލ� R�0��!_�u
� ����Ο�Ų:�u��X�����Z>B~k���l(�����O��sv�Iջ�NJ�?o����f8 ��p/�6��,5ƭG��'!8!h�X�P�	��������9Vtvdt��Fr�Q��s��/iA���@5)'�<%򓣸���R��g�xu����e�HW�@��BF�(xm,���"ەn��R���Е��O8Ch :
9��o��8�����2�Z�"�1�g��AR��w�1�Hx��q�A�^�lG��+B�oh�6���ܹܘ���EH���9�w���V`�/�
h�^�w�Z��<�����'����p��������M�����xCEu��"S7]ډ���x�o?��w`4��7��m��N�R4k������~�����^_B� j ��l,f�RFE���9��޸&i���4跨^�dX[�ȍ�*fnqU��;'4�ZK���MB#�a��1�b�l3���.��U�}���^}غ�DF�B�ˋ(��K�v8/D��+�+9I;�̅*�ν�:�n �v*Z=�|x��ox���>��p�B�p���w�)|��sQ�J��ZlKY����/^�V���d܃J��Ƒ��<���G��<��VFA!E�?��
ռI�vp����� ���SM�x8��q�tx�;��+�rTm*�c�$�
Lwݽ�"hq�EHn`��|{}.�w#/�ˊ���B�[�+������ �3I��3Φ�B�>���z���T�#��_���5�A��V����ӥE��c�A:�HMy�����h��&����c�?NqԖ�dQy��������.h�!�/<�M�� �� ���q��FVy��U����S�)F�=����lD���a�(^�+M
��/Wi|�{�~��E�K��Zk=D�3-�Jn{�ue�Nנ�
�h����_CY�Q��j_]�>�3$N^ށ�}� ~��p���G�<*������8��mw���i�@X]֧?x�&M��p6�w���J�}�n�p{	�>��r߅]��̑��J&������<�H/�o>vf��Q��һ�ïR��o�j�3:1M�b�z��1��\! ��{Nvl7�mJ�	�b��CzP��۱����Ë���z?�
�n��Q�?�����m$W-�_;nc}2a�k�*����$�T��B��.@�ʫa������|��(2�F77�T5���o/� x���g�2��0r����cY�v�1�C��q���8�B*�u[/����RZ��@��>z�g���j�Ǝ���`'��R�g�2|m��g�E䦭�<��NU-���7���K�TH�E�ʱ3�?0#:BN�Ks1$,^��H�ps/���j�'Z�]��)kft)=�ٍ�ꜷ3*
�����*�\l�	L���U����ɎwA-� �\݊��Iٹ�m�1�,�ɷ��PP �u\a*Y�g�z.�w���v�V��U��p�>oN���'����" v�e{��]�!�*�O!_"쇭Z�/P�-k�w6+�ZHm9����3��
�%4��oG�᩽�l����<!�{,fN֨��:���V�D���f��I��`�+����d	*�k���5�kI�A�6"���a�[� ����oy�rt閹�Cl��m�׎^�3Yk��qnJЛ3��	u��w
rQ�6g:��c�n�,��9��}���&Ҝ�qW��R���![�4ު��P���eܸ+kyQ�e7���Mn��4X��H�fPBIـV���Y�������j�s����nT"&Pe�d�L�PZ���۸������e�|���4�U1��4fl�{��h����,�<��L�kU`A����]f��XN.hR�~����0Oǐ��x+.�%D�dDK�>�R8H�c����;�ߚ��Ex�&�J��־�����;X��΃�Q���=���oӌ���L��C4�{���TP�������8 }4�n?��P��o"b��ص���n�io@��)yǩC�m��X��CU�i-����sOw����ᾁ���}x�Z�Й3����z5�A�ˁZ�0��P�o\o�
��`Z�k� tc9�'���GD��8�{��o�?f�E��ɈI���i�k���X�풻�hR�ݺ񜋺3Ϟ2����2-n	�6������f��p���0�t���K#��t;�|-,5^tq��¹�s���:.υ���+�"���S�	(8�ȟ�ԇK&��,��"C�C41|��r���A�o;Ē�b*ҤO�?�n?s�.��~o� y�A��,>V�X�M\Y�I�4�WeT�Y\�~�5����w�ox�I�����⭃����MyK�v�'c ��N��ulM�weS~Al$"�Wc8�:��>�$�5u?+��J�1O���ç�؅�\q
��p���c>|H��ԝG#�A��!��ͷ޺W"���vۘƅ>����e���> ��:��@�h�bĜQ�����k'���d�~�G>z2&�k�m�⪝��<�9��W!݆w�a/��^C��\0�!5h'�J���o[e3�@�����3�,R�:L���ݑԸ!QL�db;��sy�S�@n�GJ�fS��o��&Dp��� 5��Zm%���������H�Ƌ���m6M��rTBY=]���*��}�sg!���Fl�_dH��׼4�Fi��S�v>���L.޶���<���9{ŕc�B��6�[,9�s�`J����O?�W��{���E�D�KבF�	�n]Cd�Qw+;�)
�}T�[Av�Z��=�c��xc�=�~��x>ćJ�]� 0� ����)ݚ����z�#E�R���·	Ukse�%
D�=8���4�Re6�u�T���(��`6/x��)lh����wÍ_�}��,wp#�DL\`���������v(��pUoP�MC.�L�c�=T����.&�(�.�:�v�~m9>!�<�c0߬��P�7���"��J�1W�'c�0÷�?%�����ʪPv�=bf�馎��O������д� ٻ��{����3���xw�gXPZKęo�=���dZ�%h�ĳ4�Q��g׃kb<ܪi���o�f@�G�b���'�"߸����`�pM���i
j�FPS�m�_?^��Աh�]���|��'�h�.���>�fx�)J���H�#Y�Ѥ>O2%R �R������������0�c�0@���E̓qkG���nB,��h�%�?_��s/�b�/(@@Z�̒ᰎ��$�S�il��NO���ϟߐ\���rf�[x�����!����(-v��nE��גr��;����V�GN;�e/>A�G%D1�ߤ�ĥ3�N��K���t��P��V�X�����dib+UD�i=�:��k����wˁ��%"���P$0
�8�Y�W��;���3��T�H݄j�g*�� ��k��޿w2�.,O��r�����o��j�!*#�x[�W�]xtDK���V�P��Ra/uŴ9�/�->�o<�4���r��M�X�*e�U�7�ݢ�E�}����>{{�'��ғ�M���R�vB�Ay�<�*1|p��<g��V��TC�E^K��D?�����.�Χu�����U`���Q���-#��D��4b%�����:�N�R���9"5�G��"��C9� �H��.�l�.��0��	�Whu�?�i;����6�9���3n�e,��&nuQ@�\�`T�ԅ�eY��7��0�&��)
���ԏ��4�`��#{�{�0 ?�85�y�=�����O��0�㴩�i���������\�7g,�zm��XRF̸�UP��6����w&�#��ƿK ��z��R:◍�A�K"R�UF��m]���~Jضh���$�|�za{N>1&p��@�w�0�ib���Dq�~߳��Աf��f"}��N��}��O�f59*ꔣQ��N�*)46����ߟ����7͑��V-1��18I;a��YA[UZ��QAI	Bi�8ר�ȼ_�$�2�Ȏ#S/�)�U@��S"�B���< }e�h>:�^��=�\F�}i�6��FՊ����NPw��7�N��M���⿰C����f�<�����&�d%���Y�z�:Tz�<��UϦ��_F �ӡ�-��ę�[آ\��Yմz�b�1��-��@/�<�� �`eX�fK���-���4�MH8)�.�G�>h��%{�=�t���oiU8>�Ctf�P��-9`��'����I�JW���O��Rk���-�յ�h$H�0X*��O_KV�|�v*�96.����T|�	�H��|��x^`�%%g��=�r����;�Q�]o5{���0Yr�`��\8����R`��B�|��7ZNr��y m���gn�����/�+Z4�-=�`	�A�b��OR��HV���b���1P��E�((�/}�Rs�S�8�?.��e����)y�d�f�e?M"��7.�B��I��H��q;[3�v���u~�7�H�m4��&ES��JZ鏻L�y�e�;=�d7��T2tJP���#�1����^�n*D�(�SN���a��W���7B�PIjkCK�}GZR�	Ag*��|�q�Iw#˞R�1�����r���]�	o1[�.Z,_Ig���>ήe�m+^O�9At8T�<�s[q��&�7�!>�;�]MC����il!{	\����z,��5����"�z�X,���Ij�L�G�Eev�Q��n��?���,�W �`�Tc�'�@�ħ0�Q��4����R%k8�z�K���{|a�U�KW��k��:�73�b$��pI%Vw��C���b!,ZD��/�u���QŦ����%뉎�=�B�!��gz��(��I�J ��ڇ@�m 
���@L�Y���i��YñQZ������3�g��=��m"��a1LL�'~*�g�$�l![�����^.)�xeG�,֡��l�i\�p��K�i�j��;���6@&�J���ņM��=+�
�nn��t�W|���a�ۂ�;&Ɨ�r�aܧkQ�n޾wX�x���(����_�9L[�%��5^�n��5��	"�5Ш"�fP�_A�lL٥�+���o�h,O��[�wj�h3t�X]����$�P{�����-e]��Գ|%�ll�oـ��fk�k4�=��'&�X���~V<�M�1���VõD�Ar�^�V����Ȥ/�7mw�k�jY(�iȵ�k�W%�e`}� � ���rp(�5�Z� �|�$�����v^v�_
�J���S��~;�>��u�ghE���
��A�0��#��.�ʵ��ڼnR��x0�<��]�ZяY�;m���W���s�PtFѕ�-]1g����ADr�h��g�GZK�N��!1'�Gˏ��?@b��^���1]4(�u�+��;�!�*��.[�]��Y�������\�%c��WX��sZ�&��2�ȡ�3@/�����a��z����.f�jO��B�G���8iCD	s4f�z�
����3'f���u�/�g'a�������H&8J�N2~�����Lm�$�p��GLJ^�I~m��E�<7�"=��TZn��nR�T��x���鿇�n��n�o.��e'Æ���̬m����;�N6�w�ʰ�`��_ʪ"6�k1�6X�p��2y�(�qZ/_v�Rlh�^|��ԑ�Fe��f�Meμ���b�kin���l�a�-F�	��Ss5t��x[:*v ��}��*T��>.%HF�~�XIU�M���XQ���o�Y��M¬��k�$�M�!=Z��^4 ��D���v��*�CW\;;��	��` ��v���zb�hN�=v1}h�dA���n
UY]�=	���/q3jL�t(��5�uYJ|����.����5	g��A2�B�3+�w�g����O��;ݭ���_�|@����@7���bږ�������9;S9_�C��hb�� �â��K�%��,�1:w��}�GP�ކ)|��9��.�'��+�hV3����{s+^��k����]��'u��)�@!l�K��-�v���iu�fVM�6��L��ښ��1i�oTd��"���,ǐ˰�zf�����}UТ��U�b�J�rh�J�]��<8A�\�8�*���:<ǣ3z4�>�K���f����-��o�HŶIJDԣ�����쿫ٜqi��]D�I��0ZL$JXIi4-������D51E�'�[��0���L�>���������9,��"��٨%~Ok�}���n�Q���:x{I�"�M��E�^v����HL�+/�jMZ������BS��|j%�j� ��Æ	��n�4�e����p��3\:��7 R�jf7R��@k�pJG���?dV��u����s�9��2]ыX����D���4��˴�刐��8��"^MBg��`S�:�*�VD��%�Z���Y�9�H ؗwyN�zO>5�
���C&��q��5��&
X2KnR�N=�{ߨ����DnYG�I��ų]!�'Q�q����,��4>�������)�EeN2\:��Ȝ��OhG�����*CXч21��7��ʟ�{��� r����kD���`��
��L30g�?1ͥn���n���*�!�����]u7��ɱ�$��_��X �,�0R�YO.��l�5�*y�oH�0ၪ���T�g�@$�$��TQ=B��q�8��cvhs����B��n�4�3�`K.�$�^.�4�/E-u�d��˽l�P��6��܄��3����� lC��/j��6�����D��rc^i�<���	�P;3�5Qg��-!��~O�ޘ\�vEv͏/��^%��f�=���SK)�C�� �\�W���uqC�c�$r�@\Scckŀ���USQ~u�7a�(Ėn�A!B�g�0<'����{]м�SLz����RH~I�/7ʉRO�.�7������c�E�Tb���kG�P�
\pO�����C�H�=M~h�Ψ��v� "�n(a�|�Y�bA��@�H�P� �<y+�L;��y�zj�F���~�>�t�͗���h�'N��#��_��ר��B��qV���JL��g{;S� ����%�m��,6H�L�ё��@��ʢ�W����#�����޴��~W�������1d������
��������*�Q�~��������x����)ߛ��>�1$�ؗ�K���#Y��\a<�H�M�KDc����8H�K�O�m���������#S´xf^z������鰅'����_�(a��}�8���J���ЮP�_�i������k����SF����pg�Vm��QM k�����p&t�|)1��_&Q�
!\��WO����+J���?п���Y�'��ym��,Vč����s�t������1v��q�ΐL
���O�>�$w��ú�O��X�̇��c��M��n��LN��VΌ��jM+;La��8Tn�:M��s���+�bʽ"^�9�x��Ě��
���)]_f4�����&�En���;��>��	�%{IM�m�I�:C�T���$��43���w�i�ܿ]�kTևb��m��	��j��_c��"�����w_��+r4ul���|���`l�Ŝ�&2� ���.�9�&U�O��_3E.W��5�ܡ�@�S�� .9�P��n�H~�z��n>H��ľ�)-��_�߳�d�����DĿ���Y�"���SC��@�t�'uH�VIv�'m�
v�+�`�DK�A{��R7� ��g5�1&Vea����-w�K�D�[�����qK�s�#��k��+�܅���,�D4��k�����G��j����崁���'�ٞ�	�j���.d߳���r�b{]Ǒ�)
Xj��Y���N������6Ĵ������%�a��O��7�Y�a�u�;Y��?k36g�B
~��L�*ڈ�:�K=���峨���#KQ�E�&��Ң�]#ΖZ˒��!ux֒�@�$?���a�"�#z���>_u��D�b���Y��=4�겨��v��~��Ѿ�mb_ǡ�o�41� ��|)v(c)���K���/R|R��1��ZJ�>,�������[>Q��v#��daZ(V���	��=��xM�`�Ŗ};;������Q��D~,���,Q�3{�1���R����/T��hǮd���H��v����7Q����o<���Q�#�a$��ڪ%�@�L�+	�c�>��_L�TԖ�ɃFν��"��!�s�6���邃��{�	�Z����R쳾�n9ߕXL�;��!Q[ə�T�I�R���#����2za/�ӹ"���I�G��R!�5�p���J�u�v�j7?mv��\������2V|k˔��޸�0D?f��� �=)��0��ajH����
Al�E�n�Q�����������|�+�_ ~^���L��w����WP�E/���)��*�B�?�t�Z D�?�TT�yq�f�B�G/L-�0���X.[�sh
�c���k�L�q#N�e���Y��#zo���:C�]@O� ���Py�[}����Su�+DjR`�CC�ɓ:�Az����3{�겻t"���K���Al��1�MWc��$��}E�s�h�~���Um�ЦYDH��L�w�m�(����3գ}��md�5�z��n�|�Ea�j�qB�H�6&;�R��Kz9��3�H���.��*�GO�L�oc�r��Ӄ��Q��GZ��D�SU������~�~T�+-�d5�%m1�MJP͗gU���<��Ƙ�T�*�T:Hv�S��4����Iබ��8-+A(�s��<�]/�Q��eW��_b{����J�9MZ��|�r
a�L�;�;H\����k��|P��u�?Eo�>`��T����46:һJ�֞��7g��{��C �9pd-_R����>\̙[��1JN����@r��a��(L����4r{�2~E���D�X��e��?��>E�D��sŊ���Cz({�x�D>WR3��ᅣP����Mk	� C����v#�z��Fft[1�``J�㼿T}�@$�/ѭ�=�40O���Q��*���g��`Jq���H����}�w�EL:���/����|�D���̳��^�����g�,5�ow�e��f�DT�����Q��#�(�Sĺ�ƣ�� �c�1 �@8�J��E�J_6�����j�&x�o S��F�^�@אE����דD��?C���X�m����{�Ӣ�q_,����?�f��"�=�*H�e�l�� �7H�X���7���yvr�� �����:������rd�	�d!`67�9e���4ˋ��q���G܄fs1��
�M����F�z��4��mA��r'����R�ciW^��������Ov��"�W�+���+��:�([��q���9� �6���_j�¸4澳���\�g�i���v���������g��/;&Y�{�|G��$��m�&����d��^�?^�\LpWH#�9�n�k`1�Q����ԅ�����V�x����p۲���&��D��1m;D��ڶ\$�71 �q�WE�A�ڒm��G�	��Q��Ւ���ԒXtmv�2���IV�H&\�t�(y�͗��T^�܎���?� �����7:���)_걯��0�sn�Hd@�L�^��tțO.��m@,��K��Y��<��7��H�W�Ě���z��D��������?��p�l5V|&;,~�v[��ўS&�z��/�'��!�(o�t�i��P���\>��Z�����Ӥ����I>I��3QS��c��>E����������yD�?�ؕ���K}�ݬh��m)�<�:	�9��]utn��|�6������c���`��5�\u��E�:�xZ*4�F��b5�{�2��%_�F?�׼b����D����k�;k�-��P��A~����{®�� o^�@�G�x�+���+��;�ߛ�VIk�Ø�~�4m,I�����B5�^��l�����/�ҿ23ऽa4��9��Yc�@`�I��?�v6�37�L��y�E�������K�!4p� ���p����ׅ��qi��,b2\\K�nC�ix��
mb�'m�D3,��Y^'���wR;b:�D4 |����)�BO��.j��O@�؈%��lR�����9��'��A} %x�@a����A����*[��C��
t_�K1��h�5��P��Ea®�DT�Q���7N5��d��2�]��^��96^�jW+���'-:��U�8��I\G������jB"'P��ލ�@0U��7�S�{�}�CxB�; j����m�X�$�O��W��w�WI�Ń��^r�:��߲����� ����#6�(tfǊ�>�P0?��(p:i?^�LR��j�JRX�O��K�D�R�N��G��<W���)��G��Lo�����7��9�5��?BGN�_�'��K��Q"o�'Lܘ����7B���H�*��J2	$�pQJ$�O8Gm��^_�U�25��z�:yݖ+��j�^;�&�/M���c�i�E#�;嫷Uy�L�փ�����Gn,��)s%b���C�4�EJ���/�q�-��S��Il{�P�No���>��V�\�O��*�c<R���C��]�����}�_� �^V)s;�:M�lq9!��w�!C�մXǾ_+{�WaK`jǵ��nU�$��2����FX�7�No9"Ď�7������aƊ����L0m�)��th[=
���E/���j��"��,��藳#M4�ڜد��&��	�Q���7���3>��8�M�oi���|���'p�փ�m��C�O(kX��ۦ���6m�R�1�K�P/A]r�F�>���6xPrLefզCG�����2����)؜6��ћ?�M�L
:P���T�����>�=�,�;�n:UR��aU�-�e]�A�P�O���A�&{��JZ�p��?�X\|��������ܦV�eL����@��$�/���ټ����XHl�=	`��@�N+&9����g�MY���"z�]f%/�h/[J�֩� �٪��%G��JR�vȃKp��{�\^vK~�H�l�tY��$����U�:6�U��"��TAT�3Z�+�\�H�$3 j*K&̓Y_�t?��a��q3d^���52��4g�Ca����_��4kV���0��M�]:g��&^�Lkl�vt>���ϓ	�x^w�u�P=����Ʌd�~���������	��wRn�����XÆ��}{��4&�WMeWPӓb�Xb�,�K4�a�_V^�A̬����4C��W��&?[�KL=ٗ��ف,]����?kY =�=XCƳ�z�܈n�k1/�XNR�|:qަ��ܹa��a�F�Z�&/ S�+�r#P�8� G��nD%۪~�G�Qz�W F���p�(�c�z���G��z����˓��S�8*��f\�<����W�N�pۥ���p�cέ�C8��Ps0�8�o��?���n8�����cx�鬾��N�6�܆a�E�A�Ak7�	f۱���";qb6�a�J��e��^�]SF���O��|!�RK(���n2lü��Cm#у��k��;m��:Z;�z�Y݀��=��>��t�i���)����{���k��/yX�T r��	�������<��,*��0�S>�suac��M��t�%}��KXC���{��9yq�v����̈́�����Q/����¾�=!�L��������dA)"\���Z3p����®"���3!�����Ai��B;��+�ƍz}��<�G{����	�	����$��٬b���%f/��a�J��a﨣�x��Ę&��cw�K�bk!�!i�KQM�B��t�;�q���y�D���W�Pj,EW��S���1tƄ*e�p�jy� ����e5����,�hn����P\��\AJ9���<�M(
��L��|k!W����E�O��P�z��p�!ܰ�9�yml�$� A�M�0{z�i\�s���di0dxx�<ɗ����.�W~�9g �8F��<��"_(C.`S��폤ҧ����~��ً{��J��,Ep��2���_�V4����G�\����Z�U����4B�*<h�#j��O/��/U��kSI����8�sJ���p�jz+�f&�����O��vh�B���I��v6�φc�]�'��Z�A[h/�����%Ƨ�����q�:n�%�w��J^��Iֆ���^�%��2�	�}���ϵ�eq%���[}v�d��c$Y�u�E�c�P�8���i�v���E�5:��4�C�}�QP;?]�"v�y6��/����}��t����E\�h�9
�:��D/)u4'-�\�
��
y����[A�Հ�n;_n\�8S'h�5����b����`��%�KU�X���j�gq�Q����].q&������ڗ��BZ(���퀵[�7>�E~�o��,4@f/�=,*st��/�L.s�1y��+?���(�da��`d�F|ws�!.�Q��2Y3�h#ܥ�����ɿ�U]7��jE^(�}9�ԯ���E�'��{KM�FX�"�S'�`��iK��G��S�h��g��x@	�x��NI=7��ڄ*��L�t��l�c��f�$/ͦ}ym���}��%�Y�֮����^3(¨+�hܷJIѤ��b��_)QW�U|�N�5��%������'ڠy=�d�z�^W|E�]���	�S&A��9�}�qBm]g5�^q��i=�q��z�O�y�H5�c�m��	�t�1R�"��ֈ6�=��/j����z���n�뮱$��OxJ�u�o�����Nn���ォ{?6,/ P?�'9jzFw��}[���^F̘���[��]��}tk�,��'�+�ﰷ
:�Q2
��{-8W��]鈸(a�wye��v�T=�n��ϙH�%�,:��H"��
�m��p?s�����}��^�Y�.�ണȪKk�:����Z�@~���̳̓�㉳9��_�,����m�dm�.�x��=��I�uMe�e�Өu�-;�<
��ߢ�c���: ���y�p|�	n(c6`��VkPЫ��ҹ��"'c�P�����]�����{���yߔw�ă�XC�Y3j�!a��M���<ݎg�l�^�G*N(;q��5f���#�:☉\�x�
cD���#�Z�W#���fc���rUs�ƭ�y�Z��.�i����f���t����Yf���m6dBz	��q��������(F����O�y֢�d"t2j.%�"�e�z.����J��c��&��i����X�p5�����y/�8��~��f},��9�>*)}���;M�)1�z9��Ecl�O��[��*�N{�]��k.�O�ҕ�BOPzxI�b^�^��j��YA�i���LS�#����ӷg�VĽ�?F��r��F���X<���,�v>�A�E��;�ǔ���};Ūp��]������pd�nc?�@����{3��gSO05Q�<#���^����Gܯ q'Y��#Mro��ƣ������M.�h��xe���}ڞ��?����G�N��33R(�yn,����ɒ`���2�^�˄nC+Դ,�>�hd��AhV�Y3��E��
����y�ݰ�b��E����8�Z�_I��μO�[�o�u��8���v�-�H涑y���T����gA5`EO�}���vf����e��B�Ϝ��r�I!� v*���[�I���������|7g�^��[nfrSk���Y���;��#��$#��1�
K�)��Mw���t'#<�%U5��V(|H��;�Z�>��S	�F�Z@*�%��F�0)0o��n���b�����bv
��n�����9Vjh4��:&(U�8�z�\�Q��)5j�i}�[8M@���P��gi�Dd.m�����嘽���R�����Jj�d���ݎ����1�>J������ xqaAPO]Q��FE�I��
g�c���͇O&c,幊��D���N� k�9X:Sm=�<��]���s���X�~7�j3��$�����Y����_z��Z+�D��_�)he��^��O70����D�	vRx|y,���`%Ű�l��+��|���_m�w�I��DӂO>�O�P���c<���T]�t��c�|Z����Jwc6���X������WI�@��2��}Y���q� ������hn<|�+r�:��@w��)������2(�ܜ��i�@�7ͯ=�(O��~�W�+kr�o��Ex-�q��7xU|u�C�����cP�:nm2"m�=���:��a CU�r�7���PF'���I�]��V1�5�fr��}���t\3���K���'�
Ir��/&E��TdMvnj.��np�	:5囂\����à2���!5�����Ȼ�6�Sv_wY]�2��9e��@�m����쮖�!�ϑZ�����â��+�vK�ż
�Z�J�[+��m����F��V�P,���5�����u��-��T���)�y?	�X�Þ,��2g}�J�Ò��h9�/T�硎q�h[��5���=ں�޲86�I��0Z�|齂2�q�L	�3t�؝�>�j�[�+W�Q��5 �E���f�)���w߁eF��Ea����M7��X4�ĉ�J/'�5�N!�R�R0���ƺ��575a���-uM����#��(K�Y/��Q~ɖ%�T�2��M�X�jk������&���RX�>�1�� ��|�V0��'���ZЁq�Z���0��
5C���� ��a�r2��������X���C3q,�'h�X�F�(1��8�7)���v���F+cj�W&�:����T��� �h�Uᥙ%����A��M�*����?��,��Z�ܳ!9s�y!��r[��wڭ]�b��R2B�4@�&V#�������<7}଩��Ϯ�\]u�/�/¹r��U�e�\f$
~�Iu�%�-�zm� ��np�t�b��\@mc�����J�K�8�5�/�ohO/>�Z;h�^7l��0C��j<��̀L�ʯ���t��J�z0vǬ���H��s�X����!\,[��$�p��t�������s�v
.-�=O��+��b�H)�]�
��9�G�'mӲ�sY|s�S͢]��d����9՝�v�6��	�fؾ��6� (����o�h�	�$���C:��mFͥ	��V�����no��[���&%G�l�7��>���xv�MKDi� ��<��� �t��&I�*a���U��g��A��w ��zŗP���CV�&���6ľ5�çL��4ωj�*	����%��(�R��)��;��P�r���M��9�r��y�!�Am%2����\��h� �A���a�����y���h��tJ^�׉&{�\N����{Y���ro\���R��l�)��l���2@��sg
F%Y�@k;��	�;j�{�ƒ��������/J��!��LeOmb̻���Pq��4QUtOY��O���`@��my"ys7q�p٘��/[W�c]�^p]&�3�G:�7ݦ��&k B�~����"�X�HX�_*=��޴��Gk�f��ˏ�j���L�^ ���l�\8/�V�_��K�%q��6�~7o�&�B� =�m�N푡j���Ң^u����M�.�T�����O���r�6w���>L��uo�u���Y^�i��@�O2@{	|��j�f\,_UN���|G��7�=��g/������z�Dr�?$��h����!�*8n�U�ó�ph�F���=q."��,.���hb!�g59Z�˰'��Ð{PA�b�I
	H�)\��s��#�a���MB�.��/��9��]
+�|������ĘR�V,,�ʧr~.9kx_�I9\�t���p�D�S�Z0��#��X'��l�e�5��C�<Dr�M�](FL��kc2t~ �U�}69���tk8��!�Nz�w�U�m,�w�=Fڰ�~�<�&˟��Z�SկY`c��9�����y����但W��q<I�E�Q��<e:�c'��๠��� �����_V�ʕgq;:(�9���pCH�i�|pO�������z�ɿ%=�x-Жh����T��&յ�5v��q
��������x���5,�����~�o�~�<.aՙXR�|W�u|�ޕe�h`� Q���Ⱥ �Ki.Ϥ�!ֳwƒ�R �|�_�e8���Iuc��{L�.��Xy�¬���*l!�W��bW²4�d��K����Q�)���bӲ�����z�?c*�>Lc��� ���XM�N���q0>/n�Q��<%�tW35_�Ido���������y��X6%0��sI�	ƥF�����ԟĦY�0�)��������,z���d���Ok�j�֜���wL_c��{��Ĺ�2m��::���2k�s��V�Օ �/��OM�����`y (�I*ߜAu��QA��;�i�!��B������Q?��s$��� ձ��B6����F�+np��Xވ�*�Se� �:��Җ�H�ou���amn	 g�c���kuIb��pST��#�f�ՙ��Gc��z""o؆r(�����#I9�5�m<�u5�HA�3X�+c{�{���x�rg�#��Y\�6|����-.hxϣ&wUO%��P��MeZ�gI���CE��#��3v���]��8V�X�3-�v���l����;`@��>�/,�'+�+ט��	(Ͽ*�L�I��5Qy��{а|T��U'
�-�@3�t �����(�7@$
2��K@�e��N�s{x�ރ�����t�x^�`y
�I����� ���5�v��[��W���I��bX�0L�&����������aF����x��O�eޏ��o���q�d'5֙Y�g�����	�ߤ�m� Hzo���ue٤�OMy���2��*xK9��j���_�(H�w�������2�d����M?]�A��ԓD8���R���S�`F]٬TB-}�U�I:>Ҷmk�T���a��}��΍
2�U*�w�-���j+�T��
A]�1qD� ��R\Mc���ȯ-K\�[X���%�˼�mxO��R��C���})�F�����
�d�L�ב�8�fj�4�]g���V���{�A�26`W�-k�h�C7����n��7ܿ+��Gt�cVk9wG��':N���Q}pNWT[�4k�U���ݠ���w�/jM�����h�Y�N$��W�!ю[V�s�z���7:!�1���~$������= q��qej��d��zs�.�x)S�[�_˵�/M�r���9J��'��LS���Y������7-�S@j��7��D)4��@�Es��NQRL��&V��(������G^��j�T~��g���>z�_�U^��Kb�*��Q����P��u�A"F}�;�����Y�R��G��0��]��s�w����Ȍ4z�N�-Y���%Z ��G�I����6E;X��56�Yy! �5����������H2	��ܩ��� ��5@�1R��H����9@azo��ڲ/�P�!VJ��آ��'S��7C�>]{@|U��]�2��ߕ��1�����	m�$��)�:���3�~������m��6X��I.�d��9hj*vz��]�_�Q
����ԏ�6"ӈ ����;���_�JΡ��H���۲Pꭠ�`��R�Ik�jW��X%���ޖv����`C,��o�>p��cz��E.b��
 �H(��G+�0x���p�M��L!:�ѷ�s�Zz�<�o�o�>�FY(�����0V������'\)�	���"#��9��:J�%H�g��QtUf$�&�\�V��5�"͕��y-��E�*��df��f�"tdcgW�J�.�\�7���K��n���I�'A%�P�vL��H	�`w�a13�.��g3XI1�����-�\#�Ӑ2i� �L�E�u4�&̙yG�ӽ��Ƕ�P��IA�*j��{G凌a0<�HQ�N$f���F�OqB�ɖ��v1���U�5&>�p�i��SřM?����8����8\���rƽ֥�yl��o�q�Q���y�����	(�Gj�z��%\AG�{���]z�)�o*���+0��>.W�%Ua M�p����y��2^�Na���
��b�����%c���?/s��SQ��>�׭//oHhAύgk��U���X=���n��o)z���S��*I���;d颿��MY�jj�sTj���	�ZX �E��<nu���w�]s�w�E/[dc�5	n��	"|�IX'Ӆ��?Y$m����I�bg�<e�w�<<�JRQİd;�n&F���hq-��)�s�D/�.��=��~/�Eg�ٽ�R��AB�}�xf>2Z���v��<�5��|st?S���T4��,Lvk.8���-����u�hι��BG��:�5��]kF�r���?����+T����\8Oz����!���w���>^tZ2� C'�d� ��b�c[!��Y�FB�����k��:;��B�1}q�;uA򃟦������0zJ1�1�|XP�#���+�4"�s�*�"*�gAg	��G�`3��?"�Iي3晉��ij~�3��J�N�7�(�I��dQ}�GqF b��������Q2�N�t5v��k����15�5O�)#h����������������d����/}�W��ŝm�WjO�!um�2�`y��V��S]ũx��H&�=

��Mo�ʿ J���y��؁�)�+q�͎�Y�X�Q0��I,���eW�=�N�����E�٥Kkx�~$J�V䲙4�����9oN���f�K�HJ$�o�ӽv�?`�rv�f�-'��|q�~����=�֭[�΋�+?޷�R���w�K��a>S!`��)�b�_Q���E�&'"���?ݫ}�i^�E��3ur���Vc��To:��OA��������5\�N3��)���$j�5��-1T���]�Y/�%��B��F�V��U�I(�.`ڳ.��-"�1ۈ��;~���K�8.}D�?��"�JQ��_7^�L�����}���'kCh��SM�g�!P�ҽ�O�$��E���� R�5s�W���4Ƒq����/Y��.M����*�@�޶�@�5V앢-m5?DrU�����?���0[Ʌ�hxf*��+.���ǋv&�[<<�K�A6k��b���{,����r]0��*$�&HT~g%dVMF�4�UP��j~�A�<A)R;�i�DV�8f��������Pч{W!}�yc�g�ˀw���Q�Һ���O�F����1���X6cWd���j��V0���A��߃�Q(�A�|J�U�$�3�[
]ğ��Gv�v�o�Ǥ%ü��+Z�d�Y^��|š���1-���������s�6i8?�Y��[e��Fө���o�;��i'�0�YM�0��f~3�B�olt<޼���%xlSaU�<003����c���!�愭�% IB�̡w��AF���/�M����/dFZo�J�
��C�� U\)�r^�N�o�Mӳ��l
�p{�ݛ��f�E���(?<�[�>�w7r�GWV�F(�+�R�ğ��#&1ˣ�00*��@.x�`a���y����<��:U��,s����2x��l7���r���I�1Ѓ�Z��;蛆b�2�A���@����%8��BU3��.,Ej�^�����tdx-��?�W��<�o��������JLX������9 P�=�"����{�<JB�e��K��-���"�X�>ޫ��K�]Ylh�JҀ���*f��{���
��:GSLVB�%f��\M�O�q���z)I��&�\8���f��r��M���_��  "�_���3��,�$�|K}	}�*	�y��;�&�>���8�2�[�pB�m����[�����M������o����wV�I�G5��6S�>�cȰIh?cw3�tA�e�S�s�{?t����`K������`��w#�n�ZMJ�4Z|����
級JC,��G�f)~�p��o����	T�^!}���o�̐���6F�+;�Ų�Y'9RbI����U�lE,�9��TRX:e��G��B5�<i����l��+� �<���=�����l�����ƣ�F2�WT�\#ewAE>V@>Bf��%�/���]�A<U�Jܩό���������N�:V�F\�ϼ#I_��'���!
��0b�����}�1��p����G��0�+<��VV�X��]��<l���b�"h�0?�'���	?v����vBP���LH���x+�OY4,"��FT�;��P��L!p<�gF^a�x\�8?ڥ&6j��lJ�vD4z,������~�Y]�#��Yn�EtA�	�2"4$����FA�eq	���	��f�m4�@[לE5O�'SJ5g�0���l30(�q�e���J�w�*�����g%-K7��5^Ý�Ӏ�*Z�I�'Y�^���^�`�	ς��;<DWy����_���HQ<a�l[�h�	!�R[��v:�U�?L��ӨI��k���̀��?���z�zG��щ��u�R�r�7
<#�t�SO�3\�N�7����N�}����A� u<^�o�TW��Ж�뷶���(�����4�������<��B�[Ӱ�{��/��2�u�{�Thek�HY��U��h��R�x��q�*}�"Q�|�A�'�y��4^ M'�8��6u��do,Z�lKY��"Ϡ>�4P4�
�AN�4������
�d�Mv��%$F̂��Μ�-�Eږ`���U ��,I���9ʈ���sq�B��N��C��݁V�41��G%���'i�=�h�#�cA�&�1LBnܫ:!]�<12M|��A�f�qG0*|�y��;1~A��8�^c����i�%##�0��؛���ݡ,r/�� +�h7>	4������b����ZUT��&���'`h�Wf6C���$v�r���ޯ��"��M�F�H�s+�@b�3g���5�2�g��n��\��n��$~���z�eV^����+�I7�[٫�i�jê��E]G���Rw͎���R�R�\k��,$կÝҳr�2�\�KN�s��>���h�yN�jE��ϋ�Q��e>�\��(4�I[5tυ��5 ����[��"
mb_��gJ��C"�i��$�,*�}T#�@�z���2=��`�\R��ҼC%qft�P��U����:Y�N}O�o醷íx-�4w�D����U蚻���Q	5Ł��I9��$����q���X��3�r��e��[G CP�iH���}�*i.1����,�=��V�]7�e�#���6�: UpG�6p�jȆ��������Btlݫ{��^~?��[���h���:�肶΅���]�"^e��h,?��x@��l���d��k��Ւ>�琶���@j����0��>� ��+W�;�n𥠈��[R�a� �4� q�p]w{:��5��+�+������y��~�~�zeA}���Y|!�J;��(�M��=3�&�ӱcG���e5���$8}E7���9�X�Nc\�HYк!H����ŗ�t��S�i������Sq��������E#rE�/�[A6>a��`��ҩ@c*�p���À<:�ƚY���%��]jˋ�6Ǘj����S��@�w��6F�l?��c�	�+dE��]u��E��-�m����TQ����zK�ke��hN\�΅Q����^b�Jb����m�#7a�H�4�Fj�F��'aK.1RE(E�'�i��$@̿�<�;,C�M=�����]Bs���{#���'fP�����
bt�%�%�?M�i�|�v���lFw�8�8�(��z莳K{�^�b�*��rn/�޲{��	���?�F_.�RɿR�����vt��(:�hz��f�Y$���)�W��]_��M��Bgӂ��$�zS�i��Q��#2������F�~� oᱍ��~W�!��b���{�]��q�s��,��
G���t>�)�.��呾���.�����q�/����ׯs��1�3"����x�0��,�� ����&{�6�x���@�Z6�P��k��?%ɵ���|�4l-i6k;�����k���سsn��+��SFǜ��ݮڇ{��%[��9�%;��ň�يxOl3
a�MW슖���y�K}6:x����|�s2"�^����b�_�m�/����h缪��|��/ꤦ��������)����&��i�L�,������VI:��u�v.��z���p���up��l�jJEѨH� �J>���ܤ@���>�V��L�ဟ|[�z��f��Bc���Z\� �f�$�Z#� ۀY��Xti�2wȼ�Hw��ì4�ɡ[L{Tm�?��,�jtsC���������L����<��q���US�v�f�`��M��S	tYW���U:��N��{�|{�M���a���+dm�k��Ζ���)�,E6����k��FQ=(jO��Ǉ���\��xM.��[��r���k��K�����eF��A�f,�{��&u�TY^N�J���dy.it8M��Am��OoF������>jB~'�bHy�O��^�|�(dA8yK;ng��{53��\���`���$�
M�!I��_�~mre�Y�~�I��2��^�a�7��y���R�r��j]̛Ђ��x�����MI���BM��~jE��#�:R���jgav����"����~:`�wpa�2ܮ�Jp��1���,yp!��#���������M������+p��݅b�X��y&�9.6|�#�
s���
�H���ˁz�})����6�e@��$���m"�n��T�V:�v������_��WT7)���r@Zm�nZN��o�j`��4�[�&�(�l�}T������ZD1�c�ќ����n�,+���������+y�cj!�6�V�\�j��oS�/34�aK*�M���h����s{mCz	���b�n1�g��M���@�����s�"n�SM��U�I�h���{�J���i3����Ys��,bE3���: �}�*M��~۠MM�Wm77��/4s�W��~�x|�;���N���1�\�k_&HK�� A�>��I��׆�/���O�b��'|tr�9�7��y����E<��#4�6T�,���������c�K�����)�)�Ո�V�s�6U" �
5%H�;��Z����u�����eǈF�J�}BpxQJ��	�%:f����蓒2�Z����y�_*���g���[o���4*mz�=�鯛�]��X^*bo��V�El��f�MU���b�u�t�s�
���͟��X�� ��X&�yrU�(�pǾ��DШbFz�)�m��Cm
��Slt�n��4����D~�7��m+ n�&��g�m�:Pu4�d�����٤m�,�q����q��ބC��F���U��򛼳올'��e�<��&`����ciRN�-��`��o�����Cݤ�k�/]a�D=��"���J�Z�׮pg�]ç���yQ�N��g��TR�� �8�J�p��_�B��q$7�V�l7��������3H2�qv�nI��t��߂Ǒ8/ǁ���;��/�L����8
Yi���� �S
�)�v�up�Mcwj�T�X��t���%����>Y9o �3�3O�}�r�+�o�s���tcЍ1Z���BԖ��t�B�v6gЭu}N�0BEr/�Hc�<&+����lY(��+N�7���H�M������SPmoL�}�a��)���G�k�u/j62�o[�����6f!�p�v���T� �z*w��D��Z���L��SޟO�
�GC��W�<��kBg�jf���⇹/Lե�����i�<�*ui=
t���^2�b" ��j���=���"�=��-(�*���|X�cf�g��sT�����R�OQ0:%n
q�V�ժ;���:X7�"Hi�o��@Q��\ٹ�z�;j.�I,�ZF��Ov\��k��1'2{M1�Ȏx��?D�ڏ<��� =g�-��
O����(�Y�;�g�ݲ�����'�.��uY�`~�\��3ҡ,?��࿩]1�����$m���	zm7#�mu��kf��ᄮ��Vik�j��0R2l2���ޤ��A�~�Sq�߹rM��J�|,vWX��s�[�#�<�1���8���b�U5���C)a���.
;a�rjh��(�����"� _Q)�P]���Ӽ�(1��+3~>��g/������^�W�Ҕ����X��hz�a�2� ��:$�-w��DZ�y
��G��\G��S��5���l!LT��`F�%6���|=�x��}�xM�� ��8fL��s{�_A6[E2]q�JH��%�Ӹ��ӵ�s�W���١������o𱶈�崑�`�C��\.M��o�fX`����B���M�Ҵ��&)�E>"ܙAc<���^���	��z����/�f,��ME@�����-9Cn�3|�oiI�����Ӷ'�|��w��j�,C�zμP�Y�͍`}&�z��]Ύ��8��d��n�ơ����e�w��.#�b��=@��pbj"��D�Y��u�ٺ��n��zsܖ� {ku7x|A�J��d,��0��	��}j���C�gȜ'f����{ܻ	��F�����QX8ӏ,DBiB�CNI���(1E���?���5�nE�$��DG��{�P~U�u#����<g�v��;=���2z��jZ/}	���8�j*L�w�9���q����*6�әԱ���d�8e��Q�P�Ԇ�@��ܐ;�*jfV̽D�{3�s��z��P�����_����&o��*�Ez�����A17�7b��6p�1��Up�����M������y��r�����}�?�>��R�,�������QgC52���NY�R��e�V�!�ݠm�$��
�~�6YY� ��|�-ì�-A���U�-��_���7M� �ؼ8����7���C^R=Ny$�k�YO�i�
��G������iB�z�Mj���Ĥ�t#on��I?�*�;�1�)��z���c�T�s�`�t��32$ �l.����CV����[��vcmZȆ�Qgv����"/N��O:�.�����FR`$֋St~ʣ7G񁽃Fa�1Gs�4F�L�Y}"t�+	�N?U@a]]1;�?{k���!�b���˨���-�,��Ŵ$�mP���]�PX�9U�<,�1��mL�B;��<qE��k��j�����j-��U�w�jBUZ{���p��WC��\~SM�]�O.d�^`�"�qV�kk���f�Hq��!��g�JTi��+g�w�f��txR��SWl��GV)e^V�\{���.Vԓ�O��
DM��^��C{���ːY��w��alX3�	G��-.<;��)���&�E�#���)��\Ȳ���d�Y׍ �R�U�13�+]bCx�&c 3hJ��H7w4�;�Z�@~GgQ� ��AG��:�W���'���ޅ���P�R�'����/V�lfލ���cf�=���P�-�K�>�@����;���_C3����!����F�g��F������p1{+��Ȗ�K�f��B��<DJ*Jk:��|��`������������IK�LP��.BCHPW�;�<��n����r�����Z1�EOR"�ȹ��xl� k��τN�Z�������e �"7M>�����A��;�[o���0�R�S��C�`W�$g��^D<~&bB�A�F)˟�������������2Ce$�� *&_�iZ��ϸ�ҋ6	��h�Rg�@n���>="���XU�V/����9;�*od�#�WCUx���t�� :Se8HD��V��ꁠ��5`4%2� �*��+�_�	�z�?��8��UY֊Qe*Ȁ)��Z���a�U6��o]�	`׃XP��u��E�)��EX�ʈ�C�)*f�`��0/��q>�5%w�F��݃����Zn�v�<����77U��6����b�)�������ġ]��(nQS�E-�A�zy�9}gN��mM�7%�Ĥ&��¤��_�9��cc��<FP��h�u�&�U��Zi�r?�J@��k�s'&ֲ�{�r�J)ݐ��w�_��<�R���{��Q�u��R�Ꟙn+Ȱ���Y�33���K�&�gD3g yH�r���L�v��N��&h0c�X��7@3��3@;h��������R,�����d7{>�jm ����:��MnXƳ>[C����y���7mo���	����Y򴧽=ڡ��5�������Y+���ӾҲ$�u���^3����'�jG�� �l��P@ȯuB�LuvLk��s��U��5Lk����'�\r�;u�x�തh��<g.�����q����BeF�0��4���=(��B�/�D�cc��z:\�kp�:/a�
���9ğ�d�Vo6l���|�1�2�uI/��4�W���`GAw�Qyk3�))���C�xA'
4��>&����B�{��K�B��x�����÷������V�ҍ��B��Mg����wBB�jG�'����[R��X� 9�S-qt���% `�1c�ߚ���Z[C��[=��i%�17�:9���I�vl��a��� �$)�1.'g��)%�K�<�5Q��d`W������4QJ|���g˟66:j=�	�v�z�#��i�;���������{�4��ӝNV���^ "�.��Pu�䖇�8�U�R31eB7��>�����82jgnT@�x૞�cWz�V1�9����:��?���R��Y7�|���8J��K���n����_AN�,>�.�p[�G*�7��E���:5`�sџЅ�^�ܞ��)�*���׏տ|�Hm܊"Ŭ�j?*k��1w��G���z���:�?q'>Zn�w.�o������`���w����r��Tr��{�g������EYl�[�	�v��e���d����9���u��a�WV	�� ��4�^^�@��5vɟ�	qT�37_��k�7��@g�$ϰ�n</k�I��X���]���`5���b�0�X>�}����zs}��̵
��1��}m��\��V��д�;���̂���x��
�?���2j���ov���J�@����b�Nm%�o��U恩�H�MI��O�쬒��z�o'9]���v˝����x��=D�Z�����Ǐ��w�_�R��,��^����g��zk��~Q%Z�m�~Y���j��d֏Y((��9��k�6��M�>:��	������FZE{i0��}n���a�?8��MZ(s�d���yǂe�o��M\�%6�rx���V���z�7P"�@8��S,��a?�jer �:�+�Q,�lR���:&���Q�Xѧ?�6� �e��<p�Z��-�!�~�v�����ƞ�afdߴW��5�e�	c|I�O��z�� rdiD�}��6��Ty�N0'������"Omյ�(�۵���/"��G�G�����IN�Z��lX!�D[H�/���PcOo{��+|��lۛ������b�!���ތ23(��;�~���mx���r�Αt�>�e<}�yU��O�g���.�g��sF/��rSy#5�9�;6-O>�Q0�9D�>���õ�a��� �E;����^�c��9_y�l0��Qqދ樫�.�h��Q1(�n������E�i/�G��A�i�ⵢxN�?1��n	G��7��P@���һi������ԋ ����*լ���+�H�ئVP��<��'������%O�;6W��bF�.ڝ5w�Vx�Lo���By���{�5�Td�����������!w�#?H+���Z�"G�5#+�|(�B����=�0�BYM�p�q��w�t� &E�Zw�+di���jE���������0Z-�Q��jL�fL�����ʷ�ڮi���K� �a��\�#�<Ǣ<�'����Ɲ�$�^�o�#�!��G��qK���S��b�iN��	�ӕ��FXuoN��J_�~S�B.�}Ϻǣ�J#��.�3|&K�W/+=��KK�	��z�;� ka�l�Q�J�k=�+��S�#W!y�г%4E#/��j���fWA+���~ZP�'0��f����`����fH���ľ<z��'�1�y�V�-��JV�{=d97��*� ā���?&�)ѝ&�Xr��6���	�^N��H��L�f��>��f����(�e��`zE��J��~�V���Q���ܛ�?q�qsI��0�J:����k��[crCj��>߁}D�ZZ�Ԃ#^�m����C��ƣ�퍅?�:�j���M��IQ����#�Or�ȧу��;3��5Z�쀚T8���,]� ��f|���t���0F���)T�<E�:�T�!:���@vKKY����������<�`/P�G���c5c��8E+b�h�X#~^�e�s���B]3���/�&=xdyzO@
�����@�yH{�E)��M��ܰs�@z�0�^G7�O�@��gqgi���_:K�5�::��� �{�����=T�N�7����\g��#O�в��D(z󗓠�NW�fBt�6uLc�R8�65������:[�Ȼ�	��Hq��|F{d�x_Z ]%�� /ÞH/�v%��c�c��M	<N����U�,?Y�{y�Jĵ�/T�`͉��Z�����d�A��|�fFNً�Ʃ[{e�08��UA�΂z�k����S�&Q@PwYC��64-_����o�+"C6���5q�S��ٔ�������V�>�;D�9[�V�c,2]m�m
���q�97O���dwj�d�:`y��騕!46�3�u��j�Ơ,I�e�����w��J���,��\(O��J����u���r�b!��
�>dD3 ����֨�CH�OVa���|<���E�m%c+r0��c��U-P��c<��������'a���"�*����O�g! �@U�p��	�P�������T�O�̼���Fo�q�*��_8|��Ñ�"#���L����7A��W�+�������D(혓{��3#olv���qH�<��n�N�l
�&p��X��8�u&���g��!���v�Կ �弣q���� �}���i�yC6K�Q�T_T���k2h�"�G��w������"4=�c�n�@�܂�|��=j�'��3�Y�a}ڧ�&���v�`��H�(�������g=/���Խ�k���6� A>=,�Zɬ�]���޸P���"�f `�ޔ!LD���Ȣ'z�,pt��k�)n�z�"��p2�. B'��T7zT,� ��;�H�Q��Q�_����D���̄�S���^@�����f��LO�ג0V0MI�7C �{
]��9��К8J|j�n��DX���/���"��>�~v�,Y��9#�#�#f/|[?�t/�U�,�>Ub<+����2��>M�갟�!��;����Gnw�P�/�ϴi�����'5�lM�>�J?q��D�ļ�$��,���u�N��p0�kdD�Z��uO%�ƍm�cn��@j�C� �(O��a1P=���.��H}0�mhԤ���&{����D�a7z��Z��F�bNтfZ�q-0.(����S-�ry8�B�X�s{A����S��\__"/�L��Q���<@��Խͥ�~�A�3G6F��"? t�d
�p���'���.��e�`����HX2�ޔ��s��"�͞頛�\�^Z.6�C�������'<ڣ�gfAx2Ӭ��x�叨�r�9��kʨ%]�����8E��<�?��;��H�B�Q3��� �]�8���
�~�}5\U7���ϑw�錿�(4�	�m�4-��>�%&�gn >f��`p�}<�
��Bh�	*s�w/�u���f����m��[���Zwx�,8���Cx:��܆��0�6�*���X��f�Bp�!>�s�V��Wn�?��Y|}[dTY�%2P�%�Y�藯x!��9� ȳ�X6���҇����Jd_�c�e�}%rR yI 6o���G��;l��Y￷?I`���j�Q1}\��t6���<���R=X^�Nˏ�ГKjYQ_?b��D]��}��uy�6���=P���� 1��o>���뢘�{�/j�2�� ��f��
� dʿ����S]��9B��.�O�?Ӕ�D��ף�NC��(=(�0Z���]�Z�?C>U�i������h}ɷ�'�rl���qO}�`�4��|=nyee~�@��}r
U
̮�v [��>�p'����D܅qs��FN�ex����3�l׾�=*�b�z�>[Tԉqb�Ƈ���������֎�Rc���t�k�kBN��p�_�^���PX�8�P��G�.�M��.vt��|�qva���j/��F�=����ĵf�6�������u��u9�f��4�ks�����ֽޭi����3�&�y,�/�~�e����
�Ǎ)��v��}S�������l�H���l*�b_d�n����/G:�K&Ϧ��?u,������7��ǿa�)��~�	ѐ�� 6x�i!�I��3�vpC]B��["��(����:�G�f�'��������Qs_�3I�e�X����	ԕ`Md�~�t���;M/�Fщ3��V6.#�՝6��?�znv���E�7a���3c������4#�����!\���X�ٌ�%Ͽ13�n~?��<�a�va�a�m
�Z�W��`Ж?�Wۓئ;�퐨��䖲a�7������9�=���MϡN�J�q��xQ�޻gς�����棒-��H�g>�o^i�ݓ��Qr۾�	[���$�v^��TiV��c_�/��!�cihF	��8�FB)�r��� r�J�� v-P�jf�"�߼��X���d=W��\����U��W���A��[: U%I��/i}-qߛ�}>��p��l��l!9�+�d�R�R��<��!�X4�R��E��y�J� _�q9����PŰ�g��5���SN�1my�q�3/&���Dh���/��҉$���i�',�*�U�E�����[�t�91��6�qd/�&w�v{���I�A�H�<�Il�]�t��3�Z�,ڟ��ܓ��`���}�ub?�W�pr����b��Y��i�	Uey��S ~ �Ϭiz��,o�R�QA�չG4퍔���ofX�}�b�Οy�X�<;��q�Bw1�A󵶗���|~���}@� �Z9���b�T�Q|����g.ź��0b�Gt�#irr�g�p�q�8�]��I�ǥ�iǺ@B��?<��_���
d!R71TW����{��(L�vO"%~�|5��5�GL����EV��9��&�:^�ʌo##wn�����s1�=�v�|�D��i��u _���T��.��dQ�)C����׷{�U�}��C��i����H[~5 �&�>��&e�#�R��V�I������韘uڶd ���ds��7v�S�Vr��*�w��	���ر�[����y��80��gA�d�.���$�|}�Yc�I�hf�����P�n<ɷ
f 9iV��S�b|�4��3��,s�b�k��6������v$��'�5��g�b�� �F#�D#���'_����6օ����~*�l�O��p^��$���7Ȉ�BiX���H�J!"�GV%S��|����۪���Q7;z�rP�L�V/^<��QYmqK����aΞ�3A	g#�r�LE��s4���y���$�BX�L��T�r���`&m��+���A)���fG�b���"o(���뎿o[(� �{�	v�FSL0&g<sa�8C�\O���R����۶�e}�	ȹ��Ey���|kᯃ���Z�+�?����.juH��&x�|���O'ђgc����yT!α��d��CO�3����Ab�����je�|�X�a��x㔨�R�M�'�A����C[ji��P=��j3�u��]�#�����p��Xƶ2AkL���q��Qthx�W��SA=�4-߁���1^ư�K��u�3�)˳�X�<c�7���j�k<lİ��p=n�Hnf��j��w`I��q�@!��~���1G�FW���!a����f�>�3�Ī�~��������q���\�Lt���hȽ�xH`	y�s&o@ >�`���s�)�k��<1�"p���i%�sw��N���e��i��Ǻ]��E ������7۠#�o���ꅒ��80��x�[	hN�6�rN��N!	��@�i[��e�ZR������[�\M�͈&��+��H���֧3t�&^JkŚ��Miݦ�l������0�2��ΓvE �n U]5�q�R8�0�֡u�i�Hc@����K�V�8�H��n���o>�	��/}��"@]۰���h=�'�*d�rW�g������]/�}~������6LPnV��87s���L*$��Qm��G���b���,���_�z��j���Sk����Uh��kg���xM`PV�̃���<]м��~�<1VJ	�s��5�O�p�󭄣�7���ɰa�g��*3��XsL�澁�zI���8hZ�@���7tn*
P�K�ƭ�h�aږҔσ�֥��N�x���V��q�Z�2������28��X�9���i���N	M���<ل����4n��YP'�~���" ��,/��W�֠��yR��0��ǔ_������ա4N�d��#�t�mj	�_�������v2�M.�Xs� ��	l;}�aZ$�of鳟�R�J ?��j�/�2g�� {��G���{Oy��>d�_l��s�Tܳ�&�֦��8<}�##	�KO�f��o �����
l��4f6��䈇?Ն������˟<�k�y�"	w�YC��l;���U`t�d��՟�;�׷��X�,X���4VD��\F��9�=����wc�X�)X���r}<J��+iI2��z7�˂+D�N)"����C^'^
�fd��#C�Y�J�,��-�^Ø��>�1�#��3jI^g�ʗ��~��g�V�A�@��j�?�o���rj��),�|A�`�\�Bv�����Fh�]÷���C����Tq4tc٥�*#/�.o���PKxO�-p�0��m7����2�{����ذ�|v��-S���6�L/?��U�Z��䃳�A���+}K��,c�w�k���5t�dT?I�^��X�j\Gs�T��������6�ǝSQ8-L4������TA&��Z�<�[��&�NW'V�,��%��bڂ��
�0�_ҹw�!t�6����e5�@ˠ�6�l6��M��"��4��&l�I~�w��C��ݼ�-P���kLwB�E�̭�k��e��-3Q��O��º�b�\2�0�Ƕ��?�)m�����x1��H��G wO���6��ūS��X{��(w�񧷥�v�/�O3=U=�*��E�!Cu�\XB�DL��;��=����;Z�$0~���0d1���߅U��@�[���N�Q�D�
�ףq�3�E���}>�bJ1��a���#��7�:�[�b�dc̰53.�{c�.�h��8:H�)ǵ�g��%TYz�>v�&��+%�q?����Y&A5�~�_ơ>��"NZXώ���Z�*<��46e�D�]�x4�e����j��OU���D�F�Ӛ���S����og{�qK�0�.Rg��SǴ���KY���]����a�\��CB���0-X�H��3�AؖTL�����	:?��Cn)�<a�w���;%���ħ�aḔ^"]h@�c��c?�_	h��M��~�'%�W���ᴁ!}���8�Eu�苑Q�?��B��r�c��j�� KV��_�9kO�D��):�W~��=@��c�]���C��:)��"#C�V�6��l}��������x��ޯ'�IM��4��p��(�4e��5��a���R�6�N��N�����T�6I����X��[K�F!s��������hy7��s�L���c.��R�fM��^�G4Okj�P�v�H�i��{N}ѻ�����aHv�����⸳� ���.0ڸ7<����ȑ��5>f�`D/�L
L��9xu	�,j���SRBQD6{f���e�?�q*>��<4��p�;8�4��2AR.֓���`)���"����O���n̷ ���G��v���˨�������m�݅p�{��o#@�Y��X���H�H�;;�h)7aىl�3W������|��1�~c�Q`�����ם&�|�f��ў�����b�V�UO�8k}�Pߓ�/d\��qrz�_�%�cd�0�s�z��J��j��j��B�>|e����Ƀ��NG%@�x�c�.�]�cs��]�/�b�Kz�����$�r�F5�:��k�]��lq�t�+aR��w��*�_�s-R�6ඏi����CPw�]8mu�P�������_�-�l��-3���^������
Z&�Sn\����mv��bH�5U���Z��r7������������2+:�Z���X�s��?!�{;!�a���Zkz��fɽ�j�G�Y�)oF�-V�V	���t���z��-��  ݈h?]��V�3��tVy�%F�-�L�`I��'�����x;?������D�T�&����&� >�$�zq��{��Ƣ���E���-����[���'�σ���)��&�pgN]W���BdS2�v��_sjp�r���jbӳb�Y��)y!f�����H,|��d.��Й�r+�3�6܅l����٪j���k.9P�[�}��o��R��o�[��t���̤�K���Z]%F �hX,��'5�qW��}�U������Q�!r��`�	}�G8���'�F2�N��- ?`Z9�O�\�J	>��.DK���ɰl�qgk�kd6>�F� ��@d]O�?���B�WFƓ�<2�}�q�rݵg����	i�\�-���Чܲ�b
��@AN�g��c@���Y!Q~����KŐv#!�_�B?5�~�ƩNʛw}fw�쐦�ڡ �#Ѕߓ��
;}f�g#2�$�Y{�j>�ì4������7�����}�]G�̼���Sr�ە;���b\3F��8�M5&����|P�]�k��L57�o�G�x�&��%&|�k�ЮD����̬Kn|����$��p��඼�8.���%��N�c_�9x���ٜ��V_J�����kv���˭q�����B�E_ZI���C'i�Ǧ�@H�?*�F�0��(��"��N��
Ό���q�����lV�j�֍7��;��#������4`X�6��T%��.?bk���z�r*�-��<�|)���	�#-��HQ�(���e���К��j�9:���j�B��"V0�����������[�5�ˠ>}����K����UY���-^c�q�St�t���?
4b�dI���8��!�ٱ��"�]��Q��z\LXuiC���V(u�*%Lʴ"}���;�X)�5йw�ey����?F5�����!�	{�/���ͻi��M��s(��H�+�����	G�O��3Ϩ����Z�S*˚+�	��L@'_5����rC'��$��zf��c����.�3$y�����0�zM \J��p�����a��m���>w�&Jrp"$"6+�Uw�;Ϛ&T*�:���?S�oNf�5���s���Kv,7.u�u3��V�w�NOk�_��H?Y^����|�>�*vv�jԏ�6��K����yA��F����N�Y
j�VcLtV�Z��]���s�>Z(#����g�K�)�T��GFk:]�%�w���6���L�ט�'R�T ä����up�V�q/۷�}�p�8�d �<�%�g^���~��n�$�"��jm.�$$XE�r���{<���r��D�>+^�7�/~4��^�ztl[1L�����;9��D¡GOLe^k�a՞���h�)�E]��L�s�uK�Hk�O���_�%a�餏B�/.������N'�d��ϝ�VӐ���W���C~Ѓ]W&�E�ψ��0�Q����h���o&�w}�l�{3nmk[��"�p}�:j�=|�{q{�@�!�!��kY��F���v�����5�G=�wrJF�zm�@���ɾ�&:����Ȓ�ÀLɐ;��w�IHk�C��p�U+O�rJ�Uh��]���BL"���L�Y&Z;c�!':iO�S��C[h���n�i��,�[�#��Y�~e�Ԧ�'R�wԾ<�VK��v�� ��G���ɫ2�O��a���1�o��^A���E�JÜ�ψ�� Z�֢�U����	ξ��U�q�i��<dD����x��f��.}�P�˖k���}q�E(v�z�X�[�<�#n�Z��zÌ��U ՕMm��J��5��]^��y���<+�/�����0�,�� >��m.�tp����B1������#�q&�t?��Y
��s?��cl�)w2��}o�Ϯ�j����:�i��|�)�G�.��Q�ku9�?B0�s��<�iL���\�.��A�F�R}7�v��OB���R������!^GsAMO�L��s�֨I�t���P�}ޔ4U�[)w���n�&�n`8�/����EZ#�iAȬq���pӆ�����ġ<�i�*tؾr���?���s.=S+���L���-�kc�d���R�J���6�%�S����|�n�]�7u�MǺZS�y�'2�ߏ�����s����م15ftYW��3��h��:aL65"�ɨv�7rq�J�����jTVw�o`B:�ũ��֝�"�y���E��J�:�p��&�c��8���]��&T����/R����������[,��|zs���(u��o�4� z�?����!�>�Z��<�]���v����d��#��8�a�-v��0���<y���C�B+�q��,}V�
�|��"�wi�þ�3�4gȬ���������s�k�ɩ��V�}���n.1���������||�&(&cK�'y ��s���Ŧ?����1�3e�
 �NS���|���q1��(M�������tޢ�BPĝYÛE��3�/�h?]r9��0�P��vz9-�#�
p$8n	��e��)��>�R�5��e>(RO����-�1pqe&Y�im��4ԥ��Sx�rT�J���o�wf~zP�cD<"�5����`�	����R��.�0ފ-D>	�˸*�5O���%m�,F��)�/�O.�&m�b]I�31ڕ�����p1�`�kmMվ1��x���C�`�Ӧ?�P��K�+��P�na!|P>��fq�XKP�C��:�m8o#<Mt�;�$4�J_��u �C(��l�ꂵ���0f���m"b�z<�h�Pһ����*��c�Dn����VT�y������5����q�l{�-:x�3�p����A��	z�7eQ�^��C�BZ��k<����5;�R��:��v'�*���������Bc�H���LQ/�{?�� "+���[*�q��D\
<3�_a��D7��e���X�%��L�?u���5��V�Є���N�Di���}��q����\=c��B*�{���.m`�P���&���BkFY�V
�t>�J:*������[�7�pW�/!�#����m��Sg���V��jlBU��#0�74�<���J�����.m���#bR��P����f��$��aOZGRˇux&T��d_o��2��?9���n��Z@�mKM�PX��~˿��:���xn/�S�O�% �*1k�;3\����P-��k�������欓�)�s�V�;\�n�%/:d���U��U.Ǖ+μ��b>�v`��ׁc�u�٧�5O��Q:�}7�&/F���W������O*�/�;�������7U�9��*5:��:�6�2t���L ���AW�9���*���yNI�{��8�P� G�l	�FZL�k0\�9o-���D�'S�L=�]Np��x��d��,�4ۺ�5"��?���B9���N����|����F�%���8�yy�r�X^�Kp�uOt?�:������~�YUa|r�Q��(=����[�3���#Z�m�}Gk��,�>�$��'�ʎTD�g98��N���u7h��ۇЕ�@��Ȩ:�:C�ӆe�A��B�ƶ���kv��@��������d�<�l��G%
�C�܉�hZv6�XٞH�%{����ѝ�؟�a 1�.]rM�d'"��,����z�Bb��gbX�_�EM,�S֓�f�4j��w E�AFH��#�z�H�t�V�����j���YCZ�TkŔ(>ݤ�|/8d����}��S�����_�V}L0���EíT��	��w��r{ۨzl�Jre,/�T..d��_4�ZN���_�'�~
nc\'3ϡyv\ϊ>��롐pG��fő>H�M���3N�t��f�7�|#�~�F&��@�k�@,����AF��X�̷;���ޙn���В�k���R�h�Vԕ�E����E q���"��å����rg:Y�d�R�[G�L=��[�+4F��0齴��繉�B
H�Hc" ʡ��̰�.I}��\%�  �=���1�$к��ei����X=镯�eOoa�C������vP�y�<z2VϬ[$�Y�6tXښ�-��ZL 1���CÙɒc�:�j�{4.����$�l�3Y^��L�����PT�F��(�������H���q{>����=rVW�V���En�o�|�v����*VM{ަB������Jɞ[�4i*JS?�SN�J��A*X �6Y��*�j�qq>���"�1x��m ����z;�!ϒ���a{��_���h�S���4*��iwp���;n�4��Ԇ�����H��ׇ��(���10�Qc٦�8#:�}S����_/j��m�����w���Û��k4Pϐ����6H��y���3=�y)^����u��r"5|4kDF��&�g�<E2 �I{��ϟy*~b��],�M����5]�֊p:T�'�4a(&��*�6"��A��r>JD�oC>5�Tj��=��#C��婰2.ލ��}L�Z��m����Uo<I���$�������Y���j>�^��#?��DT������{�mj�M���|oD�5�f&¶x��0��X��í7��d��L�<�-��-�O���~"\�k]"F�w��yX�8�G7���"��r�-�P���U��d���r�p�)p����)Ss�=�9��^�/i>�(�ƚ��<��'�;=�A3�7\�*ǯ/�T��䅻��x&o��r��"�-iWg�82.�1��0hU+�y���f�3P>�Z`X0��)"�>�S�˱��Bcp�^F���W�ǴiD�����i>o���d����5/�"�ul7zj����ViYQ"��ey���!2�	>zU#��-�%c� �,�% q��~1C���VlR�"rF�-KO�S�d�
��v�B`��������bGQTꉶZ���������4"���׸����`'^HT��	ԗP��-|��--�ew�A� ��־�.Y�'�#�$W�$��-�eKNs�4�GPGL��[jq��/�Rx�:Uf��?�@�6OK<�������}��B�����Flc�0�EK�KJ!r����N�lg&%�2���˔IH�����%���3�Z1k_��d������ѥ#!K���}�r`�>M�V�M��/)���S�0|��u���{�؍�ބ�gbH��U��)g����{;)3d��L�Y�FT�E��u
��ȄT�q��u�y%� |�|7S���'�T��L9M?6��6���ԓ�:�t _2nc�J�}�S�n{�֫1���8���0v�O8�ɣ`��lwuT�u�LolH��%Uh�Z<�T!�ck,��\�?i��x�%��߭1S.���H���U��DV�:�{���j�~�@��Zh�,���!E%��y�}�9�}����";���	ޠt���~�[��m��
zL��8t �	n�X����6���9n�W��_�p�g���&uSK�	�I���-o�-�S�U'�*�����UI���9$s{�rz䁐�m1�B���4�Dú~�]����&�+6�,t��`	��,,��2-���4�zjɘP��\*89�r^G�[P(j]оj�_�)�'1� ����	���T]�d1o�Nn@!Xby7��u��ku�H"��`%���a6�b��-%�R
m��3Pq����h�=����9l�C�n�<ɑyŜ��o����"U�e����X���Cٍ���k)�JB�}0��iX	�����đ���!�4Oi0��[߇��
	2���A ^ ���gsp�9� y���B��Q֫�5ۯ�]t+��IS��*NJJ^�VAf�� YS�	��б�W2I8r�Tg���$\���r����h$�SZOx�'��sC�'ѯ�;<�rX��V�@J�]������5��q>&�|��*�
���T��"&|��2��k�_~i�k-t|Ղ��;�n>4y`��]T'��Ӏ^������Ќ��`=*��5K˅��
�W�^�jMSI�0x�������0�9�x>5
>[]K��9�3��Q�Ӂ��X8�f���i}�^m油!Kk���s)��E�(�������]��Q�Ԇ�yf���
#�����!�Ϩ�2��b�,��sp��z���x�;3�Q9�ΊOޤ:x��6�h��مpi��1�T��h�a.B��Z��ioVp��}f�d!a��s^~5q�!�c���+�26χw�a]s��`4�����7����J�"��h�y5�M��,&���Lx�Wť��n�<
��&�Z�;aXb%�E�6`���~d"�w�7BUS�����<K�
�gwj{IR9�:q����eUs�4]�А����bp_��\(}�@X�o�2=��^�m��!�E�j`uW+)�?�JX��#��}�e�	���Nl&Ca���@: x�jw�F�q�	�z��f�!�Nu�l��sJJ��w�l2�|�.M�*'����*�q�R����
�T�;z�~�K���MJ�?q<	ﺢ�0���z�|�y%u�b��w`�ݢ��aGkN$B8K륨T�n�UF��?>/xY� מּJ
��/Ȫ�(���Z��sd��9d�0
��G������JJj��O��Rft��ȥ��w?aY��0v��~Z)N�o��$��k%O�|�
��8�6M\�c��?#��1�������o%��EҜ_� 	����+_��"�;Q2GS/�
?Ij��-K���wjLP�6Xf��|t �]|&��J�}���߮�]O���%�F"��(�r�~��*����±.�q���ۻª��(�"�Xђ��+�'n�l	<����T����5v�q@�K�lg/��3��)+�6D<�},6�7Ux4i���TjQ�����c���4�qE��6,��m�b,��r3����Y�'v��	������V��46^�龇2��)�͓3�ya�ǀavs�m�a���F*�`Bf�6K�Д+C99�EP�,B�&�j�R�#K�x ��|FAHt;�q
1�]�>(��5EL6?���7�tQ�x �[������X_���S��	1���L�(*u�W�#�ߜۿ�}�� ���g�0�9��<f��jRj+��6"m�v�M��Ȍ�J�?jg~�vd�������Eq3/P�.�<1��1I������{2-r��n�l�R�� ٭�P�-�Y����3��79�5�}Vh��U�nk	��=�8�Jy���y�^6�v��/ļw����?��i�h!ւ��#�H���	�Z����-A�<�gQ�V�!�����}�%�8��<���ɔqy:dbg����B�n��+�ړ{4��<�j��z�Җ������(31Gh�����[�?�al1}��&���P5�$Ā.)����;HL�>�E{_�~�^j��}f��e(�� g�|�aՄ(���a�G����9�Ќ{�u�y�<
�s�5���Kʯ��l8��YW�m$
i�\�B���S�����0b+-nF�U��k� s�H��Ɏ󴴗,7��� ���n�\��x� G�����U-��)t��V�o��չT��O��2��mæ!�: 1pl؍�tZ���x���G���9�#-���ΐ>���o�y��{7��7X�OTF�AidFxJk{�t�?�0�S�a9�D�������(�
�*Y�'FK?�{�7�?��Qئ�%�xb�M�զkG�b����*5\�n�Q~{'l~��w�K7'�P�đdŅl@�՚<�wM85K7�8c�c+�"�A���L�G�|�I6g��.�,A�f9�Lߵ����A�w;aaB��8A���E�ɩ;,�=��/�E`���7p\1�0�fN�������~Y)��Q{�8�����9����r"%��Q�����/�X�w1K_#2��S�����E�*��.��0SC�՞�Z����8��'(9��n��[,��������0rb�.I+D�\��ɣ�k���K��mE�8�^8�_x���-���8,y��Q+JƜ�g�/�N���z�X��d���>��!��k @�,)�"�&�[�+��x��zsXG�9��f�t��cw1���x�T�VǏ��X%~��T��C(1�:���@d>܇%�!��M"�D�����*�p8���_jF�w�#�$��""1�>��-P�B�������W#;�VbB}f�L7v���@C
};6~U���t�Y�JT$ÿ��:	�}-_X��F�j�&��Z0}b���A����>d��[��������!2��a  l.	�:!�,�Jߛ�|@��c��)_�r�?��9׽'|��ɮ/�2�׵�#y��&���i�^�o[�]6V(t�	�qȑ����G���>;0犢��-a�W���9F��p�Ô�a�������J:P׋݃�o���sy���~@����'k�)\,�G���l��282��UB�η~ �I< �K���C# ��}�E���qSW���(��"+=E�MʺM|��u����4e�u����~U�Gڝm����NM����V�Cd��t��ׂN�rt�u���N����_�r2�����g���^H��B�2��� =P��6��e�S>!M�Y%*7U�M���*z�s��-J�	ڼw	5þΌGX_��P�1�K�5�WE�{t��9�7�� �:�5�����KM���/�c� �{\#z�^�-NJv)?���:z� ��)�.$&Gs*�{Ջ�$G��c���"Fnd�i�m����e<�(�?��Fٮ���T�8���f���5�MWG'�.Z��iȈ�V����{\�L��Pw����	+�����K��[p�.F��U$׾"^��"w�hL�,sg`jW����;���4���(H�E�3�,l%�,Feѱ��Ҵ�7?�:��xXk~s	V��u������9�4Z�Xӥk�B�,��0�eq7&��!�w.�q��?�1��b%��hЊP���/~.�A#}��Mc����}Wg���vO�r�y~5�m=� �ۉi���>9��	��"�a!j3�=n����3ӵ��A+?��tK�pӝ�/刯�?��y����U�%������EV#g����A�]�YU�N��.]� b�Qᾃڣ�3�4<�O*EźBk�'���H�T'L2]pPT{�=���?ԏ׈V8��)�9F���V��uE�q�:�%��o�P�_��x9��� &azX���YمC��2Š�Y��Db�4HȞ�&��m��w,t��a���ݏL�B%�*h�R�'>,]�|:&B(c�_�W��	kĆK�hV�6P��)�%�g!���6�����[q��)�O�o�/��zX�ki?���^NX/�'y�W�1���+5sѢ
?|�B�&��/�&<ȅS�!����0�U�O ��l��\D���K��O�m�Kl���ۊ"(1xA��t�k�|̓�W)o��6����y*�"�v�����RU�Du+�Kf`3�)�ȓx=hU�/�j1j��p����K^N8mg|:���*X)* 0V���^A�>�NN�M��0b^�l���Ɲ1��e�ء�[�s�D::�䙚0V�F4��q��&����^��lo�3B�ė��]��kR��|���,u��������?��~?YK�77������nQ��v>YZ�
B�d��|�s�=�x�C\���ik�Ŀj�Y��uQ���}%��*�G���b�N�]�a ��;�IIA��R����^�(v-��N��4lҗ`��$���6��P}�ԇK���K�ߟ��r�dZ�6Ե��6��J��A�x��mI�K�@1bw_E}�����jυ;��w�����H������3��1�Y����b�NxRH�sO�7��\�r�*��P�-��̄��ɚ����:�����`g��1����
s���_m؏�>Ǹ�"�߆:,�����߇��8[�dτ`A�h�qsGQ0E��7p�Lb��P�}p�P>�Iѥ�A;9!����C{g�v-�R���Q2J���������%�NZ��� lB���A����d�5k	}&���x�et-�vsQ�?G���;.10�$�T��녊W�,��Nۡ��5HMg�->���1-k� ��Y7��I���{}y�F�9��d�o슾�~`(�B˭?��H�>N���.I'��)�ڦ
g�V�#z��P�{ʟ�
�1�j1�A���W���Cb`��Q��[_��F���mZ���y��@\�:������?���ŕ���E,�e��X<1��0t��qz8�`<)X��2�����s!�&i����тz:����$���M&��~��.���?�Ӆ�;`Rgo��xO�Qyhܝ�6G�����w��Opܦ�ZRV�*�"MTu!zM�3�V������Q%�t4y��H��֛�x�D'��I��n�6WW9w���¥Gt-��@���J%b��;�C��nJ	��Z7S�j,i��@�f��6H�I�`��K�K�s��#-��ٖ�C��8��7b�K!bՃ1U_�s  ��=}6�YH���b�_�{GУ;���������jJJ4E����Y}
��|�;`<���b����d���biWD��	R����}���7��=�K��.��v����M�Yݫ3A=����"���˲�f���ޙ�/^�����Qdb�}�7_+�{tE݋&ޮ�)~\�6���O}�Ru'���8���>�%��d��{ uA��G��c˪����m=���������o}�J�H=��Xͯn���������'��ޠ���7W�*m�5׫�oyD��W<�T����"<C�S�}�ˍr�|�Z-?�o��=���\�	=���p���c����^,A�B����)KT��ƃ���Hr��t�0�m�h�k������B�`���|����}ڈ�~9�	�0�|�mC5���"jb�2V��s�dĞZ�@\9F�V�Y�vw���{6u��k���B�$�֧^(�%o�r�
��4��3��ʟTq,8�aqr�,�#U��~��*Z�;H]�� +����JO��U����N?/nƫ*k�\����ة�v�[���t�u��8sH��}޿�Er?l�6����!f>'�ybϸ�Zm4<���QV���J��9^�H~e��&��+#��|:���}Ͽt�V{),wG��t�_�b>>TL�7��qR�¦=��I
��(m��`�dС\���(�}����pT_�$�i8:�A��V�~�v+�|�R7��Pw],U��ژ�9����)6���cD�TY��D��_��3mMf�ܕ��x����gn��:`(�H"7�1s4٦;'�l~�� ����]��;	ykO�&��׃;��>'XV�{v6RQ���ʬhG��Oz�0���%�	��u�Dڏ�O�H�<�˶�Nʚ�C����X�_��*�(;�@zM��D̜���{ɂ��b;�	��蒹��%�:��v`R��Ƭ(�;�p���R��h���C�d�H�Z��2˭��� �˅y��^��6ojrs;�@��ͻ�JC*���Lr]�? _��ҩ��CAW��WY�+��M] ˡt��� /%ʋ10�(�`/�%�
�����ha�yV8f�,s7q9���]|F��qEs��ّ��Z�ޚ�&ƻqҗ��[��[U�W��!��IVd���:��S�u�)�T�x?�0+����o��	1�=÷�>)�[���Z�һF��t�
^�����J�6#)E�7*�Y�ӄXӺ\}�|�؆j���/�2����y���&�m�f��V�-�~��.R�G,��e���CS�pӯ�H�~����./~�z���$ҽv1���S���>���,�s�,��>?�����G�H�Y��y��(�Z�S��_&���d�����:���X�+_���ް.��	����fqh��&��j��� 9�A�Hq�Y���K-�a�5H����;뢇؃Fӝ���f�.Į3�2�v�3KS��d7��EA���lg)�}4�x���I�`����<6���j�ms90����"33��t��a����vۑ�	�W�z��<����Dr�j�\�qi��*��x%��i�o���CtΎn�e�sh�
�܌�Ȟ.l�BrP��&$�<�ЬBAa7n�\�vy w,{TC�Y*�Y�\����ME慚��R�Ac�k?�����7��ǹ��5�p,ee57����H��+��ٻ���hP��!g��c�m���|�]l/d����[@ࡶ��W��VC���i���@��-����Y�/
ۭ�g�d]Hϝ�l��	]E��2f�U>P�k�����'�pR�&g�EC�'�3��;�Az)�%rI}%�&]�8`�V��a�������~�T��/�ꍾ`:�rI��'�[������ ������'Q��3��*Q�7��
X	�: ��"�J��|���>�{K>�f�+|BlkO��Q���x TI�0H��,:�|6�n޷%V�e��h�$�e��ޒD^*KW�l�m9
h}ia�6��{�L��Sv=�Ǒ�S����I(i�@x@�w�^\��E�OT�g�]βb�&�ӈ�����)��v#�!�J�A)�|�����^����rl�Y!�]��U\@Ӽ9B�{������ ���47Baj��<�l58���A�4C�\�r1�Gڙ[��m�׸SnttZ�'U���h%�jh�ߛG���b4q���H�����9�力ع��ߝڨ"��,]�o�@K�������.�7�`��8�*�߿b�b�j�l���H��K���J��5�\�0Y��b��;C�����c�Ҧ\��P�<�cQ����g�k%~�~���ZQ$ڐ�ڞ`Ϛw=m�>U�� �B/��z�ar����X��4}�
�+�jhx��a��0�-��^�˴��9)H�]��(����5�q4a���1�1��}�oS����!�,�oל�D����K�0	�+��ü��1>�%u��`��`�΂�`�OL��/�.���G:�I�����p�Y�',L%Y0ޥR���v�Cvzb*�HǢ�+ X��t�®4x�,�.wu��z�.�����ڝ�D�5KXh"[�3fW����o�����A2�D����R�^����Jw�KD����7��-���ty��!U��.ٙot]BH$��Ǫ��U���p��h_0���|J��?p�M��E�̫fH	y�c���a݇���Y
��'�3�.����4��>G�7h*��
t1���ZL�X%�� �O9G����J��g-�T��n�A�}�itB�$�1�ɞ�]��D%�Z�nB$({�1,m�6z� 2��fE��щ���k��yw�Q�;M͉gؒ�px�/���v��7�o�P�0��y���v|�jsS<�$�;�j`&�u>5�B߂2��<�@W��&��/���e�$���i�e;�q�Hqj���%�#���I�&j:�Bà]��A�r��4��W˄4�)�,p!dsu�1Z��v�������x-M���#hv=d��H�&�վ]��@ơU�3��+�N� T[����n��{ q�x���{��Dfqz�ƣ-��R'> z�Bɫ�L��М�Ҷ:��Z��x����_Y�ќ�خk���E���|hB�@��^veOvx&$U�E���A� ��"4����-��|v [%s��k��g�+�3Q$�.�|�O��]ƪKb�]���:G��ƀf�@����O��_���LΧu8f/,���6��l�_
/`�K����sFk-��O'ȴXd�6��:qb����NGՁ��?���j�|S�����r�*`��|��\v�$L�h8�F�x�"g�`�ٗ����=e!�T4w��`���"���'�� ���|��GOQO[�	��a��/3N�*~�ƺ��a��Lԥ���8�8���|�zn�ޓ���,�����z�j�P�\��;��$����h�o�{j�o����yt=N	�Nh^wǄ��%?�8,�V N���_�����VT���a
s5������µ���X
��p��C���3�_ ����s�P�Z%���Բ/X���9f�c;1^�|O�g���}%gb�ߏ�/pW&8�ú��8<���X�4J��;�C{����~�n+�}�r���)�Bp�����I8��DA�b}��A&�Ӥ��c�ó�d��c�zV��[�|L�LR鵀p-R�4liZ�٩��ٰ�f)��z���u��2�_f�*�"����2[��y��f��_]�XpJ���\I�sd�QQ;>�@RB�����x.�\-��J��-�-7-��?��E��Q-VH�Rw>���O���[�t N#H46��o��?Ʈ�KJkrm���̇*�O�>g�	C��[�E���q���mR�L��q���*�F:��M0��njFw�!�d�K{l>��1�oD��p�Ow�j�z�4��pe�+QK(O��L�`�wYى/�A}7�5����3�h�Ђ��I��^� kH�ߟ����v��R$>�F����i�#;o߲Ne�6��)l�0�q�Vr+3�^��B��� �v��0�x`�{O$c��ׅ���P�+���Im���{{�O������x����h��'P|^oǯ�H���c
ng���wq�;띒�X�W���@���w�ᏨĠ:�0#��#����/|0���L�kKZbP��rZY('��-V:s|����t+�&�Vj� ��D�s�\��BH�l�c`;�G�6%r1Hw7�g*?po��S [.�1�P������}��w�jp��=|/bb-���Z+�>��!���8Z�&ͦiR4{��6 Dd�2�6O��"J����H�apr�!ϊ4i^3߽z��# U��(Q�ջLމMhΒ�?��j �[��}����D�
_}���ʦ��C�/�#���YyA�x�G��bw���a��vF�T,����E���W���o�]�1@�E(<�t�'�x��D:Y]n��l��{�U��3L����!�Y����ܙ��N�]�t�3(@m�������������DR�tP��[�ͅ�L���qD|��{�2}�п��pn�_�XbOy&�%J�񠭝�tȳ><�0�����������Mv�Q/�t[)z�)�o��ir���!��a�ئF�ȱT��M_��B�� ȉd��C+$>�	��~|k�Ų��w1��+��'�����0&?=&lD0�v2�$S�s!��7Ü,�N�y���� �iP�&���_��G�`<�6&���\X{�j�:��r��(� E��T"j�`k9l�Q�2+�
V������Vc#��E�E-��<`f�X<�RP�E_���j��$��I�"�r���	�l������
���7�a9�1�X�5J�q�J�xGOk���"���D�p�6�|�V�V7x:�-T�U�v��[n�}�Zs3��NE�J����
Kf��\���-�Ǩ0a[>�ᜭ H�*�"?�:�J,��Q��o���7+�Wp1/���Ek�ե�θJl0vX�:��&e�G��/C�d�����FD6vz��-B h|t����D�:�&4��d(���tcc��ܕcg4�Ѡx_;�^NØo�:]�K��y�XI�������A;D�8�N��]�w.�rv
6v~�Q}d�;O�#���>��s榌���NΚ\(��b���#���K'MVB�	Uǫ�M��oVz��iBk�4򳏳J���<�C��	깭#b)3>����P���>i\q��e~s���Ԙ�#�{������̀�쵤�AP���s�Jl^���c�̱�����B�����D��z��(Sē0f�O)���Ǉ�0�ˍ:a�w��?�C�/�u��F��\�bDZ}��o�=�L\c���G��$�1v8�7k	�ԋ�uo�;�̿���:��c��#�L+ `S0tQ��N�}� �������x�yd�@� �tK��%.o��Nڵ�'�X\a15��e�:D���F�d�[)zUd.�/��ޭ�~��ʷ?��tSۋzKQ ��uL�	k��@@�y+�hg�BhP̞Z:�DY�1��s���KE�p�	��ܭ�tC���(c�G�E��8f���tJy2��cT/����W����]����5���m�$�#�)!����zX�f�̂^6��4���n��\�^�/���e"ͩ��Y���%���O42��f����8�XΔA��/K�$�
�Ū+�3��u5��:��J�]�a����ӧK�d`�}���1�)D��9�|�^�Gp�d^�e����?f��u�?}M*��kV�i���:���Խ˯�� ��8���lH�>��8��С��@7`[(���A^��d�0�7�.'��<!�m��p�����&�C�+��ikh��0G�C0:;c�����t��5Dm��ښ�(f�ύc8��M��Y][�~h�[� ��R/f5�k\�)��/��v�}f"����&��g��ʓ����Khw[�3��l�Q��h-M��HC�dԩ�{4��&�B�ߒ$uƌ�@�H�v�ښ�2Rp�����"��2RG��:P4u�%���phU���>�������|\)���?m(�FD�g.D��D�x��w�։+E�\�����^�ݘ�u���#��"C�A���zR)�
�Z����e�O_E1�ݵ+�M��Kv��y���+3�>����p�Ѭ�.SU$�� ���	�h?
,]s �Xf"˥��#t�p�y����íI� ���u9I��4��uo�C�фՖTN���y����Bso�����sb'�?\f�<�%w�����h�Z^���V+i	p俅��� �8��#���:��ٺ�뎜���g�C]ܙ���6���P�����4������G�J��v�D��|+cu%99o�Q��p�؉��V D��d��<V��|�l� ƞ��]������-��SW�4]��:%(V_���y�
OsRn ���vb���h�p���i�㏷���C�
���;>��W~�7�:�O�f �h̞N҄�.�G�����uG�f��4��>��{�	|�D���TYw8`JB��}��SL��>�4�`I��@����QvFK��䟴C-��73G�|SДw+l�h�}��F��u}��+�:R
���r��<��:�uֆ�!3��?Uf2�@�H�¯��>���_vs�8+4$�T�D݂�=��WTLi��ʉ��7t�\�~�� O6���R�%-<�>�<��y-C�m�ϮoǤzď�������-q�`Y�錮���"�����E��s�x����g�,4o�$x�ۚ�dڦY�\A,��9���A��4��L�_Ϥ�g�)�X�YqQ(���i|9��z"W�~Y�DN��$��.���ث���TK���'*��$���֦::ǚ�qO�;���_>[����_'p��CvϲU� �pIj���62ׅh0��Jfy<B�p��쭸���}%���Б��I�\AV�����]�NY� <�s)rh�I杊T�}u��V��/�����(p4���=�|�J��]�"��*H�>39S2��q��q�Y.m;���l;��e�[=d����´H^�%�M�B�U��V`R ���ע���&��F��@ا�hZo?4v����I"'K�����8 �������M}�XeF����:±�ؚ!��4#�.�,�(^�������~l·�<�n.s>����|�cAt| �TN�3$$�{��qn�$��z��V2��Ctɵ)�N�"j��i��-v=	ͅ�6{4^�J��O�{G�k;����+H?�+Pjz�5ء�
�zGo�U����^PB���׀`����~?Ӛ�L�G��Ϥe��i���AWi�?^#�d�]I�Ty�f��?QY��{+k"��J%�T�Y�����$<��[�r7��gZ���g�G/��qnHoy�����N\^��3w��p�[^�%�,v!��0�3Tl`�2���e�+�&��0�l'p��
�y=�HJ��zu_
Ǵe�&� nzw�|�K��ˍŻj'.n]�/[,�m�X���ɂ�����?1�c��QSL��=F�L���:�˾�G˦��v�d5sÞ1��ֱ�����ʤ�]������u5��i.+���&�Xc�3��`�g^5�(V���+m���#^��� �K������:��QAܳl>U蚜�s��Ka�CLyV_̓Pҋ J���`�x�{9o��Z���*+���g�����"��`���KBy��ca�gS��̾���'�����\�t�v���eD�'o��5�� �������� ~&�1j���VHB���ˣ6�-��k�91���!p����t�[����4���$C*%!�7�>"�cΕ� �@e�E۝�'�RyC��35&P$��<�`G����}�Tg�D�nX�dq�M�p����`��C�I1��ԨD����3����a��-H@�52�;n�eT�[/��U��f�$� �$�lS��<U�o�&��a�*C��|�p�Ҕ�1���"�Ha��<?��4Rj�
�;�I��^��ݮ�ۥ{��}�\����5��7J����B��˦�9���J���)�ۍ�^��A���,p�d�����F�#�3��Q�=-*bx,O���d�*�4C�^a�	��J�b��J֭<JF�7���X#0��\�GSintu��ղ����6O������ݠ�Y�959���h/����ix)�MO�Og8���}�ʁ��� ��f2��f�^��>�'I����l���lȖ|��>P��m�oV���=��G�
;;���fPi���e�-l���	�.���J�r�r�zq��t� 3�U�ޣ��<M��.Dl��HH�[/g�K_�� s�0�XQ�@Z���^� [Ь�;��D�+�u�~|��U��Y��1@>��4 ��o�� �F��7�S�,;�;x^�`C�	;@]��[6Z�4�> 6�ڰ�\Hl���Z#��7�A�;�XC�H�A�x�`R뚐�� ������ZA��}�y������q��^�G�@��ʳa����}B3ܵ�\E��\�+"ֵ��"YA\:���9�G�`�����[�7�_�Ι�ﺗ��w��m��ڥ�o(��Z�{I|2�H��n|��l�9����� `��)��G�'��YX���ԧaO���z��b�L!QThQI#�NgC��ڜ<Ev;0Yϖ34��p��ey��V�J���𫚔�ӤR�)L�9>;�Au���Z�l �	hr�w�>��x��|U�с[g\VlnHV[r�TNK��:���)���	�B��d��>b^N���>��	��4�Է�s�\�ޤ���W6�o�s��_��9cx�m�pB���
@�C�2jLY֧8�����+�]���	M���W�Q��xAZ����.%_Ĺ��#�efC`"��~]e~����R���d²���Wp|fyE*U+'��l1[N���!��*�����h+P���,�4�m�!n��"K\z��K&��h��>���w��$Wp�@�Jc��Gc��!�ɼ�s��T�}�U,]ಸH����J�Qʛ�K+�W���/
�2�\�^�ŏ�㱮P�AX�v1\�;���z�<�b۰�j_��t��ղC�C )l�T p���g����0pΒ�~m~��'" �� �Q�K�=0\6�X�u%�4ZP+����]�*Ω���P�f\,�̬1�Y� ��YHؕ�M��*k뜾6��DO�=�k��ژ���_�nZ�zAQ;]2=87��-��pi�X>����V���u)�5Q�e ȆW�j�}&.c&����׭V>L0ZqC�Ț�p~^��.5�=�|��17e�XV���u���=5lGI��I?y�w�Knx�����B�qX9���`o�A�m.����� ��jZ3H ����r�-7��7��V��nޘY4����DcYΎ����<�=�����������4���>�Auδ�	�t�[Hݺ�	�L����r��������(��RE!
w ��{滏K�,�r���P���4��|8fu�T
\2y]�1: "D����O"���?��Yƿ�t۱>�M#��!k���yw ��G��  �<�i �EL�{��s�ߤ1Y3�.S7Rך�u%����g9w��Blvȏ3���]&��ǎ�C��V��c8�_a���b�75v!"��`��H�X�{��Z����br��&�=0z� �*���F����߭V�#��b����r��-a��*����4+���ōg��7�K�?��H�7T�7oԪ���^�)����:���f�$EgV@��`38LZ�֖0mSJ�9��%�kA�G����j�,��
��ٚ״�N�Ͽk��jJ�����}Vd���_CA�YpǶh^@�
�
o�i"Zʩ"?o�1��v�Z�h��#�vU��<��ۼ��o��ݾ⺠�pǗ��^�~>Պ�)��]-�E�4���}!5\`��#�1�g��j(&�}�Gk�[����ʬ�[Q�Çm�r�U{�� d�j4�����-#���
�z���;0=�)7x*0�6�X�Vvs�/eV(��w�̰���+����\���:�l��CðrWi��5���hϒ�U�&�zSԟ�k�ՍQZ�vF�ˍ��!�3Z�h�L�H����0�_�r"%nW�Ź�=��+��OX��
~��M���32p�i�|qP��v�R��EU.��U��S��Ԇ��hb-0��!����<�Y4��|O���u��e�46��|��ج�ƀ�U�.5�я��n��~�cX��A�����D��J�?���7����-6��R�+,�n�.>A��������5�R~0�ĕ�Ú/�b{=�/�0��7�I/McK�U�ExH�g�T��~X��������6'y�n�t�oPuM��j��;����e~*2�"#�vA[4�<O5A�`�����Ǣ��8a2Z}R��\6� �?�+���=�zW������4�_����7�TU�
QW�%�%���F�<5����àԔ�[��x��U�s�)�ց*S�S��p(q6 ���*��ck��OB���lH��1wukl��nX�?��R"ǃ I�3n��L�Uf��O��߉L�O#����39�ڪ�	%�
��f��F��e�|vЇ�?�R��q�/�Z������F~O���yY���6��C[��pq�$~H���!	��,
�B���9l�OV�F|�$طBqD��(Zj"�?�i>������ 7�f���z	�t���s���!o�h3ۈ�UZ�s�
�,�=�I�_�Y����o��F����ղ���ܷ2�3+��L�����v1�sX�8$C�*_ˍ�2���HYxYء�7��sqEӷru�-�T�qS�wo�3�K'�p�ÀbA�]$�P�]�:����4��1$xV�V��;��'�m(�-� �?�,�@ Xu�*l�{����5,)�E`��_
��O�ǫ�1�2`����ңE�)%��4F�驡^���ř����]y_:(#&��C*<���fO�<�����H�U/N{��2���T�4�'�H7)kW|�Ԇ��dm��8[��:��I��������_E>K��ƕ�12����u֦`�U3����Z���r��w�:/�m�+���uU������x�\��4S���m�I��[{���^�*�K����k3�����f-���Z �El�o��o��3�K���v ԘM�����S�`�j
��^��(��Y���:֬���+w�(T�<�V�1B}�Y~�p��3i.\/�Du��8�PҼ\!#kz��R$��k�Y�1ն���'�b-ICԎM�>�Q�A����={�I�˳H}��-'Xӹ*��X����Cc;q�����'�2�c<��S�_��y��T���K��kvQ�Q-*�A8���=��WO�H,�z������7ݻ�� ���p�MmO��������j|��*�H�d6}>R��<߻�����M��*�����?�\���Z�D���	�����]�j��?�Y��y�ÏyޱW���\NϦ�V&��Q����P��u�_1�.�@�F\�V���4b�5�V_��V�B� �80��Y�'�V�}J�L�-�[o�s83\�03���SU�&�r�Rg�bb0��.��[�H�O��gľ�,.��br6�;�D�N���t
^��F��9«5О��V���к+�KE�f���L�4U�J#�;�F�o��Sa��H�CĄ�n�k��׎EZ��,���`�!?���z
��{{����E���I��*����>�/dgDF��t]�USژ�������]tT��d�Sn�1D੡������a��L�8�\?V�������W�}J�Y�3g�O+c�¢���a.0HҶ���pY��͕?F�.wֿ�ک�<��z/ȴ&c�<�,"�U���u�N��o���S�Qqю�v Vd�c��*)*����ג��c\�Q��c��_�-Ю�z�<e?r(���!9X-˓<�1��,H�$mѪ�1m�,�B��6y�o��P��L�ӁɯܒT�4�<ҧ��]nT.��4t�"
��މ�su��xٓ�3�Ʌ�nc�H�_���rK�?�k�g��bv,o�F��h�AR\yڧ �r�綬�L|@r�� �ɦ��8��R��#�j�.�w7����jf��a��R'�#�K����ŏt�q�q��S*ea�k+�FS�ne��u��&6��
���F��L�wFx��܇�֩h���P�Y ؽ��>:�6��k��?�e������S<}�.�``}Zh��ZIN��'�q�߀U�93y�/R�K�a�.�Jm���٢�������śN����VO��� �����܍^�P����w������`�ZۜY�t>F��U���;���L�{,h��4��tv�������t�,�v�1�s*ׅ�@
C��>�� `�T�-� #��>{�Y����U��heN�����w||@,�����Y��$����<Tj�v����H�|K�mX#�;E,y\�eC=歘������HP0Q�q�-�u�<�녠J�T���WZb��?�`���g=
�W�'�uo����|Lo_õ]^ARBOg�������X&�ڃ�IJ#|����
vߗ�����Xd�]V��|�般�i�y)��b��s8�h@�ًn��?��i����'2va�;_5���,u4]���ض�V�/Qo�X�|BOiK���~��) ���
V.���=_��uܳ��q�ih��*#?�f�C>���x�ub�%�M�
��K������u�Y��U��v;
�^�4���F�\�P��������Έ��Bc�([i��L�܋c��a�-�$�Y��u&q�����c�o�b��o�Z`H�>�KW�CᒘS�-T�p�N�iZt͐��l�z�!��OtuH��R6-�U��� �]��$Y���g  v�����l^1��5��˲��Op3qw����f��:����9�[F21��<<y�_q��=v.��A��h(+��|C� )�|���=.�7�LE�%��?���>ߕ�L�|�V��F,�r�D?=�;o�(�q���dO�����w|�:���v��h:�7��˽�T�a�$�m�t���W�� �Ri�?���ׄ0��p���Yﾯց�x�����-lj�S��jf�jEoh��E���a�ʔ�0M�x����B�(�U���4f�V&�	K��_�sg·�u��#oC5S��
:��_���sG�t�t�K�rw#�������ig��dJSdή����P4Q���pV�X��~�K�՟<䵉k����l1���}l��hW�Đ���V:�m���*t�NOnWm�S�|�Q�.�z��8v�=\��:�4��PLԊ��
�0�yD�t�1�����ӣ���=6Ό�G@�qM��=_����8���H�v�Z�"{4�w� �)�����V"D��!�Ơ���ͽ�!����l^J��~-�C��UH�|c�[>�~t�<�4�s�W~EN�SK|�j��z�x�8��?J��<�ʩ26&��f����[ty���9�/�֨�N#J�~���~�J��ӣ�Z�=�#A�]���?Zr`�vIz%<@���?�Sdp%Ja�E� o ���U/�2��2o͜H��,H5���*�9��7�����C��h�JO�����d���/	��b���!�Q�a GJ�W�*��s�g�L����l�#Bc�K�
�����Vy���<�Zl���Nr<x��VgZFb���{h���W$���1F��\�3����1[lbGԂ<�<���"s�e6��&��A�F0��N�:^���d'��R�Jg� �E=�KySF��DԞ\��3	+6EmǬ��#�B�m�;���^F�v<�����g��<,�Wj���"��n�F�P� ������W��.�����T�*���!f����ȥ��w���ȇĥR�? b`X���V��ː�����xRc1�U:&�=d9��s���SZ&�u�B���a�����+�ZĤ�^�=��L�S��t��$��vW����j�~�clHDWL`ꮹ�`��������\�N�f�>"�86�Q���t@"���v%���eKa�9�����e� ���G�]m�i��0h�I���5�;�U��Gc�N	�n{�(wǫ�������gn���6P�[�YX-+"%����ˣc�1x@��SW�_:���hDt�ZV�CD��O0�c��O�8N�1�'�Uv�,$
���(�܍;�K�B/4"�k,_��h�֪+=�U]�k�7�,G(�Շ6�<�W� �%4ܤt�Y1<5�0]&���-���:!1�r#�F�;պ���"w����[�>%[�V�r��7�?��͗�^\�=�����/�@L��P��V@4�����$ؽ��@��0�������x����I�A��4�x�A4P�2"ʷe�_���"#5��Ew_��2�f�<(L�|ڋ�dF�mh�/ c��\ؾ8d�z|@xKSb�QG�v��9:��L�����}!�9��I7�����T&Z1���ǧ;-�|���]�T9��z#. �$p�\%�z9���Uù~��	`8s�.�/l��w��Uv,�=���J�M);�@��;sy�����t�y8��e����1/K?>.�u��Q���І��L�Jg0�߽X�s25s_˕�R�6S�/��>{u��Y���f�U�6v�$�ZG���'%�Y&�`�u-h)I�ed����޵2ױl	'('G�5�fn����X�ʟ�����o�;-��{�e�[��`q�~���ޑD�p&�lr�e�?���C���yy�|֏c���)��s�nM���6蹢V��v�@a�tČK-鳧"�{��k-ݣ���B�ڥ[��g�u��h�C���Qj��H.�ZUa�N _�gɏ���U�/��	X8{�Y=���~5׺��aT�s{9�!39c,�Q	ab�b��Te��i��
o[}����x=ڵ�q��Y=�%I��G(�{���q�(mx��
^��#!�[��!����J�GK�h�%��4l9����A6Mj�Z�t~�	(��[jR@��n8;�3���骜��+�o���L�%��kS��Mv�K�A)n�?��;��^7��`��G-4��:���bW�'/�}���ʫ����.Z����U;mR/�D�qÀ31�$-�oI�\쬽}��DJ4JӅ��P飋 �vm�P�B��u}6��ۋ�
�<��%��r�����3=Ѹ�eR��La��6/�O�3w�F��[�nj�X�	�8o����1� ��8���hꕜ�^�P�گ_ڻ�����)���X�f��ZtQM�L
��;��j."]�-�ۧN���P���i�n~O��`n<wEN�o��*ɛ�mR���;�e�&(���2.��E��j)`�g�=,j@�-��a��w(Vч�i(S{�<�"ue"ΎD|�����o�	���ޏޗ�tKz��^���ѻ��M��q��1%���FDmм1��g��o�9�a�	��q9�x����g8��L�csnKt��*≇�a��U��]m�݆�As~뜰�fS��=�����/�^�Ф�Hl�lj}�>��{�+��	#C
fzPU��C�ǖ�h����W������E���g<��U��'���Kn����;��Ђ��bQ�<�'��=�����|��o��3$��[����vœ�f5Ec�I��-O���L��Tp'�*��\F2�Mx���ǻ�"�,�0ŀf�+����)l{ڔ�H��*��s��ێg�UQE��Ys~ƚ#�-�n���[�ka���h�������9<�����!^i��g[im���Sw�j4ɸ|Hؔ�O������/�3��ǿ��v�{q"[a�R���M���\��,`B�❲$��=�7��k5cX��2v�xYb�9�2uׂCm����f��!�2��+:{���އq�z��^����c�� ���Ч�.�<X|��O��$�ƈ��a��]EUVњ�n��2�^��>l#I���^��|zN�5y��E�!��Ic�8�r��/�V_1�H5�:�S'�g�苯D b� �c����JM*}k��S?c�j����v��dp4MT8��U�e���) ol+*b�4�Ⱦ�T~s><$\�e�������rc ��#?z��e;���π�#�[��_��t����5�`9�*���8N�7K��64Za�j��.S~��
�W�|�@�|z�a�Aa�'�R%߱�\b����_fg��R�6E�e\li����J8ȶHU;P�̏*26(,J��u�_���Δ����l�@�� �Q7N?`�`y3�)q���r#��03�E����}`�\'�
���Z#�A��9�����#.ǑrХw�����C~ȣ^�<���~�{��RU'�C��2h�����|�#�U&@F2�ޝz�y�킔/QPm��ؙt����ZotG$G)��x��`��=dT��&�bO��@e��z�_��3:C<�́��N�~�.��W��1�wĪ�/[i������X&,����\5�t�&��ޭ�r/l��l8[g���D�!���rMO�ۈ����I�Ż�n�?5�EV C�T�o�.�w�H���,���#�E� �C�q3z��ᶙ�z�<f��K;�o4�'77u�m�^'�]�b���nZ�e�	+��j[N<\9ѫ�!G�
pF�5�q�p�@ʥu���1��{���ѠI�v�x)1�i��A	�&��I,�gA�
҈~3 ��-a8�;��߻=�ubGo��-$�^�F(U##d�w��;�;�KX���Dx�y�MkVB��P�6�S�8"&s>�'F�7��"�����i��O�Pj<�k������S��l� �Q1Cnn�r�P��G�t0����<1Z;B�S�m3�Y�o���^��+�c�s)m	��k���-��'s%��e��R��%�Mc�]��G����d��@ߋhO��܄$�;y7h��t�����'�B�V �]����'���//u��.�����a"�G�� ՝��XX�:��4*�W�ifz-�+�� �/E}�u۴�iu[�v��Oh�R��=Q4��y�����0ߐqs3C���XW}s�Rr�u�f?&K������~���(��T��n�=��r�ne�B$�����]w��\��0�S�l�Y����0w�b���fx��v����6���ۑA��$X6>��^�� ���{�L�8�UO���?Ӳ@�v�$���T��"ᦦ�UO��E:��~+�R�]t~���1xA���+��N��fʢ]�*)Z��06nZ�!h�G�irH}|���-���B|HjS�T�[�i��K��Z��V�]f�s,-(-�_���2�M��` ;ۂ��h��S��5Z3�:.{[�y�����A�E���g�j�;����Z��v߃<��@�t%i�rJ�������P���t�3�Jx�H*�����VF�Uǫ���<�k�z�F�ב�9�HX�z���0U�|��?h���%�]ڱN%Hv̕�;�������?�� ���b!�.�� Q(�Rۡ����~�U������c��:BV��s��'��"��>zb�Ft�!N�������5��<��Y�b4�]*U*4��`޼�57��yd�εVI��[�MM��M�1zյj�����m?�<Wlx�R��RE�����w�"�<tGc.��������u*ބ�ǯ��9�?n���9}��M5�MKW�4��6Y����M�G��$V��ߧ��mg>�1���I-�?Q�����須��]��g)x�=�[i�~N5wT���k+*�q6rHاA y� mY��%���ޛǝT�{��>��~{)�s�ߞ�5��wz���K��) tp������JL��Y�= ��� �4��!�Wa�1:����8����jBE-Ц=�!�V��㐀�[��#�g�O��U�g��:)��pJ!��:�bV
Nf��Mq�@��|"=��a�54({e�~�#ooi�⌳b�:eg+�~p�P�_��(j�X�q�|e:Q�o�õ����yEy��>�B��`\�C�PTz�ZMlr%w.S�6�Lp�K������ӣ����2��W�6n�KC������ij�5��'�6� `k��<��Ts,��|5V� "����_��2�u��c(2آ�����za3��g�m����d��	WM� ��C�)�:?��7�gd��!_[��!!��dٔ�w�Xճ϶��0 nR�	,c��N̡q�Ǭ���tۢ�^��s���~N8`�jJ�pT�e�����//\�X3���=��<^M��r�����~UL3q�����疃�J@_����\�7v���p�\V2��h�q9\X�s�#�'Y��'�Bt�%k۬�Z�L���u�^n��2�+ j�f�x�Y�ṑq|kN'����ф���A\��U�3&��XkJx� :p�"U�&Wt1�P�?ڧ�|L��0���{pI�@��^�$8W�j�I�8@v-���w�u�ێ�'�Z��_0W�eW:u��]pl^4�/��4w�\��[����1U\g����h��k]�qvݣ�	���A��&�`؉��m9�}TJzl9�5��&�����HƠ,޼iv��f��p/p�Y;&j��
N^�u2�L����֖Y�IN�H#�YW���XJ32T��ے_�&WJO�o���H��O~�-���?f<�%����G0"�Zŵ���s��S���B&�Sg�Dzc�RA֕Y�k�I�^�#�bv8�,w��1����ݚ^�Z�y�Vs�?4)c��JGM8�d�ъ��-��-��]� �����{\9hS�sT^./	@5CxȀ�.[�G�Bs�QvGzds�s�w[�6"��W<���@��N�t��G�v9�Z�d����[���䨽ذ� ��(W%�o��_Ѭ}߈l�kD�q��ǶNn��$~���2���1`?�ݦ(/Ի�%���A��hﯫ7Q�>u�BN���R`��=�]��m>X:�4�(�=A�4ԛ��2��9�(�SC*�fSX��G�7�0�jHK�tt����Ð�� O�x ̓�ܝ.ߚ��N
Wl�W��J��t��1u+Q��r�^�7S��V�/�Ǎ�jH�nQe���+��}��8�}��Y��$b�FU-�0�I�/��r�C�\���m9Ԍ����r3��&�)��m�-cܤ�V؎�U҈I%옍���y�S�_�U� ��wU~{=1�}-�����G0<:�k�m�0� ��)ڜ��5�*d��z�oBEk�o�-�p��DG4��R�,�A������|�f�N#�*_M�rr�(k���|h��7:c���Su�t7������Q3�u11���EK�6s,����&����i�`����k	�Tlw>���C`�u�EJ���R�lY�yZl�t���U�hM iKb���D�p���:��Rd�Of1���;\�'��10t�h�B��PٛxG����~����c{���.#�d%���q)��zH�y+��<NQ���^i�÷B��AP�Է�eq%��mY$�ҩ����*!�Y���4�����q�3=��`�(o@�=Pv;�����g�p�K�4Hf~�j�� �#-X�􉀛�9��(Zq����U���T�j�u�*�IQ���@_��	Nδj��(��u�0 [$"�k +yx��RÿoK�¿n?iyz�2���|b܅V�� 8N[����U�Zõ�`�oʹ`��Kz�2"����=������ޟ����_A\�5ȉ��E=ZOɞ8�b�q��ȧ��������..O�����5���i8��KGn4�t�o�ε���,)J�h4�g��Hӛ�%�����!�)�̞u�O�.�ԓ$o��\q�2���~�QEr�@��m�=w]>�g|�1n�w3�8WP��8�?8�a8��3�J�Ѓ��N1��F�5ذN��*��!���G_[0�܄k];rF���O�~P=�9�N	�P^�yvK[�[D�J�h��d�F��(H�@�%ɘFk�ۚ����!���i)fc��Hoܐ��~�`�R�x�Jf������m��d龆��G͵�xe�pӏ]� ���b�Z �
����d���12�,u�C���"�����
�b���,B�К_?֥��ug��M�"������<�m+��rK�lk�K���tW<_٬X���֯��~��V�`�H�i�d�5��]1!P"7���X�tV~�qln�k�O�9����:H�Җ�f~Am�QG]��xq�UĈ̀_=[�����`_Hz�!��'3�����z� �H�c\Xcp'l&)gl����$�MP�d���~o ��JTVd{	�Y814P����4!B���������$Hz��C}x���}ĀP��T�*��r9�Dws��h7�*}w�:�v���8��ď�e|�!�].aE	c�mv���J\�aXߜ/�П3Vl�u�W��q�9<�j	��^W;�_���U�ȅ�{YG�%X1�� [�tE�b{3���5��A��H��a�RQV�hp3ÞPܬ|�:l/��)ܤ���R�&
�b���o����=ǵ
w��jz�%|A�]Щ
�Mj�{�Dy�U��z�2@�E�x�}Pk~V�h����~B�U㩾�?�v��~ZUv���O�{��0���Hw�T���F^��6j竌�A�s�U�G`Keei�lt��r ��cp�7�sI��O"�q:&���T��]v/��g6�Н/�� -��<&oʧ���c�g�կc����E��܌�;q�'�(�L�x#l�����6�q+P�^J��;�[Lx6��"��,o��WBۣ���0�f�L�P�5 ��rh�����IؚB��E��ݾ�x2�>��GS�|�`����i�2x(�qez�	�0;R��`rM�3 ���!����r��j��(��*�&k�J�m��e�za���������Ȇ ���Z.���T�[<��ٴ�r1�k��2!���t��59���$��!Bv 	��{����h�0�>c�
�M��"ެm�OD=az�#����p%Z��o�&�p��W����*гuz% ~!eF+E�|�x���4	�O��>CXU�Ґ�[�aǟ�s ��$K���*C��4���'�TtS�+��o�7���HD�O|ٯ�1��D�cK;vSM�q#�2$��t���p~}m�)�Q�爐\#?���j�v�����8�Z�=}F��n���p,��z����F��Y�vU�P��x]�F����7�=I�5��n�Ӧ����?烊aIxw ��Y
�9�^�K.�h�����i�OQ$/T�]���L5[�.��+���[����PL�C����s):{�w�pZ��˵�Z���I���~EiS9n�޴BMr�{K
��xxu���,6=�TGE=5��1W�S������h�O4'���D*����Q�Wb���~.��8��SDjc�*�Q�h��VV� ˆ���[��F٤%i�o�8�«s(��
�G���Y1�cs%\q^o�2��wm���?��a���N����g�G���Ę�5��lci�>�W�1$�s���� 2Jv�K�G,
O�ԋ$�$�ir?��hy޺��[�mz�ԶB���L�t���{�G�T�����@7{��@���hۯ�����A�W�H���exء�-�1pL@��;i�#C�8?��'�e{|�֍�f�Il|~����d_Ȋ�%�_��s��6���Ŝ��y���H��38!�]����,��70�^������>�K�ؚT���k�4�̭"r|�ߧ�h�a���+4���nٕ�BH�?>���	��)�)w���ȷz��x�OIؠػQ׋/�1�	��&6☧!���[J���Ք9k��RiFb9��
��82BPgְ/��n�ZP��T��S�ɒ6 �6.>R�1G���?�8��I�j��\w��'���{�~)�Ԧķp�ә�O=b��zeϠf{�r�d�h�pdzF.$�W��gOk?*��Ȼ��K�C�V)�z�U����ɕ�	7�J���B��=�~bђ+]+�Z鱉'�8�� ��K�=p~�r�����ګv;�(E�hC6�)�ʅq�g~��7�&"�i֠�k~m�e{oc��^uݘC�D�~���-��@ؠ�Q��Y*V��M,�ͿXes�!k�9C�Щ��{�[�I?X徠����1���IYA�nmLt-�$��8l��*�j�ݙW��o=��3��E���\*�O�3�]ɚP,lH�&������q]�Цi �M�g/f}w�-���Y�t\\�-QCg���Zz���d���g(����fRD/�O	���N�4@�m��jg)z���Aߋ4����3>����p��k�.��f�a4�őSg6p���a7�������
p���f����?�n���C�(��V$�k�g�����wD�}!똮٘����s��+���y�E6�u�i�_�AZ��6������k���$���S��#+�jJy��]1[����x�C���@�/�l�,]W)��XN]��t7no2h ӔK�~k���=�7/�� wg �#~�U�o{f.�!ezĵn���'�%�1xS�r�-��隲����h��O*Z��N��+�@��Vo#��F|�B|��j��幇���w�RE.1_�G�����0'^���?Ώekyz���d5����l���s��@�O�!�w p_�&O���:�u�D��<�%���=r�u]mw���=�ʞԂ)��ͳ��4�l�_D��4����hH�-c���/�k6����L)֥#[�:�e�~c\��>9�1o�?3���h�#V��ȃ:��/}�����v����;������L�Ӽ}=%��9�01Zi�p\`,�+���8�"ͯ��d�@�B����|t��=՜s�YK�M�&�Y�?�x�%)pTb���b1�@͗�EvF#������C��*?�ţ����{�N�+��fB ��.>a�:��u̍����5˄y�����Z�6s��x�����N]����������#\�M�#���Z�d�Y��o��j���:�Y�~�7��F��:�-@���<���T�=��O�4ģ�R�]���A8�r��G�w�+���ټ�H<K�م���ZIFf��q�q��q���V�������,�;��WP���b�M�	ּ!�����Ҷ�U��/Whݡf�9u�̟��)Z���������_�����So{�����N�r@������#mK�
0#��:v��D�1r�f�/m����T��?����C�bs��[xC)���U�\x�}�/k���� ,�Bcf���)�eŢ
l,����o�e��vm]ől�ȮC<�ߤ�"�.Nb����G>�i��>nڵ�P�	j�����r����2�	���nr�&0$CO@�� ��тKb�y3(l����a!�ԓk�k�n1����!Ի�����}+#�9?�Q���T)��� �n�!�ǵk\gJ��*W�"��s\Λ����(�c��L(�K�����!T�QH����Ѽ�q��R�DP_������1��7/��$��wl����Y������R+��e�Q����/p�h���T�Q��`�Bqp�y�V%�5�P;�b\i��.���H�`7du�>�W�S��yy�:�Y�bWG����X�f'��4�=S5�?�,:v���)l�ꥋ:�"��q��"4�)o�ϵ;i��yQj��<�I���"��Z��(bZ�������_�O�W����}�0_��o;$�{�B����?��_XT�U�?+y�B�{�ޙ|���E�
�i\@�؂H���8�^K�AU]�_pz��?���f�5vcd����^|[��n(���[s9�MjOu���W��Fh0��
���!���5c�Ӈ����Mf�J����S�.���ZK�:?%,u��E �Ss\�j��OȤS,��*�вy��l�S���z������Y�U���~DT�����Y��!"u#OZ1�҅^�2����yU�1w�li��SnGsg��y��o�X��R:���Cx��g����Qm�{^��/t�̥w@$��3�/�D��6i�ȡLw.��N&�<s�]��2�u�V�ѵg�+�k�\��8��'�VcOR��ͽ/A�i �g����A��bY���S�I�Pu3GD9�9�,��6%�8�\�!�'ߜ�^���D�G�4���2�h��a�2-߬��/�ق���[��v���1C�o�=���u��?��$O��z�)��� �gU1x� �3,f�%�v��f��XA�<E�=]���a���D�� 1�)AU�SA^���:�]�wo�_Wts�a%�x�>�;VO9,u�:`�V�8��մ��W!M��|�9d���TjE��[�y��RE}��_<%��P�ށ���8߿��B��r"� �h�����ed����ap��=!?|I�~K��r�21v�t�T�tˉ-��7�]7�{�Ħ��[���*�С�H$�����~@�N�#az`I�~��U�Ԟ�j����/�<��ˇ��h?�"������lX��E��ri�Gt�N�S��b��^\�1��2�r7�Ă;!d=}'ȥ)>!C1�[»_9��v���1wC��l��^vI�( �n[ӳ��X�ߕ��1�k�Y�z�9tmf���i��Z��Ň��e�(�M�]R}�GV�I&<ؘ"��}U�V���B�:��OeĊ�qQ'S��	s��-l	��ee�W�*��F��-λ���a`�w(��=���0�g�N�ȭ�6flS���o"�c�r������ a�m�n5 R���Mi֏"&���Q�s���	�(F�"���w��)q��ihf�0�!�q�ЗF���H��|�$���P¹BE>JcCb"��F�� T͏j[�|98K���������i�I���u"-��įӋ����8�?u��W�J{<�ۃ?GB�0GJ���?�Vr���D�>�����X<�$��F�[w���m$�R��1�kL��s9�;i��T�E��i�x�X�k�=w������Ax#�nf���'QT�l?U'��&��8��	��xP�^�q������ZD�G\�>q3&�廴�K��%3�+�����B�ܔ�?�����C���zd��� �S��wj-h��E�g�SC�|�]xfm��eŇYo���w\������7_6�}>��-^n��*����,5��ͽޅ�;���-UH�M�.2�S�Hu�-��Hj�U�H{�c�N�X�.|�cG���C���]Ko�j�*����BW���i�nR�8Z]��D/���" ,Ϙs�����
	�U|��x��PX���� ��1(Z�b4�ܦ��A�z~��tJH���{[/
�H�F�ps���"ʗR���A��{�!N��yC(�e��@���:`�5
���Ψ�������Be2���`-����ƞ���C}�S��Њ{�bv��z����7�ǞQ,� -�����B�5k�&w���-�^/���=n\���V����^~ﳨ(�%��6�I�#���XƠ�������AJa�3D�5��2>���!����L+�4���@*����c��b;��uĸ�T��c��H��3\��d�C�||���rMF�({�\mi,��7�|��@s��W�[$�	]zV��^�?��`ƾ���3#sLw��/%��%&L��R���h��N��;���BO�E1cS�M|Y06}����v!hg���*��{�OA��
b׵�逸s��C����g�]X�.��$���1���D�S��U�[�\�V�A���FQo�����ـ���W�>��3|+K�����V��*�9D�
���Տ�4T���K�}����pff86�f�b}�$O��y���K'qRR2�rR�.~ZE�RMi%�v��q��(Aڵ^A��a�뀳GY�5d���Y�V���JT��uL4��z@'�⚇��^���t�sׇӭ�~��rrʀ�1.��iۄ���O�E�Yx�?����_�.J_P����\������ݕy�Q��>�ÌR�՞�����K�bq�,�q��lAU�MO�OjZ{}��s�����̢hЅ��u%�u�pĒ�A��ME�T�%�$�A�6�o�$�ȨF��W� �I�s�@�͹bV�"P�T##��y�G؈���X����Ւ�ɠ���r�),�=a3kT�"C�2�?y��i[Ӽ�xgy~�yKf�S�������Pw��2%��)���;���J]����M+`
���f�/����ڗ.�<T��0U+0#-�U*��sc��|g�8��^�.J�wČQ����}K�f��2��e&���Zt�Y"@	eB��\��y�Y�!u�l�?�u��+�o��0�[�f�)K��O�ܟ&��_s,�T���.q	 �{�Bf������Ϋr��>M�ێ�xy�GۢB&��E�Eǫ=���ҼQz< 5��u�����z(oހ�E@�A��_k4�Z$ÛpEv�B���g��F{z�t��sj��LS�!�U�8.�������s�x������;{>�I�AOΐ@R�g��ˀ��ͬk�3����8v�G���k�M���&���`3H���r�!7�S��ƹt��)��;mV�o�0�W+�����8���Sj�H�:��䐓M��Ñ�l�.ƀ�(iHŨ<�,ɩL���,$�<���ߙ�(���(j&�s��*VD��)̔��|��%}}C�U��BtQD7	�]C�h��aX����-AhQ��� �f������\k7�c�I�$�: �x$9���5S_��� �y�p6*ĺh����e\��=F�L�pvLC�j��ޏ�����QB�+x!�  J�?G��ŧ��3�������}����w�V�j0�8Ю�*�	�>v�d�E�с�ҥg!����o@Ǐ���{�!��.�a#6�����Ѱ��̷ҷ�_��5�L`.O�u��ls�	7�q�Ea`7?=6N����O�z���h\x�\�(�Q��Z.�yi h�rY��ty�͢,L��W�]XM�w=Lj5�L:�~�$����Xڕ�u���\7��V�_l��"�9�{��4в���7!�@�/����s-L��H�����h׃���&�O����������f(���$�|� ��\��)�	��I���W��RA��bg�/�����m�DkJlv�OK�_ƻ�������g)��}^w·�ϴ"\��JL�D�eȓ�k@�	������I3��Wc��!����8|�i&r��|����߿Cџc�
H�;���Q�MH�㈔}$3Yj���\�F	�TBs�Huϻ���H���{��47�{%��Hl-~����Ph2�-J�fI�Sk,�+��m�@�М�(�e�k�������Kx��=�b}j�3t������7��	���z��=��gk܆�׼������+�$���s˻2MC��#����%���Y�M��}D��*�����Bخ�(h?���Q" ���s:���~�cg�=d 8�#����x�hfoa�	HG�1��R���=���@�R�~^�6X@��{X�>��4❙��e��]�ī-X�@��qc޹��aU��Wug�̳u�x���v1d���ϩ%���g46�������Ή�`����+׾�:;���]�#2S;�sF��m��ߊO����P��I#癰�DYU��ݿl�&:(��A��(�G�(��}5�qg	Ѽ�+�^l�t�R)�h����O����X���2�)h%�G���/���pn���ռ���ׅL��JC�L*��� �U��f�7!U�I����uM\%�5�o�>[g���)��NX���\�Ʀ����=��!#uf����D�w���o��4��W��Lu���(�^�C�Jp��q�k<�����ΐ�O�F��
�\#B�9=����D��$�������X""�h�R�d�W�K!$r}h�Z�b .�?�>.C�PBq�K&����)�Y��7�8�y»͙��a0�2���3(��j�±4�Lʰ,Hh�$��aPR�
Lm��G�:Xw{�������4Z�1	+�~�MwSd�;�����9��/S�M��u��ysLQ��uI5�E� ֏R�M�B<�w[�"�k��E$���~�%F�g�f?��(�� ���g-t�yK��]�/a��3�奍��fE�d��R�(Ntx%,�M�S����P�P��h�dF'0��N��Im"��g����[�6d�Ӽ5ꢆ��Ko��ۺ %˙C���24@�y�c{����Ţ~GKy x0'� s�i��IW�5�|7��X�so�C�r9����;����M�*'e�H�ݕɘUp���u��� a���gym%��JJ��������_���T��U�6	�0���և�\���J-Ј������"��=�sTgZ��&"�{��ڷ[S���)pf�$� ���HY[�K�@��b#�~x u|A@�J�pN�.�:��gz'^Ν��o�;1���%n*�"�'�D��L��I���	�(�:+��^�;#��M�d�kw;�+]B�r�+0uY�R��ƃ[�u0�6��onX�9�<5��UǻQ���v�#��@���ň�Uᷨ}���ב� U mȕS3(�k�ճ�
���T]��D�n{�:�9ȇmV7{|�լ=��K���-_tA�|!�k��юe��K��D�H��>�zg�J樭)6#�_��4	/�@�i\����J�آ,Vw�?W$?˙<�@��&7�,��2�|�K��%�bj�������VU(ᗥ�g�1����g���H�$F?�	����O{t|�M�� U.F�m���׷�J���@z�s��|�'�|�����{NL/��Є��n�:�!K��;�ڪ��t�?d~�̔ol^'N�;Y'�f]s�UPIa�����V�����5�_��2oC�5�#����H�y��lOE���%Xs�Kyf�n8�i�ܝfQ�C�����:��
�g8P@��c����DRo�sY�s7K%�u���� u�mu���T�=�E2�w��r��x�U�˲�`֢ڮ���|G�~J�����Xu��=�=�ǋ�]J������> ��&��	�y�>�)�	�]��1�IE�]��t����0o�$�S���j%7���V8݋�ƥ�l������!PV��r�>��e�ȈX&tv� S�t{ڧ�8���O����r���-��E��#�f����3�9��:4�F=IE+�BS�P�Jl�d��\@�bx�z͋cI��z���6&)����»���q_�$��x�f�СM�j.�	��9�%JÀ'b�$��?xϨ��8�K۶��A�Ez7O�)d�W���~�ϕs��!�1���˫��+�/'!���e���M�4C��5h�����"�;E�#	Ȭa@jU�ŋ���A��i�s�J��rT2��5���>P}�11�,�s��`�=�#���y���f��s�1�E��!#��_��ck��zd�U�/Ad��7fz�@L�!���:p��Y��'b�������%,�o����"��ҋ1�Z���d������L��z��$6�8���	j<'�@O�
��Xz���L��?
1��zɰn��3r]|I�א\��~�B�p6����t$��fkB-��H6C <�1}�|b�wj҆mt�� �B�^�W�ZQ�3��&jk��z��=�&Z�sw�;���6�<�)�S�1����֍�,ļ]���f��*�*س����g섓R,`��n]�ք4���-q��t�tx
�7����NA /��-�&�P7��Ek�b{E����/��d�Qq&1��<x��.��Y�bn�8�C��&�"0P���`o=��3Gg�=��ՌI;�pH>_�9M�qq�5�(��N��&u�k��v�~U����}�2c����dim_JPr��{8dAt���DZ�<׫��LtAÞ|�2ǒ���5�K��K�o!�e�Q܈�;y=��J���!+ꡫ�Uz!y�㾛�2g���_4� �Ё��2_��tx���P�G�H�����X�Ez��U }֕����z�PA�=���YU�&�
�>�`�QlIF�����P�o8s�vy�?�]���JC%z;eO��\��]e�&�
������P?���T^�y�J��Z_8�~�ݝ_�i��������A^1�i�D�{�|���}��ȓ��o�J��𺡂�S�{{�C�A�],(4�����!�2�
k�xC%����%����0W(Wtx,�1j%F��3����������7e���M��f�R�����R� �}�?�D�;a�ʿ�5���{���������'�^�Z�5���xx:_�	���j��pB�!g�*:����{XR�kQOC@����*;� ���>�����໚dǽ��^T�� �[���Y��X/�E�V��1�1`;�ؠ�kɝ����B�tޔ��9?�J�!P�4���Ұ�~V��2�D'�ZT�����6�!\���2��Ic�@��0��3f���0:.ON�(�s�ps��*׾9�<�^a�~�|9V�~���~��6��Q)����bgm��+�1����`��F�py��$���Z��C�����`N��rɵb�߽Zm�ɻ��� �݈������<�V����렻:��Hl��K��c����������mǷi�	j�z	_'�� !/V�ff��#�s��eQ�'���l�F~�,[M�1������1�(�(�G�f~)Ga��Z�XP]���l/���4 �ȃrTUI��������!g�&��]rs�X�ҌlrA�Μ�L�h�n�U�o���i�"~���Muw��5a�&��QN�h�^����1R�V#�����/���������������˦�N�:P�w7��<�B��+�M��c$�+���M��������Y�­���#ަ�)J���4�H� �d�O�P�V:*3����� �$V���}Ē7S� (��#Y��W�ɽzS�*�s�������`%���k�Tj�!�5��Z*X:0����o+�s�����^��Vh�3�l�&�Ƚ�R^G���=���V�-#޲��~nf�ç�n��<��z�j�L�p)�}�0M�"�$���󆒲�RU�r���r�#`�C��9�{���h;k'���y��.�t�+MS u� ׭e� _0�&��:�$�ߦ���zF�
��uT�XCࡷ�NP.DO�3g�לR�A%�Q��e���K"�RҐ�~ɞ�3�~������i�n5|^��	�3�xI�|��>�&�1��5V���5����YBf��y�>m���c��d����:^�)λ����`�3����8�+}M5�������+b����}N|s�(/�T�w�s���Ȕ��Q3(���:�F�����2���hh���|��&����3����bH�PbWU�D2ヤ�a%�
��6%�;�Ec�^�k��ǡ���G����W�����a���G�t��n�i��73�����v=Kf��'����5 �ti�i3\E�i�Z5���	F��tF�P�a�zI�oS׊�"�$��G�u%P��]�v���>���ӻ
\�����2�R�SB�����o�a��1k�nᑚNs�%{Ct�?��ǌHj��S��I�y�[�Dx(�P|Gc��I (������'6:�v���VG첀��� 7�0I�_��r��~�����l���E�'���� ��˲ܧ����a]�,['ſ~nh�?r�!���_�=[)0({��APZ	�&�����&��in�Yn��$�6�	�`r#���e.����>�)�Z���Kp�[�;D��@9�c.�ZxG���+�uE� �Ib�6'��h�|Q���z_���xQp����#��`�n���_\�@,fu�/j��IE��Ո��Mm�
Sgek��wd+_�X�� ������Y1Tz�Qc�A~R-`�1U'��
��Cy�D��QW��ǟJدhd�3rF-qS~�����6p)���xy�˿��O0I3�� ��)�\
R|e/�ѡ���b� \��������ľM�z��&o)�{WE@� &����P��'n� �-xE�jrNP�(E��t���}j�엧đi��@��?����ǣloz6��1#�ٻ?N#��`w[����"��K�_�we�E��v0西^
����в p�gs��.��@G[uIw�B�AwI�mԞ�5:J>z�;��PK:u���X'��jiR�Iq������I)��f��Q��;��Tמ��i4�mΤ�sEPs��l'B��\ڧ(�ZBKҍ���~�~��cLD��?A���u�yp�[6��Ü���Ԍ�1�{�sV�	�҈?��g��R��[�Τ��Su��.^�j�P��o����_Ҟ�I��'�R��h"�:Fz��j/ϳ�b���zߠ��X�$]�>�ˆ��~�u���y��OM���/_2) iUA����b� v�K��V�>8t.�;�e�XrZ�� ;j���f�U|���t��(�#5bJY�f��������s[��4�`ˮ�^�v�f{���%�G�X!M�� ���΁rG��S��7ᓺ��D?�G���Z�q�*R��#y�Nq�H�.	�oe�si}�A<��g}�(��<� ���X {uUY�s΄���&Sɦ.�����d`b�sW~c�$D�G�R����nN�n[2�	"g=U3�N�$�5*����f��l��D4o� ���(9��I�ɤ�kͨ�|ה���M���Գ��Ԝh�Ȟi�<O�If���mzv�jE�2YbT�+Uu���wC�*��6���9k�`�/���=kS��^�
�-�1|E)E$�O�Q(�A<�*Ydj��ȿ5@�M	�S�fH�N�{7[���?�O���ց�c?�K�\��S�B��V��}D��4g8��1���F0��#z��Ys����ޏk�K���T���[l���W.�D�|w�xk SM��`Z�$bO1#��f �*Ǚ�Z�I�锌�oQ�TQ�Ĝ��#j7�yL��M��Ò�	��:�͙K8�붥����&� 
w�����K�}t���ҥ6$Q���xt�:չ�&U�?\�	s�%c.��}�-{?6c�Yg*�������N���^��V9a��&�˨����"��^t���Q�D�kF�\^\jE�n��Z�����u
���o)��J1G֐Z\`��l�M��H4^�̰��>�v�^�����v i8Ȋ�!�"���?k��Ax>�� {M�vޓ������u �ʗA�t�;�s�wr�s�D�����R@:�CJ�?O����#��<c!$?�EPr"�R��s��}9O���3�St[@��`ةB�ݡ��!ee�W�T}Pm���%�ͦ�����.��	�A
"ɜ�8�v>�`w	b�n6-I�.`n������(v�l�*���k|}A��M��Vު��P����"4%[R.�p �`����>��[N �n�����<���m�8�M���0�ױ�����!Hݑ��<#���j"�
�K��?�8����������2.ˣ�h�����ͼ��3u�>,�,�\Q���`��o������BOBo�̥Tk�R��.n�N�/ef�+�-������"���?���'ly�&
>������H�?P�Չ��_�q�t4HE:k
�6<��v����85�=y�F]��]i	��i��\m�
�i�������1V�rn�d�U�87�i�EeY<�1��۽�����AE�t��^f�������N���U�g
p��4��_�5&�{0�mJ3�0o)ݹ�v�/<������1�c�m��;N�U�#�y}@H��6 ��.9�1}�����+��	�FU]S��y0��{��mS�ַ4 oy��h��O">��������Q��q�=B?N�[G�6N�(p�wɉL7�u�s&�0�)rQ���AY!b��ȒF�A�ۯ�Y�Ep��&���#�Sm����|�q���L�������! j��꿘B�Q,u��BŬd���A��s���<r:�N؀2x��,�U���,y&
�#�#_��]ГIVzیS�ގIZm�蒕�Nù���ʮ����84� �/J���Z�EKi�]�1�V�a7�Gk�w
�h�_�VM�� ��%)�<��� t�${f'�X�:��X!|>�V ϻ��D8E\�QA�M!vK��p�U2��}��c5�Nt�cIc���%j����o��@��az,��}���F9j2W�h�8�~�x!�x�N�wj_���h'B�M�=����
�p��G.1�\N���?���a�QԵ�}H#&��������D�1ݩٺ�i��ğX�������̐�o�oK���C���}5�.��Wj{�Vu���7䌱�"�����w(K���f�+��*�0]Y�t�(O�������>(���Ȗ�V�i�P���!2����ZV���:�� ���U&��q)u��I�G�;L�V��U���0;$2n�j���H��|5p	�zQ[��(:z���.AGN�v�,�E�?�In��Ç��t̷�疿9�u��0��D+b�������:}�M��)�o����SÙ��#�o��T���lFB!�'������Xco���,�/?�Cf��"8V�c�� ���aIx3CB���h0�L�O��]����k�-%�[�+z6�@��e��-�>�c����ȟҌ<��PH�t��j�V��j=qƱ@F}�ѿ��1TmT1Y���0r��-n�I)t@^���dǅ�}���b�Ld�<��^�x2�P:�P���#�&�+xB��f��EU����4�F3OZ�Y��pCu��v�#7�}�p�i|X�υi�9���+n�����A�y�Th�}p����ɐJ��S�x&Ƹ���HH�3F�kA�0ˑ%R��U��J��|�W�M�D;h������K ���������[rIU��1Ι��4�B�4�5�xl%�P\���+��ϋ��`�5R�mN��2���\e���̬�V�y��c������g�^UDs�^-��!<�ԡ��m���������NC�B�U��i������>��yQ���#��2򩘭������o���p��E��6�y(6�RU�͹}����U��cZ�b�VR⶜%��w����ڑ�q���t۳�7��Ϣ΢�.�nI�����4��Ŧc�w�}����	���.�Yn�ۭ��N{}���C>H��yy�� �T�l��M���i$,�eb��㌷���Oj�
���UO[�~Ŭ�Z����>G-�o�������&s�58�O�2�NSjh�~Rܭ$xdUi3�C���2����	�Wzcױ+1�@ĠLL9��z�q�T���;O����p&�wp�?�ؿ�ϣ�c�k�3���aDZ�cnb��l����������e���^-�`��T��x��GKL��K˸�+��׻���tD0��J�����O�wh��R�I~ב��`Y�%�T{�t���ꕾ��<��)�,�[̓��?O��.�(�*�n�Zhj����5x�JI���Z
����,0-D��Jm2
�X
I��/"(���w�_�(V�=�� �+��^�
��y������������`qX?��㗘��@�'M�ʇ^���$t;j��5�-����[6�%���(
�-3� ��-�"���9������#�{E��v�u����ϬLzظg�\%̙d5g6OL�5�E&�KKpZT�]�4���}�`�7���)m�@K�[�9a�2'�!���p��ԾY���<_�Se�5�,Ѯ�lCZϝzjn��ޞ�ϸM�����㭳o^�+F�ܗ:w@�L/�&sz�
C�	�P��i�D	��7�����`�����B'p�ϒ���,yrC�E����p�(6��}���-�l������4ݩ�F��>���N�v�hd�����ͱ�����i����H���O�zmIF�~�l��m�S+�^u��W[�U2A�?$��fC����{�P�_;����cI۝fV�N,�9/PB��
�'x���bEE��o����(:E�[3q*�4f�1���$�?���gv&|���h���h�D��uʠ���ޭ�7���F��~��@m֪
~�H׼b�ސ�D��]��˕ G��Y*���/s!����L��9./��k������׋���5DK�n�(l]�I�-�B�dl\	X����J�����t�|�Ȱ�W���=@���Udب��4'V�ڷ�~V���#W��_>����>�a�+��?�;����B�+CH�Y�Vn�N�f-�mc\�f���gM�&�u��kG!�!���I�M3ģ����{�� ��/�7��<R�utQ�v��f�^�?��p$�V�[	`1�g0!���nn����]�ON��ґ��]�.��&��������wtߐP�3(�F�&FߪhP#�<���1
6����^G9�?��T�Q�����������<�PM 9�Dt��%����b�;)Q��=�^yɈ���7�$+�u�p�Ԝ��6�����~�OI	����Z�Dͦ����l<���%��.�2l�:���Z�s�{�~U*�J4x���_-�<�:���a�
.?�N逌��Ը�٥��\�*Po���
砪?�Y�ҍQ�9��@n��z�Q�(*w�A��so�6h��rR��5} d�,�� �M�P�&��$('��}��*���W�'[��/�`HZ��"��2�?�a����X�����y3��y�ޗ��F�P��[��#Ͳ�y��ݪ}zs��F��}Y1��ȃ�B&v�g��5"����0����9-���A|1\��x�v#E�UT�£�ϴAǺ��΢Xb%Z�i�i�.��tZ����z^": �B�8�ƺ���i4��/Ȱ4��K�H�92��G�3�4�R�_�>T,{K�by4u���#��3����=4!���WR���R����_' �c�T�;6�פN���$�<>6��⸖&_̬2X�,��>�>�V��J�mt)�Ģ5��*li,���y`�/� I`Ai����p�u-��V4@��Ro�x7q���a ㌲5G��W��+.�n�yDx��S[��j'0+1?x3P����_ 03��w�]F=���A��e�_�z��Yw�D�p�wG�rF�m'}O�������8&��FԳ��tݵ]->ik�����e��̂�A���8*@�Ve�W������X;��\�!���/Q� ��;k���S�(�*�sN)�h���q��9(�j@��3�J�U���`��|1$��^8Op�*}�l��"�4䬡.f�aE�.>����)��}��ʠ����O��Ql��� &��ev��{U���sc+��g��6�S�m�pI�b�����e��i��{U`R�ױԛ
|�D���ro�g ���?�O*��g��߹�f;�o}p�8La|�ܚ>(��qH�3y�A�)�w'	��P5'���-��N�C��,G����a��a�_�h�C�wJ�
+7<�|��'�Z����:[Iѓ��T��m�1o'��^�sC����\�KՈo�S@ݾ�/�����hR��V�U���Cvn1w��W���n��<{q���泈��?R�h�w0vp�7���ܕ3e�嘤�۾�W���}��dfK�7}�Ǎ�����0~ĄZ5q�^�|gs\�M�ݽ�����ls�a��I�y1���m۪)l��n1�l���J��)�0Ɓ�5�D�y��=@ �a����|E�ߔ�Z)(6��/�vX�`��f�������k�9Fi
����66a�2#c�"��J�,�� EtQE&B��y�Eko�~.f<�RC�D��PK@Ct	�W�;1�L?4]R��>�๕��e�*���0q���hj�� �e�ap��OQ���(�^�ݕ�H��cF݃ҝ#��ףTC\Y��f�>�W��|����(>͔�kN���}x�|I��a��!���ʗ�����@kJ���:��4��j9�!�QY��&Y��x�8l�$ +�C�}�D��F�̸S�[�����G~b� ��� rH���G�����+V̸�ҞUk�mɮ��*ٍ;C����ԥ(��n�,����;�}g a�(��[FH���͞�,���d�}��K����;>���'��m���o��%Ŭ1�u[����r��^tm��_#��	�T-�ӌ�i�2�L�f��E#@0&�U�Y]�I����n���u8����ߎḈo�F�*�����rN�uN~�̛���I���_1��+m�E�X(ć��������M��-0C��@�@��'3Qy���i)�|����	�O+J��ʏ��wO��4��z�%�n���z�nwΦ�����g���y�����5��Ix�Ǭ��\�>�y�M"��O���sg�Rw�]AX`~6AJ޵>����s��	�@��/���X,��y�RDq3&�����]"P�� �� t\��\u�4��LΥ�AO��c6V�](L��&[Zq��U엛�.,� �}������z]T<��D�/ck�o���)_ g�?����c|�:�;���U~�}
/��er���ĵz���k�s��M砞K'=�'G�f�w��FU�.J��\�8�wf�oI�U�B�
y�]��S�p?Vq��ڒ9X�r�G��2�� �k8^��1��nQŝ��cB�T>]�v��'����	��1n��2k���-̱�T�N��Y���ȊW�HI� �AfR��!�2I*	�+��J�̈́�ɣH��0�G��1wH��qK�������r�_�~V��_�X�8)�Ozh7�y��Y���n��IK�[�<ydY���s~V��w�Ц�e��Ge��R�Y� �+©[�	_�ܨ�����bnG4oof,�>�a}���(�Üh`�o[0Jb�D�	� �b�*�Q���kn�G�B8<$;�ʸVk������F��a��Y��Q��2qD8M��3!m��x$�C��r���j�s[���(귢
,09G��p�l��\3�����Qb�?�l�x���Ki�2�aw�5�o��&lB�N6"�⻤��[QZ����]��}��w�cV��������� ����_�zy�1A��*�C��5hF�G��Ɋp(XY�3`�itS��!����ti[w�@
�$h�g���ԕ���[��h.^=����q��L����CjP;V ��+z��B݅�'�9
K�V���rw4�t����i�&N�B박uYh�Ŭ[�:!����x��U�s��B��:/�e��^�Ȟ�m T�&������0c�I/@^6Gj��c�Z�m�`鋦4A��#�Č�t�aE6��[�=B��?�'$6�3v������K�ț��YvL<{�$ �6PF�<R�%n	���T3
��.��g�XL�[t�gu����In�E�S����.�����@'�]c���fjf�n�}s`nԌ�P�Ģ�A���9������S\�;L4��<�Ɩ\�c����V�b��[c��� �ȷ^�H��]���rr_1��T��/S8p#w����P$ RfN*WX�b�J����#_�k@uה���U�m�{ШAf�0�"��c���j�Ъ?C1 m�c��['o���6�6�=��w����t�ԋ�n�2�H��Y��������������GbT�A�F	��
G�2N8����(e8��C#��_&�	�t'LV;g2� $�Y��=�Jwl��;�n����	x��7��O;�ugn�g>�]"�"g�8��� ��1����v�4���k@p&�G�6)�Z#$%[�=����>2�$��1<�*��w"A�M��פ>o�6��5ά��"��vY\3��aj���i2ĘR��?�ڇ�t\q�p��-q�J^�r�0)Pm'���e�݇�3D��\�/���其nR�L�~�G.^� ������Gcc�-߶{�[r���6�߮V��7̵| �����É���X$�:�
�-����{<%�2�0�:CV� ����0Æ�;���5?8��
�t�ԛ�h �\ƣ5~x�
��R�Kx*Sep��~�Mj��������X�-�/�K��^5"o�S Pv��اu��J_�v�B6k��|�@��&.=�����Ac�>�2�����G��!2��(�������=��@�WG���J��w����W%��d��4T�	5��ހ��$����9IiG"'@ۆ��M%N'#�������S��m,a	%Sh+F�����)$��*��	���/_V���?h��MH"j��u����_[�n�\l�"����-��<C���j�ۛ��������c��?�h�$�	pb��y
��'��A4�2���� �լ�\��`>v%����f�S��T�������y>2)f��L�f�\=��М�}��X:�S�0P�R|����i�B>Pe��~|I��пi�scI=�tA�)Z��_����C�6I�A�l]�f�ۚ����Xۓyا��O��K�	�l�0�f�~���^X$Ay�'����A��0�4)���$d���?ß�d=��h�x��z �N������s�]��H�?��o�� 5/�<*`zт{�Ȯ� 2R@����`��	�a�SR�&k��u'w�$N���d�̀����h��{gڷ�Ⱥr1[�Ņ=� �fB�)ҚG�=�����n���/R� ������?����G�7G���ݷ���'�R ���ivL^F�k��3��@�B���h7�9�4U7u�N�#���_˭�	�4��0�A�\�8?捆dg�R/1.�	D�y�;������tc<Y1D�;��K����̠�]y�������i�{�Ȏ�+,��IUe��E
�{Wo��o��/�z~��US�|�C'MJ@�	@rp�fh�b�Y{񇮝�UR n��t�-�PS��!Ѝ�I�!gi�R���0��?�����oDņL�f�%�;}�]i��z��	�h	����Wت�Q��gi�|��e"�Z}�:�0V��G�@�����[��H�BY��}C�=r����4���	?ru+�a^D	��%>Ewwv�yEd�Z4�� p��X.��Թ)��^L�֪�t�u�Xl�C#U��S3�Y/s,xU�c���N �+7E�z�D������䱙.�h��+��"ܒ��	��/N�f�ڡ.��1�@�ؘ|W���	Y�Y �V�=
-�̅� ��w�0=!�Ԃc7 �"�����C��8�r�"��l�@R��l Ĩ�h. ���V�{������
�^5w�&z�����vG{��3�5 ��G�+,�u��ݚ��eF8�7��o�E� ���.=����-+k'Ym\�v�K2-n�U?�_�t,�"�c�wl\w�8�	��w��ވO�?ga�C�h\tbb�\��yx�>���w܎�)��j�<��Tx���Z)	N��L��lY\�q�͙7vx�y"j���� 1��D�[A���&Q*s�	[�'�(%�SD9x��ڀ�Sޑ7O�?��z�����ګ��fA9P޿b�Jls=�9"1�����0m f/�2���N�utW�T�@���PcFW�-��AV�)oL��7�	���0�L?�]���7�A���ʯ�#���A���)�x����Ց�e��Z=�w��-�ku�� l�ɱ02�(�'�+A�|�o����÷�2:��Ai?{������1�26�k|���{����"X8k�#Wj��^b����I������=Y$6]�<�t�
xN�s~.��؋�-�&H\1��FVɀ�@��6;����j�#J�5�?�Dۨ�
��tG�sl(�Kh	��h�%v���h�V��u��k��9gA�W�	�:�*����dh���CNY=`�0��"�}�fc��y&i�s�e+<�
�я��豬���jt����fuT��W����yU��.P���'�&y��>6�m1'��C0r��+�@��^p��/��'�4k,|�� �h�0(+B����� U�`%�����tpP\��F�z�&���i�d�[����`%a6��k�8ҐH@r��o�Cֲj�P���h۪��y��ʢ�A\s��2;�&_~���GN[�jk����o�`��s@�hA6����M��#�ex\b�|���C~-�^�@��鄭� `��^]KK�=�[q|�H�9�i�͚��VaV�s+߫�O���&�������&��/� �Q|��ު�6�EB�"��"���W�����q}����K,׋��L�dJ՝Y�(/"�PZ�����Ϸ�v
fz.٥����ݣU����e���8��c�A^���)�1��kEG��ɶ �	�����[�+UD��l�eB� ��7e�=�H��ߜ"`��K�R)3�{�����$=z��'��=���>�ca��.꠶&��⧙J��S%�pys�i�����p�^����*y��S���1�%e�M"�0J��h�K}���Bx����|��.R�,��"�W��{r~�o��?�Ƀ�8�	��`�6+�R��!�I.����ba*�����Ps�z�@���AZ�R�{�R[��<J��
{��z�-�5��;c8���w���&B�;��w����ѱ;���겏�w����g�Pp�I�7��t>.aG�2�/�e_�����
-)�H4�-�:�R3N�iqV��3��U�Q^@�a")�r>�/�c�!Y	s��˃|=6"m�&ی�� ��� ���
���$\vs�||ϫ ��j�vg4�cQ�kq6�w���V��"�ěp��mS��Y�o[�\�j�)"o,�fb�4�h�͢�� ����������]�9�q�5���_L����h�)�g~{(�r���4��e��g�k�~쥂*�����GF��Y���H=����@L�G$i��hl�TH9P��	�	R��S��
�-/I%<����v��ȸ<X�\Mg��.���oF�v�t%\���ё}��%?��Gu���yB��!C�V���[NoV�mv/����L,dw�C1V$h);�c$�*E�qa�t�2[�Ųl�`����>h����ޙ���wE	�����S�O��~�nM���9��+:��{������Nav	�Xp1�6bU&t�hq]�>9�g�pQK�}�TkҋC΋��F�7P%���}�D\�Eϴ�Ri0��~R����F<�`�Y�t�
P��ֈ�P�MN�u�x�8!s}M�>@��<��-߅��?�]�����!�I�mh���$M����Uؠ(?�@�q�q��ÙL)�Z�Y����+S�)]K�p�KIyR-����eC���N�^M��G�\��4fcQp���[>�&�Ը=J����b�����
kN���� ���!��c
N#��W� �48�����銔��+�0�|�q����-CV"c�T�3^�WW<����ƾ�q���\4�jT���-����r�!ٟYj��i�H���I�q�5G����2X� ��g<�ˈ#�{Z� �[�ͯ��#[>
T|}�vYo� ���>�b5M
����*�D�,!OHHL�c97�u�3�V*,�~ l�<��;{���pb�R�Շ��:��1%�-0IUV�j��m��B��U��{j �G�b�L�r������ǿh��Tsgm�8U�3����"J��"4/A�.�/,T2��1�Q.�IL.��z0�Z�M��}5i�ͽ�T�Q�F�I�9w�*y&�n��O���K�첋K�N=h���)%�1�e�����=I��H��7�怗{�7s�tŬ�0F��,-����W�y|9�7��������w���BRu��������#(e���"�$��E�g�"�� 2D�#�aKA�È�aC4n�,�)?(v����j���!�DֻR��[��|��C	�-e2����\Q��`eܥfo��N����X��Y� @��_o�e�qg���U#`	���!�s$�-�ck�f�ʯ2R���.�{3>�����k��
"�+�	�^�p���5`̦�U�%��H$5��1|sA��nX������鏥kֻ^�{"	�&\�4Y��կ�p�ﴎ*5%��3�Q�]�o �qc�G��w�d��Գ��G�v�c�nC�ˀ��$�n�����'���I�\M������B���kuED�3�>m�/��_t��[��^��!b�=*�5x��p7�o�Ane��a��:x\?3���W��0��Fz2���R���X�SI�x�6O�� H3���$�b�uyd�
M];���Gf����#��5��
��g�O���!3?;���x�P���բ�/?Ǧ/���u�B�H��PPv+&�++�[w��\�2*��&ȶ�k�I
s��ENi��?0K��\� �be�͞�Y�(
آ��/(�XM&�s����r��^TI���ѷ��)>���(N�~9��KG�˝�F��!~�ա1a�����!�e���m�}"vV��?�"�v�������<�MFU6]%.���e.N`�+VPj
A�U���м�f�.$����ʊYw����W�r���X��`"t��Ŝ���h�OO��!F;6B�S|�6 �\
4�+'�W{^ݞ�0v}�X)�o+���8�B�^�w ~UX�oT�.CZO��O#
p��Ovي2��
�mǿ�$3��y/�hl���O�y|�|��%�?ZD^���Cd�X�FA@����po-����D�����κ[��X��6e� ���녢b�Z�g��y��c��+^�+r��\��u�@���r�#��S�f��f%�K����Ӂe�a��GC/������1�~
c���2�l�;&˓u̬�����"rj�V�-W����M�cVu��+�W� ���G��!P�md8k]�c/�WLP�4~�g�/a��0s���� 7a�Jo�E<!�W~�wgp�h`h�<���{net�Sf;c�=|7`�T~���a�+����x��/�+4O�2d�Cޟ�5��hv��Ͱ�r}9E�@{\|d>ة�ݑ��*�6u��:�ʼz7����&��:����0�뱿Q)I��њ�4*�j���*���ToG ���W=�_���غ6����eJY��8��6�k	k���	~�.�H�	HG�+�[�b1��[�i��a߽���wV��6#0j��V�;�لp���:9�4᧽ۨ��+��G�wI����I�� T�0@���|[����:����Ǧ���BKB	�O2V���Oe�$��X�R2�B���f��Z$1��%l���;�5s;��`ב��Hu�a@v�����Η��@
4ן��o�-��  �&��
p�͍ѵ��Mv����S����5�-^��A}@�e�@+�h�~�	�NūWP�������.Z�艹4%
��p;��H��`�kg�/�űjQI�EX���,��CT#�*���g�=�����N�W�����d��������'T)g�BBo:�KFW)�UK6L&�� ��s���el�A����5s� ��NSAHj��;mt�1�'��=w�OR��ԅ󎯩"�U	��UB��s'�S������R߻vQ��bx��^1{o�	��i�A?����ۨ�r����.�,�]I��5�>���Y�Վd�i�Q���AU���AK���Aמ�����,R�Gt�m��"a@�]�$�ߖ�G;�V�I�ؚ�q���6T@ĥ����n��Yo��[n���>�ǫ�ﳷ��ҳl��Ƿ��z�a�����,4l�:B.�f'b&�����'SI�,�[���8���"�b+2���A$�����'�ա\��4.�Tđ#u��W������܁��g�;,��"myH�)̓�y8r��D�z�9k��U��X���t��K���j\9(B�����8z��=�8�.uK6��1����|֖����"�U��,�����؃^�0��ժge�*��d#�ꓙ���#�GN�{�ԭ �)	ac�� w���l�pl���\�@�C�d�+�����欦@E]�y��_����DB�)b	�CƵ����AeU>ۆ"�c����=.��w�&6��\�k����i�?۟D�
��i%/}�/(S��*��Y�|i���r�R�/)�nIx����p�����̋皁 �p��B4f�����_���hS@�����9"k����h��[�`�U�m{\�G��[di�b#*t�+j��R�1v�j���`�⃧��Ӑ���f,�܉}PO��Y9л��w9�<�eJ�|z��NG>Z	�����X���-��&�� ��� �^?5�"�CM�d�z$�f��U�2:����,����6���%���=��qˑg���&;����j0�wҿ%����@_��AZI�D���8K����)�Y��O"������J`Hj�P�,�(j���� �b�J�7⟆F���ƣ13i�G?�#�o_�oX����82~?��P��:M?GPAyBS�.���f�����4�O�3�Y&޽v|�����dP%r�b�9�d�I�m�Nk�q7X�AV3�=����Cu�i���J��w�кL���ș��7c���Fǚ�E�����:��ն>�!a�D0�:�`��T�ӥ�L�K�[Qd��-~x�J��<)������]6�=�#�-*,�w��[v�A.}Σ�i3�]xb���Ș�d�32�I�����A7Z���N����R���JeT��	�'���T��_�($�C��BN�ii^��|�+���j�uѭ���'�Ua���Fġ����_6m��K��{�F|�G���I�ꑨ�����>�g��S���R,���|7st,�!�&F( rꗄŝ��-7�����pk�:�����pF#�@�K�s>Ϝ��.c�{�ѷ!e4bUj1�6X��>�*/�
�.����I��� i_*^�w�nx��Y,�}��^w��Z9G������}Y�l+��5�Ȯ��J�miX�gD�L��"rɤ�*jz�Mh�[�L蕊�Y^�I��=@��6u�w����y�e�WRgԟ�6�5�V�����N�<y�r�av$�Cֺ�Y�n�٦IfʼVK����S[�l���0���"|`����$�F�Gǜcg��h]*�{A1�JJ�)I6�	��̆�"ꑛ�y}���(�XV���ow� uG���O<B��fz�E�0FtJ#}<>�x?��)M%z>K��k�;;��n.b��ᆶH�!��~S^�����)g��c��_.D#0a�1�A|�Ϋ���'k*����C���}��3��7u!��(��<����P4�	so�%�+����/ײ$\J1���c����pE2�rJ3�;���3�P�����g~�`���ֱ�u�������qv(���d��T
t�̴�C����f��G��A�NH�cS�},�)s��M6J�Y9;�Bsz���^��A��(~�L�^Vm��*z���yؓ�ôt���vL�A\�8S�CS��K�wO j�o���q��Z���wBa"3	G�'�.7�������e��lU휳`����v�J�����"�-lʹ0䄉��},T���#(`G�x����0���d&�]Fx!�8Txi�v	5y_I�s�q�����ܙv��?$ !�C��m�o����������R:���h���Af��_Seh�+���S��"���g����껣b�ΒwCڣ�XU1�~r�I�s5�'Vtt8H��"@R�%U*�j�сV���`�*[?���\�
���Cl#p���V��"x�P��r�%�������j�E &u	��p����[P���#dϸ�/I)�`ŧ���C���t ^*�a�Ӵ%i�hn-#�آ��֭{d�HQ��V/{Bܹ��w����2G,�>������>��);�\�Z�Mi�*C(�A3�'㌯��W=
��3]�O�J�^��0O�0��mX���U��srg>�Go�Dφl�M>#r�xIST`	j����O�|�f�6�?�����TBˆ�j(�<n�)�J�/B�Bzc�{�P_z��iD��D
�A��!�\.j��]�\Im\���^V%]�<��s���y{�4��8�I ��*�0[�0����&}��"�f/��;ȗ�� �q��>�����"E�_}'�PN�Yi�9ڧ�*11j;��U�	5�E��\_D�#�`Q]����g�1�lc�de�6%��?�յ���������Vs�d]шd��*� ����Q����m�>�,A�y	�s�@�9�>�G��l��Yvh��l ��\Er��o+Fł����!�q��T�&��-Fz��,}x�^P86OR��TJ�\O�lb��]J��u��3V����5Q�fĴm"���`iSɉ��}$�8q�2���^s�;>��P\2��b)�GMcq[{��0����	��G{��=�#A�����D����hӵ^�7�����X��j�\��-v���|�F������n����o�<�PӜY���|�_��W)?����<��qW+�Џppk�GR[��|��wq��P�լ��XZ�k>�K_q�p�ǺcV���υ[�Φ��P��ʲ6tɭ��I�J��@�����`Q�8�b���&�b6vY���E�<Wϧ�U�8�U/$�Wo� Y���
˭{?��n�W+�Fہ��� R��}(վsܱT�3�m��	�n>������4���P`-�����h����k�^6�\��}^��|�7;"+ڜ
�<"V�/;^!u��m]�W��`K��+�O� d ��!h�_O��MN�v5�F2��DdI���'����9���g���E�����h0����d������0j+�R=q$O[PF|��V�~��r�-;��L��`�M�*��Z}bfЃ3gE� �dO����
��J�Z9nBdgdL���1��Ȃ�K�y9Q[)�+���3P2�A��`��h����f�F�������̲�F[�sHd%�M#G��{���,���k��'أ�*?G�7�E#9�}7JtxʑU�C����>����3���]a�?�S\��`��_n!4$Λ�z�:>J��1X{ E�>�VvW6c�*(���y��;�w�ɖ�p��id`�>3��:�^�S4��H����&�v��݄��?����*����$�`�+IxҠ�\7`���8醞�w}����k
��X}����l��M�i;���d�cH�����ଧ��,>������<~"d7�"��}x���Q�+��Y��LBO���9P��i�������_�7�bD��hKIU_u�U|����|&�9�̺�-Ն��T��O���sum�ኺ���v��y�q;��U�>!**����?W>�R�-��׳���z�ϙ���
9�J�ޭ�F)�;Y����=�y�.�������n`B�U�~�	۠<�	־.N�r�����"����jMFٹT�@��_b��As�xP�6�ke�3e�A]Ћ��hAKy+e�"���_dY��&��Ƥ����b_��~$���[��v-,!}�K�2S�5�-?�y9�0��%^�ݤ"�Ƌ�-�kk�}.t�^��f�j�q"�*�u��ȕe��R]��Eد(m�9����_�������ζݍ��2�t��4$�r�N��Ux� �8�x��!DP�P�u��Mŀ�gj��9v�qH[PF�f4@g���jC�ڮ��35�<��1:�#?~d�K�}1�ޜ�𭣪�Z�_�0j�a�z$��|��>�Ԥ48��)d�_��e��pd�%G�F�S�:��_���J7#�BV��j��mݞ]���;wL�la'貝��D��6V�2l����0��4�<��O�g�E^Cݖ����������)*z<���(h->c���� 4%������cA4����kC�f���¬��n���&���M����ߌ�45��;���4;�R$�{r�N�<L�v�(�b�w����K=�^Ud�8�u������?���6����p�R���l�ھ�]}(ddrZ�X���n����Z�����):m��q;Ծq�60�_ �di��o��%��7j�PI�_���o�Vg�N�^A��8����}���Eߝ�0蠤�ب��6`3]u,;��0�m���Ȑ��8L1�δ��!ю2���ZK�O�
]5�&M�L�=nl_p�q��i��}�o"rN !�(L��1����
�g�l�~���2;Lz����>!Z��j<;��LKަٌ�9�r�y)�T߹À�<#��OD�)𤔕�"�S]t�CoR׎6,�B��t�ٿ�M�3L���2�+��d�.�7�[���Dv�0Նd�-O����plI8�Eެx�,j��ɩ�J0��&8�r�4T�Wm�WJ!�#�_����.[����SZ���na���ܰ&��"�an
�%>����ĕ���A�*���h�`⽻Ζ�x���fjo��{�HyB�r�ϲ��8n���*m'6��w2��;�vŅ�$�A�#Ikqesլ���o���z���At�p���Z��~G�_���������H�	��w���(������<�"��-��#��a�f��ڱҽ�7�`_L1�k��d#�u�F���k)� f�5��E��v
������/ރO�o��d{��+T�|Kdd���\�9��G`S%�Z���bw�F��~�Z(��oA移+/8�٫4[� l����{Go]$�ϐd�D�P|����]�|� 8R\��D_����D'Ge��#w��T�� s�NQ��͵�����I �&B|�C��/�0��캔қ�e�Ɔ���?O���e�6{y/��@�w�or���HL=Z��X��7������C[n�R³n?4��6�H_߮�=#�P�����F�R��1J|=��36��5%���ȍ�`�'�cmR��'8�1|������br?V���n�J�R���~H�UO����0��5��̸�����ւK�JU:l�(Y�������	~;����[�����>�h�TX�7斓l۞B �*�Eh�r� u������E�C�4؀`��6Q�P��̓���kp}U��[
��k�����a�����̜��=��s̷ewA��{Ό���,�U~-���{L���T<i�A�Bx��ul��'0 Hz�M4�;V�9��6	(�
-�H�����	5�r���A��F���`�i=4G"ǃ��w^�$P���!��kZ>"��I���J!R���ވ���h���.j���5v�Tƽ�[�B�6�?&|aE��=+�!W*�ȭs��������{=�,��o��4)x
����]���|ܢ��7�w��A���E����!ݾ��~����M��xha?D�ou�L��p0*���	��s|
;\4y�T��L���isM�ߔ�mK�+�լ��s<�n�U�U��宙�!��d�d��)����m��'%�민���T���Z���;�ܷ��5�pӸ%�b7��9��.T&/7�Rq�ώ�Ȝ��c�a�"8���� g9bڲ��>�Z�STh-��tni�.X�fr��@��!HYCS����w3c��:H�B�K������A�^��8��AQ��
���f
��Q7*L���_w��a�bkř�Ѣ�����������(��JV�8OQ����|D�}S�5;��3.��HQ���ٜ�"�<�;�2(td�.���p_�{�*�e=�c������x�h�q���3l^+o�Lը�fN�y0�5��+�:iI��Rv�ٝ��D���C�&=F�Jb	c�-U�
N�o�e�����_���w����Ȇ��j/��ip	s�%=�O|1@�y0M�;$wy�c ������h�P·@L��ӡv�#Ŷ�窭-DLzһL	,��%���24L�ѥ;�C�?���o3�eRۅy���0ɢJu��f�+~�!g�U��D�#�,��vV��%O�#��6���?5�2Ȗ�;ʆ�-�ԏ�4٢Z�wr��|#�����a��pK6�K��p�����?��
6�+���}
�G��Q�ӭ�:��yb��6$,�����,�"W��Tv�۹�����iv�㺑����i\�����M���O�=RJ\j��f��X�����g�<���NZ���E�~��~y(L+L"#���2.i�����J���)��-�^�Q�VB��;����xȫ�$���j��R��<�������:����<��L<-�ň�@O�P��ӥuV�]�V��@QK�h:p1&�yuuєɎ�ݱe^:�{I�8[#o�Jd��o�������DJ������9�ߋ�-���(�uc���M�d���=�^b3v���'��C�q]�c��
"����fO�T��}�눐�MW�L�|�3G����t�,�Y�`�B���jA}�>�"�ou��nE�\���6��(��fM�()�������ͪw!AK�v��C�q �O�.���ip�(����$�܆d�#��w0�/ۀ�#��t�b\�8H�X.���1�f������^J�+,˘� ?��-+ �((�u��G�&-q�QnE���~lO��;���0\�4���8ݣ���&h��P��؞b���W�o�M+�_���D�[j�2��)�m:����k��k��zGN1�~2Q��γC�0$r]8LqM2�:sK
���5`��jP�@�ðvL:%���J;�U%7o��%X�/�A��Tx"�bnz��c�
����z��~�t#my�HC���X�|T��O�$6�˾�T��g��;�� ��&�\��LLq�cd^}ҤR����t�* ��H,�ح�Ż*�!������q�ފ��Gљ�f�["�s ��|��ͦk?�{�%��g�#c��P�)Ch{���w�s@��/�e�em	����s�܆�BUZ�pD-]z�	�l�n+��UU�3c[�<�<�`!�SG-^O"����j�^��h
Y� .`H�M0����9wgs$y|7J~ 4�����}����7V�-�gN�����>%�� �m�ն�X�b]�Y���_j%�+V��MyN�[�l[��_���c�	9$��r*GF3#Ԃ/��Rm^�/ �~)��X��� �E�:�G"�L|J�m���͹a.�`/a��B�|�E�:����������Zf{G0�c`��{��jV0©���k�(�n�J�M�a��!��T�=ɋ�q��5j�z��V��a��ӵR�ߘ���-;=JWta,���
��J��)*��M����|��Q���g}�W�Y|�"�������̗YE�:W���n�*J��/#��K�Vevq����
�kFd���~����Yϼ2 ���N�B�����ҁƝ��W&��fJs1ut|fȣ}y5���M�N�[s3cg?�8u��z��D�x�:뷑���(K��e�F�z����<�Y@�1A(��x$.p���'��??B��WGul���=}�JQ��dx)nDd�f�B\qy�9��RՃ��g�}	HA*�����h�:��5���ǝҨ~��gi3m�^�h&q<��7�3����N��7Y��~�ކ̙c'.
.�zJ��+4���.�H�Q�kiO(�19 *�h�~8�b���1�D/F��j-����a��q
%����=�o~��~�ٹе���J������#����$.xY
��q�E=���p  H�Ǒ�����ʡ�����W������$e����������02��v��*��GY�pb&�*y:���G������Bv�m��Wrϟ���b�p�d�#����BSh�`=!���2�O�|�����ON��RwUV�>"*ѱ`��Ydf��+��gыV�+�3\��Ƴy�������樍?1���b{8�tz����O6OI�x�R��Vk�ö�S�sdaQt��Dat~I�%��K��@ͼH�&�Y�3�������ژ[������ƚ]g��kEZ��O*܇�;N��B�4��ї�H"��6�F�Y2J�!M�?�G��J��4e<U�������A�={7�&߻6�ټ䤬L�z�t����(Y�{k�ŀ�پ�t�*��
�è��*�L*�h��7� ;�cw��(�&[�c�\��9e�uЂx�ma e4U+������Ϛ�����q��i�^������#���]�[!�����jRE2ŇFl{)��S��c��Ϊ8$�;�KMOF��06`t�����|[�eiT��;��H�g��|����f��J���r� ���$La>3j����㗫�Pa��ȱ�b��
;3��(?Hrwh�Q�]B�]c�f͵~�M��j|w�Ȱ�N���CY"�J��hA\�j�>J߶fᕲ���2��吼�a��c@Kh\�O��c��Y�tЃ�����(�rR�:���G�h����t��8�*�[��?��M���C?Ek�
���5��-��l3��V����%����
�r��v��t*�����'Ɋ�k�v<z���F��k����h������&%Uq���%�Į��@��I��痸'v���g���[�و��f�4�h���,�"l��ǋK�=�.h��	������#���p<[�g�j�r�b��ֶջ��8#\D���MD��.�_��8��Y\�A0p��)��E��[��$�H�+z9{^˫�є?c�	┍-b9�&~�i�9��s�%�.�a�W��A�V��i�]�*�'0�������[���j��<��ϣ�G^�_��Z��E���h�^��ۡ]��#����6�g���m3*HY�
���+k��lJĒ|;���b��T��x>�����N:�d�����b�ԭN}����ȫl�,�f���q��RL���+Ô\���%.�4�6�7I��r"
� '@����g�n��?��D�pWY2fī	�jot'F�����$|�vDM2R�D)g-�N�۸���	�z�!p�2���eƝ�@� .���
���E�Җ��n���
�#P�>(#����+b�ϛ��"�IlI��v{��#��jӆm>���-\��K�v���ژ�>u����ܖoY�ݩw�My#�_6�����JC�y&�*���}�����Ƅ�5���R>ɱ9��t{��r��2�G߱Ro�<��?�������>�kȊ�����|�K�z�+����h��Y���rCI5����-M����;T� D�����A+ܩ*uO�S�rbU�� |�.��
�W���]>3���P�y�YF�UZZV��������h�p}�#�U��_4bt�n�������Q�)�+��֬w��j�"�)9b���RA�oJ�O�fp�?3.��m���QH9Pĺ�;���H�|GI[�N�-@���ϑ�%�Cof�����S�w����-6l(n�%�]�M�����cG������,�cDt����c$e>�d~��Q,�q�奅��yB%��d���4꩏�J^��������ߎ���/WX����h2mY���P��{�9�k��I�C�âT��7���2�#u�3���%GEժ��ǍCy6B��i�J%��Q4�s�h��D:�D�`��E�P/�ʌ�O�U:�"r$��O��5 \��'.�C�m�{!����2��l�NL�%%|<��8J�m�0Ԗ1U�(;/��Ps��$f|�(F%~Te���Jy���U%�k�.^��ć@;��L�)���.�\����M~���-+��P��@�yg�_((Ru/����#߲�����?�W�2�8�IOO�_2��	8���C�f�ЅV�����޺�K�h���m���͂!���Ba��;6~:�Ϝ�jɿfs������A���#��wZ����>֎��W��-z]�z�8�f���1N�Ûr�����OM��ن��fYbo��1~�7s�Φ>�vQ���i����@W�<a�|.7�e�[����p��ԏ@�p�H�B���p-��|��h;�0l��������6"�ilv*�7:(P.鞦O����ߖ};�Ğ�W�7fFAx�[w��[8T���}^�)X���0�]nNKi2GN[��q�nA��ט�R��T�|�$-�x��6�zU�od;��{��G	��o��I�NB��U���A�s��m��0c��!	��̈́�l���i�A�6��!V��>i��&�{x��'etu��%�i�����zj��C�CY��{elO��t��eh�d�p�6ӥ�,)^�h���'�0|�J�
~�4��*�;.��d���� ֲ��]�ϱ�C���H#f9��'�/; %�U������tX�`&K��:-+�LĿvɫfIb�Os�̸Z_�'6=H�'������C��&��sB�\�S��t6\ISߔb\�e�a���F�ߜ�*}Dq!�}=Ǫ2�'v*��o�|��H�+�͝�RZ�T�����`-�I����'Ωg{�b�0V$�wZ�p3��	�����]"Cs�@�N�o�T��g6�����(��lW��������?Ū=j?��&P��%kmF�� I�%���8w5)f
z%��5u��PB'wěj�����@%h=a>m�1��^,��%Z�@8ٜ"�sh7��ГmU"n����d�� )��_�\7�A�iSL��[O������3I���xf���4�ʸ��.�>���J���;�g#�Tԛ��?}���Y��i�0y��Kw4�ی��@��S"؀�g70� ?��0\j�P���uf�2V���:�F��R��	�3�qS���!3m���[�S���=.p�P7Qq�͕m_�(e�ٳ��C?hy����E~]������>|��U8�����4R�nq���󵥄��r�x�̊��_x�EHtA��+T�קc�4�֗'f��t7�^��9t��I�Wi!UAi�-<�O�ôk{")�
g���@�L&O^�u��~��j�'t��������*3��ͬ�,�=3��+!�I;=3��;����nM�;��E6���2iw���Z;��,S����Qg>�X�s�X�k�ɿ<s��Z@M�I.�����:h��C��`�g�*Z1�����]�~s��@���Hm�B6�f�����au�O�heK������1go[�V�\SSq� -���;�T<�Č=Y���{%���%pd�ؤ>�H|f�T��2��GT|����. ��0����>��۲�DT���P���rO�wq�lm�O�߬�#�����p�'�B�$G��#���x��_�˔<ާoOaг�GX(�sT�-�
�9���%X�7_�xD�d�q���/�_��볋�*�]�Ոf�`��{!듙&uE�A��`�jR����=�¥P)FȏZ����_r���}T�q�o-( ۿݱʦm��.�]�
Igk��Lp{�S�����|�ӢzK��w�8W��3��	"��C�_BL�Pᇵk��A�|c���o���e�ϪA�=��IJ�@�q�Vۤ�+I�R�R#�0�E6=�K|4��!����j���l���n�����:�K`��9E6h}�6���6l{����l��ǐ]qh�`_Ϳ�̥�c����wb��w�������n�������ݡ_�#�I�]p�
P��������L|�)�^�%�id��ήG���7|;�����PK��T���Z��dΥ"2:�����/��z�0��oL4Ll��4|8}T�Q�D�j0T����x2�`����2��#dO@�wC�f5�����]����00���+���.a��=i��w�V`h�zP��'��[pWp��O ]��5�n�?���J��\�>���z�=��7v�9�Z��ZF�X5#���T�&�Y�	�RY[�nk�DH�$Q�� ?�}O�?\j��:b3�����]([yV���~�,��<�<n��b�����Մ�7$��\ܑ0�OQ���4Fd���h������ш��S^N�kOz.�4b���ȸb����� �lc��Q_Ne�ʎ�`�)�6���j�a�)4�5�,�P�G:�d9��|��r�����fU�7pxOg/��� �lM1n����]��2�dz�;�[Ĝ��J����>�V>@����J�g��A���^ ���<�SҶp'*CHZm��^h��棙5B�%����<�n`�cbb�8���?���V�ԇ�F��V%�o�D܌ ��M�U�Q�S�c0�7U��3v��&~1�_s˨E���D��ǻ�gG���nȜ�~�X��7�[�rÿ�{Ot�x�ˌRx�h�gG4{!4c�Yq�!��{�T��3l4$�`Mo�)�M������;o��0�I���)�e�LeD@C��0�N�aA����xr�Jb�T��WS�Ͷ�I=
=Y�槔����F/�A��/�A-��7L�A@���m�{�-W��}�˛��r�_�"P�.�7>_ʏ�*���C�������n�	�P �`N�1��K��uV/�*FwƷ�Sk�[���#��`v,x݌5�J�7���:���z����jE��9C��&���(�ɄqH�$��8k$K>s_>,ߪ�WH�=�����XyaҤ.^
���?���{��7�U9�T�-|(ީ�9�ZO�B4	�+�Ͼ�&��R0��ƴmN��w�b�������V)c�i�eJ��7����C\�M{��j�ܕ4<p�p���zcf.�j�?�M�Z`�������ؔa�,�]O��|IZ�'���12X�^Pr�,������k6(���QS�,�P���M�o��3c��,��tCl[���P�5B߶�u�sO��3���!�T��|�h"9�C�����t@ѹ7h߳⚃��FG������=���K_���TE�`%�����~��Xy2|	z�&Ke�L���\��b�{�[],o��dR��ǹ6@��,{M�[������]�
jE�#V�Y��:)z���N���d��w~�'���:
�*������VgOB������9 ⇓U1�n����I��;,��p�/!�V��p��p_}��Ij��eY��l��r���Y���|��oQ|@�������!7W޲Fm1�	8gۢF0�1�w���{�ȩ?s%���� �A)��I�C��G�����4���Gʁ�?�8kK���b`���r���\�^���C�m�M��]�b�@63l�:�J�*eܲX./�BPd�����btu��PV�����ݰ8%+2Ȥ��9w�ƃdL95�$P@����.�Z���v�tt��l%���
-ߊy�yRt!�l ��$У7-�m���h�l�gQxq9��Z�E��YL�uD��9���V�'�-H��&�>iV��,��W�-�F�x��;_x��`�[���V���8BWe[�6�߇U���PM�,{�3r�x�o�Y��{�?��(|��(�>�3?j���7`������01V���.TN5)��0����"�W
|� mqV��2v�Dk�CīI3X�O{�-e!'k����RDz�!��ѡ�C�_`3���V��l�[������N,y��q�w���0�J�,b;�Vͧ8�3J0}g��+Y�Q�?���v}�9��5u{Ik��;��m��a��+B��ܮ �-������!>=m�0)��C'ց��\ރ���5�`��� Ҟ���)�n�~nI-~�k�Bz f��`21�������+4&�[� I��T�;m߭2�p.65c|{٧�^�VD�b���a!���(t�l'd%�+Σ�v�#.�ܤJ<۫���Œ��$��%�`�Kb��XńdI~i؏��7p,gcR�
u,R[Io�~�����颅 xZ�ٔ�>ka���ݔ�2��L���(���fsq)���w���X�j	<GT U�mٍ��/
���Y���e�Gc�m��W�vV��q.ߥ��u�����>6����8;���՛��+7ڡ.|��Ec��z�,�b�[�t�:H��K;<����=�0��j�8O���������vg?Х�u�}vM��A��-,�� �4�=�e�����rV���:-��h|��(y=QpK5�K`�m�.�OVt�{�L֦�[�+�ۮ����+SƯ����������P��hև_	�S�c>o��B^\�ĞQk��b�m6�¡��jʞ]b�<��b�� ��/�[�w�����	@\T���(�^�ޟJ0{Q�bbE��%���n_�mBZFOά*�Rv��K;������ڏ|%���B>����E�����Ǔz��,��b���oV��������J�{�t2h�.�5K��,�ۮ�����6������/�Y��%�h����7��������Oc�8)�:�pƙR��b��c}��-�B� �W�Oi�I�W�)�ҫ�W�h��M�[7)VDF��_����J�D9�.h��\�C���|is�H܉��� )$$Ybx����OQ�U��)�ofA��kZL�4YS�чq-ũ�(��7�Yy�B�$�����_d76Q.d4Tݍ$��qBI.�蟭��W�=�>Բ������#�<�aT^��;���$�EA�ƀ/M��7��w�	N�-I��=�<&<�ٗ9w�8��5O��Cv�d(tԑ��8i��B]]?�a�7�X���yMT�q���h�!=��y�9>���M9�~a���5��]p�+l�
�:����,���K6.c�Jd1�Bt�i1kS���l4;�G;�����l�De��F?\�F��/6��Oxв6��h�a6�~�XV䁐g<r6<�Mާ��_�3������Z���,d����.2����p^�b���֍�/ܞ�4	"��S�Fء�? ��	2����_���1��Y�� _�|��*='�s���8�5a��55��i���,���%2/u��<����[�ޖ��N�b�ʷ��2�,�L���U��ѵ�͌��l��܍�(0xu?J��iVe�Mn�}�����<�H=����ߚ=dO '�.��FO�ɒ|�H9D�=�`ʉ���XW�*�F�#�7�j�����	XT$V�r
��k�L 5�,�A��4}eu�H�
�D���3=��t�}�M��+�?E��';Y�\��^ه��5;���$a8Os�.��qSQTm ɚ�O$ns���a��RU^ i 6
��5���"�O�L�
�p5��C�����l��X�p��-vL�U��i�^�C�tr�8>�@E���k+��Q�:��W#7�A|RwN̶�� �8�ݶLm���w7U�?)Z����_��I��� Ɩe��ɝ�eJ�FoN
1�G"oi&�jO;�9�7KF��@�^���ʬ&�Y�.�1�ظ������k�Y�( šO��*�9U`$6g��:�x���J�ue�a��8�'�2b [�e��guSʗ�UĖq$���)Q�Q�����FD�����(FH �aG�S�z"N���S�5~z���0�	*����rF�G�+M�Eag'�#	 ����-u�'�@rw�`��b�����1�eg�c��˓~\Oly�i��1W���;�R�J`���e���Y��[�u���<b>[�����X�0��薈���L7�����Vwh�hW�ɪ{3��)�.MU�A9�$@U ���ć�����C�@&����{���sJ��Mh��C�2����kaq��k�Vf�hV�Hh)�H|�"�Mt�����/9Gߵ��z�n7/�6�\:�b$D��ڶ`˒�\_:Ղ�Ѩ��
>�������?\L��-��Qӑܾ�k{'�H������l@.�	��	�W*��;-`3����!O��>���J��O�q�6�\��
�y�<�L�7f^d��Mr���ߏi"Om�:.�E��<�����$��Y�����F��������p���:�,0�������w( y*����#僓~�����*K0A�KQ��h.���ƄRn�! �_��$c����*C��Pᐐ�b��ŷǩF��C�p�l)JSOζ""�L�D�**/J�	��I�9&��ԑ�o�m���MU�)�)N�f����CL�&ni2B߅��W�lr����[��r����:v�!$�9U-�
`�q��-��T]�t�[#	���� ��iB�f�Qϙ�@]�&j��Vs����Ń&Ϣ.�N߃�g�9�d>��,�k��e#��kj`5�Y��0�ѓ�W�m,���2݈}��U}@
׸�`�,_kׂ.��4s���?�/�y�$�������j;��ee�7Y9 ,��!��ޢ*��Pz�Հ,vZ�-����^�����}���7/����-r�����f$=Tus�Q�>"��4�|�⏵�=c�_(a�V��-��C[h%�#3J��m��	�(�&%(�"N�ӥZK,B�G��O
����ѷ#�4$3�nxE)���7��/Z����4,��J�2�x�	�u�RQ�C�9V˕�v����
����E*c͚�i�x~��yp��:V�-el�r�Pq�⩏z�C�c�� �w�NЕ6�K���4��֜�iZ�����p	�Ik�ӄ�R�zv79�v�fow��r�6F�0�\�RQ�p>�[�`�����E�r������d�X�YB����'������3��w�������^��O;z���Āfdژ�A�����4/Q�h@=<g>�x��K@�8:�y!�G�Ǌ�/`����g{�ǭ�Vc��~�I���8xv۰�н�c�RƩ�@)�~\\���*��o��r�_8����FuU���ܑt����U�s ��$z潍�
�Y�(������Tm����$��z�vefm]�u�Tr�kS���#r�d�]�Ob����S���~I�v��1�A����z�Deך�2�j;XbH��z��l%��ۿ^U�)���Ԁ4�����y���8����w���8�^��������{5N�I_ۊ���L���/�,�HA8q.C���$j�a�e팖=\�ᴘ�!`��w��[�c%�}H�d�[���c��(O�ƅ�(� �#��7qoD��mnS�y�#԰ ��?�4^�z'H i�JM�A�����@�J��;t��o���| ��M�8,�����M�/|����Iy䏏�F$<
���FO��U'��;f�ę���hmC3�f�O�W�%<je'Cn�l�:o5�X��G��������:1zy�#@�0���������~غ�M�og���p<�h
�&��.ڃ-[���jIcu����R+uQ�\n�X�'n/�zY�;���D��e��8.�~�'���%*����l-i$_zd����A4|%H����m�f��&;yF��R��A�&�^e�CE�,H|�(�u��w����
�+��Cҁ³Y�珬Uq8h�P�SN�S���W�1;պ���&�Tu�0G��H�{tZ�85�i��!��7d����ml���}tߙ3���yy�I�r��CK�\>�׺eOk ��Zd���ze��< �F��d\{�����}A
��J2΀����'���T��E�K�!�]�͗�xw̭L'�%y^W`d#�܊����FҢ�(m<�v�E�*,�)��;15�W枷h�/<�lh��"��8�͐�b
��ͽ۱p�J�JH[���+ dէ��*#)�Ab7PN���(&ο��$�Sax�{���6����HC��}�)%Zg�\H��FMz8ߞ~�&�.Q`J<� �F�/��[���h�(����.��� �ޡ�VԄ��7���{m/���}$h��oY�M�����K4찍wPR���6q���37�?{�Rm�����{l�q�&P��;a5!o��y)���咗 ������}م�z�^�Ő�dpIe��A&y~q���b�5Rn#�,�"A�ԕ��"p�@z��8y.����緮�|?��F��[C���{'��.L�?L>��}�y���2k� q���㘛�Ĩ�v�*�1�������M��a��$~/H-�vxP��6�m֐	p|	l����V�ٓ�j��ZS%�$�S�g���C�K}�o��#�e���;�N���C���+���W���AU�="�߆��$���0�$��p-'Ϩ$��*�ͨ�h��z >(iy=v"� ^Tq�������v�}�A��ӝπ�Eťn�O�n¶u&Z+5'�CL��LGz2�+U�%�_��ה�M���(HM�Yp���҂0������;ͧu����+(RK�Qa�K�BG�˓ŧ�3UQ�7 �΃�˗��а� 0:��UH@B����"���D����p!�5�y�ʫ��f܉jn���o'�q���M� �k
���ӺL�[Y��Y民r��QhqMC57= ��O�
ք����͡Q�� /dl1"��!{_��*²�J���R��(��+�$��b����4TM�{�=��u��&�O8��>�1
Y�q���_�N�rn�՘�yY+ݢ�G�D���{��53�%���A��e�������yӐ,��Ǜ���tuWt�S�>�VQ��t�����`�`ަ��{M7�}�Y���΢{��Uפ���S�Wс%]����f#|�>H�' 5�괼lS�T� ER����e�����&�d���U�'�p�^z$��qS�A����O�E�B�r�]�O�,�"w���s�[�',��s��5O���·/�����u^߸B0:Uy��.�Uk-/T�+��ɕƷS*tK����l��"#r&�Aa���رsb|���CI=�ډ-X��n�2w7Ae۩ɮ��S"���+��J�	<t��h�i�L�j'�����ǝ�y��k@#��������X��r�5��lE����)�I�"?G��OWHX�Ŭ8�@Ʌ��5��p���Bcm(��_i�ƛ?��E���X:<���Zp�\��s�k��w�F��]M���t��dF�V���x6&�G޶��ڳQӃ�zLq2S޽�����W�Q�5ݳ�-H�(h�O�?��W]�;� (/h��^N\B� ��j�hm�ܛ�m O+l�,��f�1�ʡ��r�O}���y.���6�)y�r���������/�1F��\U�k�e@�w/E;x�AW��ߎ�:^� o�Q0u��ܶ�dW̳���=�C�1_��w�[��ᆑ0�C�����{kꚅ`<�s���ڏE2]6��V�`�k�-S �x2��܅���k��)�ЉH�(+%�*$�0�t�:^!Q씣�1���0��=2�H��:�����cfv�1%��Hڲ���:!��k,AG�)�!�v�ON�R�3˱�id	��Ӟ+����!�n&�1�]q��M-w��gÓ֕4VH;�w-j
:��zc��37v��즶��DZ�"�l�Ӿ�F�p;��4P�t��;��Pɇ�:�������l��oc_�3I4m"�]'vne⇨�*����X���6�����VM���	���̾dX��"���������U���*KK�y���OQ.�{�@ �F?t��v��t�����S��+��s�l�VM�����6����0�^�������q�,�Lx����N\�|&�!�m��к&o��FK�����նXn��,�n���1f(�l�tW3¼�5����Ԭ�>ڏ��!
x�<�OR�zM�v�hf��Olk��g�i�Σ�اi=���=ݰ�{���
��F�)}���U!�&q�d��/ �u�5l�{�\�MBݎ�
aj&�~�_�{����j@���hϊw��H����~��ۥ��������q�@g�TE�=������*��N�H��-�s�v�L�5Z����x����`�$�S9�o}ְ뻷\�Yyx��/��j�z���6�4���=6~������"�ن�Q� 2Yfv׮L2)y�\ZZPUg��h�
E�_A�|�Z��l��ؼ_ȝ"���IJVr�>m�֣�k�X=��R����"���&���Q�^S�B����j��W���C~	��u6�Y�Dj�5qO�SQ��v&�-�kޓdn�O��
%*���W���&���|{0;fsM]�5�"����]ܥ�M�����#Z[��S�?�������������ؖ,���Њ��2[��uv'��δū�>��>^����6ﯩr��.7UWC��X����v�8��]�0���v���)Z�x�X��/L�T�G�|�GpGH�������?2=Mد/^+�'n��o��YT�y-{�	�kd��E!k	Xh��/��dp_(D�/�����;�ѴV�0��P�s��0㬋��O��~�
�v�I�t��
D�[��� ֿ�����֊
	1�� ��T��>����\%�{�j�_���88/y��L�Wv��
0n6#�#P9aZS^�k�I��BH*|�[	 ��%��S�Vޡ������գ�8]�Q�C��~���bXgo�q�&KN>��Pv��&��DQU{l*�"�vf�s��}{�6�i"dM�#�uid:�*&���ތ���^ӆ���c1a��pE��������::ߑ���VY.R�o9��k<*�6{�<+��n�L;p��ߥ
>*��rŉ�=�+���L9'}� ��p� �d:��M���&y�x��5X)�ƅ�p�ݡ"����?�D�Ҝ|{��*��z3���<�o��ً�d#6�H�T���o �}�O{ /�6��e����|��IZ�:"�z��uN�n~�y����8���%��*g��4lTn�P�H�F-��o
l_l*-��*��cڳ�	��C=��_+�8�I��Ӿ,�6�p��RQ]�?���h�����5�L@}֞n54.""�ڏ5�*��4��Oq�22��q���{n�kw�7Y�K���(�1-/<�dzD�h_�J�i��L��|Wk#�'�����?ޅ��x[�b	��g�b���U&�:Q��B� �w���6U��e�,b@)+�����s�_dg�AD`�/Bs�N�y\t�	���;�u�g3�ɍ�b�y�6���+9�_k�>�9�;��DX@�����]~���F
-�%�|��Τ���Q��_G��G����{SB��C�� 죂t�DaU�����<��*6AZvN#7m��gu�s�}�_�.ո+�R-�P�/eJ�fK�]��ΘGvF����a�����p;��9�y��/&Gy�􏋆��m���ZOg���w�C&d��zh#�:E_���-�@���ռ�f<�S�a�Us�8�t6��q�`#�(@���\h��R��4��#��X�[G��8��ʕ�WdO\F\J^�%�.x$o�a��^�fψ��W�2C	"��mgO�č�0��\�/5��^h
�B��X{ī|�M���
%~n���U5��;EU�X{�Ucߎ�|=�������-�u�L��l�~Z��Br����u'���Ɇ��	�ɘM�*��HUh�Ca�|d�����E��� �W�~��0�ө6�*�cL�(v�;����� �b��, ��j��(=h�5O��w�N���S��+�V�x�"	� ��Ei�cd�ܙ�  ��.�ihg{�������kvR�z�n1��c�U'��P���X�����}�*z��dӺ�Z5���5��أVt*ᑟ�|{+��(]M�C9jxK�x~YY<�6ם�t��o6��w�VD�[���)�l%ͮ떫b��� ��9o�L �){C�G-�{�0a pv@`BQ��L_��Kҥ�#�Ib�8d��^:�4���SOd��"Nz�I'�y#�cYVI�W���Eῳc���A<-a��,��hx����ta,+��柜�"�t����3>�J�ܐ����q�d����qqtr�s�E:�U�i=�z�P) 所>;�z�W)@m'�{�w�ƭxv�������!=R�\n[����Z�	b�`�b�N&����bM�����B~@t��cwE��4rz�y�ll��S���93����$�>�;Z����"%>���=L�3 ��r0�O� S�������<��B�
��D+\Q�&��a��Ǐ߈��4����?9�
3��h���k_�xFE���ad�����ʌ�G{Wn��xK������p0����-�"z���-���*�4p�P�fE�����-F��ϥ�B����xlC�,��Iyx&~��
��.qT�%̗��TA��O0���ٶ:�s�YB�F3&�[�xMߤL�fԻ�	�u��+l��f�;+Ŀt�/�����l�D?ia�
+�����?d���q��v�g�uì܅t���~'u�L�>��w[��=����7�R����C��;_�P���C�d�G��+A&S���vVX��u�o��3��A���xu��+���_�r�"ܙŉ1f�$1iݓ�ȕ�1R(�211W~�' ���a����b��J��cw�Ĳ�\��A����배��s���5�̐WC���6q�W;��*�����zUaf��t+�1��p��&;k:��ӊ9��:��Ѽc�wBX`mMz�g��3Z>v�XwS.o�_$3˪�j�	m%�Ά���!���VF����ǬrQA|�ک��C=r��jo�X��l��k���4e#o.x��z�=�v'��GP1J	�~�X�t#�y=	�����^�Dz�J�l`BԿY���7w�z4 Ċ{;Ӿ��Sk��*�:*�nOqȍ!���̋?KKcb0�W<M�p=������"�sv��i0T�yK�YE��򑐅��ne8�RT�R������Zl<OK)^M�k����3	6%T!vk��(F��{k��$��H���b� ,ɪ0��,}[D��95�l\�?������#k-aBt����L���fH�/1K�����v<�Cf�]ܱ�Ͳ�W}S��Q��Dos>�k'd'����B�IZ����3�{��3�d.���=ufX���o���Q�v����Fc>`ꑿo��2�ӏX�|f�!���"U	ư��+Y��c��ti{q�r�.�aB�o'P�0
L=���t�;g�!���u���;�v����E:��{Ƹ���MwnҼ	޼97ǧ]�v��!g�Cݟ�8WS4G8Y��_�d�a��6?��zG�A}�D�.�l���tFL�Y%����f�}ǫ��`-4��
���%��7��>�D]��:\|T_I���	躃��0�wr"jg\#^��.��</�M4�	�i[�e����8����a��VRP*�Q�f�;��\w��E���ߦ��-"��	���S���NX�@%�2�؜p���L�R��F|ܜ@&�e�����Rb��0�w��\�� ��)�^�u5o�0}.��Ѿ(}Rz �Fn�WDH^ǲ���c���	��q)���Vy�wB���L�E1l10��v�N�v��L��Z��c�f��z���p�Fq�%��b	�p�p
�����Y��%���f���xL�h�Y|Fש'υ�'jK�$4����ep��H��;�?�i�����.����f,,:q}�����5�s�I�Ky�xI�Ds����;���W�n����𲲹Q�h�(�N���Xۣ�$* ����Ht�@ȡ�
��zB��/;��[�ذ�C}��Ϟ[�:�:��P�O����9���ű�����Q����x��������^�k���rhtҚ
�r��|�A#�3!�7��'��7c~��+�5�c�A]�='��Vݪ���i������+>BWs�6�)�>�@�@cH�qY-�T�3� ����@��M���J9t�ߌ��^�e�{��ُ���U9�XJb����8pm�\��9��=�k���nS��d���y|�/�߭��p���^�"�[*PN�H�A*!&ޢ�� ��\QT�2E��p4λ|�g�S>v]���.T�o>�>]���T�b~�-��*�9T��Ԗj8�0�~�����!��S�����5t����­���$<Xy�!t�踸���E&Z[C�[|e#LV%�_J��*1�?�H go"u/����)(k�	�Ef�/�]�˛�Ȍ��a���	@p��HN�Q���k!���/�7��~{������-�<�&m�A�-�}��Mr�4���8�KB7�����2�.�O
��X�䳏�Kt��˱7�s�4O��n��@�+�^R�10[��Wm����u��\��9���jw� 7�Ϳ��i������跶u�b�3�1?��n*�)�wi�t8����w���&LS��x! �1��o��R�v7��hk�w��PEC�sҪ>L�tv�.�6۬��RVnF�k8Ƴ��m�PLIT�cDőq�N�!u��V4�YZ��,��m.�6�I7�_rM��Ϡy�없���m���r7�3��4tY[�����X�ua�`D*=�U�*g@$�R�^���u����5i���:���T�(�9��;3�.ͬ�s���@@�et	�B1�+u$�z*��X('��p�[�&���0SD�j!ס��ޢ5��������c
�t�r��}�BY��iQ�������Yn>s�3�%$\��w�'�>Uf�:�S)�$?%�խ{,aK��P�@� ��E	���<�}�F�)��5�>R٩�	�ϟ�R�^J�> ��,���PT���ٛ3��=�v��3�팡d��fF����0�	W(^G�)�򀑗H��Meg�KUm�שt�)͚GK��R��A�0g�."��~�x�iu䛉X��Nټǡ�7'�)&�fV��
�]*l�[�j�ٓ��G0{�2���`ȕ�)�\�$I��bύ��_�c�q@b'S�8D���`d������g�������'�"��ǈ��|r%���b|%�U���^���{+>��,�&�&����ڑ6a�N�//�D_���g�X��E�{ �j��a�A����m}wO�c���O�;+ǆs�Pp�6�h�*+�g߯�έ�V7�uM��<^��R�x/YI	T;��3)|ީ��Rc<L��h\ڭ�B�)�p�t��Y|�z�L-��ϟ�5�=�>�W7(	=˼�P�D�V%�5�h	]U���k��J������ܜ��%"aT_�Ȗ�����T���>o�iq�N�܂�^jO�C��������=Ej��6���d�!)�UgL^_n������d`Q�Bbc!A݇ �;�b�Ԩ6�=��oz����1�+1���_1�O݉��p&ޢ�i�o����8^�M���A�	/o��C����J��vq��3΀�Bv斑�d��L������4w�~_`�8>ުz�R��@b-q��n�#�f�A�3��!'V@�w���=7�pN>�2���&EJ,�I���`4	�PI�{p��������
2�~(��+:Ja�dGf�9��ؤ�
*�>��%|�_����ͨ�-��qdץd����@H�}��}%�,���kA�)��ڶ�E�M ]�@;��\�F��^�|D�٢��وw�9���t[�0\��LP�GZ'�N3y�v���`��X�Xsmc��}�*g,2��2��eS�ޤ�#�?�}l'��@OV4:p=}]��,r����I�9�������I����W�Ky�dY~`��)�t+��6)����D�JUC�E�+S�=��Ⱦ� ����^a�� H~@�k��q�:PH���+�e���XF
�Z?�]B�E�파t~��M�G��_��1���pS��3m:��G�6��s���7��6�*}�b�-���H9�V����?��$)���Xe��pX����޹����7��C^Z��!����rK?�
������~�*���}	�)��L�����ΊR9e�z
��,Y�ipX(�
<DHS��h�o�M4�pڇwJ4����qc�����9C9h�,�n%W�J0�Arp ���)���d�D�=�O�B��po�~.H���� �6:�J1�s^bU�7_X�W(�	ՍQl�A$�-qz;l���HG��шb��7�a.���m�U�8�����Pf$t٩E�K�Q�#>P���f���b���VE59��9u�}�Ե3��:	6�݊u�I�,�~�,�,��f����hi��fᓀ�M�!�0c��H�f�v{qh�A����S�W�����F��oX����Z�P1��E���Ri�f��%�>=J,����=qR[zc�l�F/�РV���U�qK�myr��=
ݝ��5�<3�Zs��8&�B�}D9���%�����ͪq�ѵu/�ԓ��D�1�)��Ghy݊V�� �Y����R��6�y���8���S2����N���vb��4J ¯�χ��`G�⨴�ގ�B}_���rqy�C�pE�nN��Yԛ3߷�k4���d���UM�^��.�7�B�UX�ݒ���;��tQ�a*�י|�Χ|Er�;%��=����?�����A�{���+�[�/��&M��������Ѳ�1
D:`]�4ր��^���r볺����_w�A��|h�[����<D�(��]A����'��ۀG���
&zo��}�������G��!��DXB+:\�H�7̽pd�?��O&����6Ĕ1mMH�O��B	[�O�1;ӦCV�U��k3��ذ� ~���[�t_>),Z�q�F�̖���7e����D-��Œ��V��w�i��C����J9oF�%I��p*R�����1�l�NN.���I�cy�4��$_h����M�C?wi��u�V"X���d�����n+����qU)�x)������ Um�;�se�H�e��oE5�!/T�_ĎM�H~'��gaet#۠�%�_��!R=0�@��[�/�8�Y�H�$��o��I��MV����B)<�tF^i���,�mꉱ�^�8u�Hg�>Y�%y�40��թEkYBD����sGx�s]�~NEم3_�	6w�ߠ(E��ܫ��^>]aQ�D*�?�� �\�>6�g'�.A���;8fz7�Ni��X��z|���p=�������W�V�K�#iL�{u,��7-s"��̯6�0z$9cr^���=u`"o_T7؃;���#
Ŧ.�w�\����WhfKԩ�9��n�"EJ�خ��C��uR�a �Ie`�Fp��o��ۋ��Q���mn�������%"3��%}�����JZ��w��d�VS�Ff8r��;�8�CZ$ �����z�x:��l�zo�qL�0���rH���jfF�R�҄��jζ��I����.wzA��roc�v�7��K[��=7'��P�'�R����S�}�>43$��i�> gd�%6!���8���a~邀�L
�`��� ;9-�ب),]�i�1�L%�¤�ً{q�����*�T��}��2�V(�،V�u\O�+s��u<������BQ'��!���H�O8@���,
H�t]�l�6���p�����U�b�9PIڒ��'iT��aΆ�����9.�����J�YywW�����:ni'{�f�f�>���p�	(�n�azZie�^����$�U2%�Z���)M,�E�~J�a�>�U���3m�I&u���	��b��ٶ�q�h��[/�oִ"�qҏ���~2���QTy
1q$0�<&5�Ē4#'q@��xH1rջ"V��HIἃ\��+��1]�/�� �r`�t[�%�ۢ���|-�.q����>�}���5� b�t�mq��J)��Z^�s|�F�@síi�?�1�C��š27��~ҧ�g_�,���T�H|�l0�hm &�*��~��V{�`�����~��N���/,7��E���`	�@0�}���S8GI1#�(��I0a3��,�x����\��vs2�^#d�"�s����K|9�z�Z���X���!d�o���D�!EeԖ�;JR�g��B�P.��i_c����E�s՟>T�7��d��V
�O~3n�9X���_����f��e?o���y!( ��r>�,��>����Gb��&/ ��6$�*9���Zg�`��]^T�>.P�Q"fO�W*7S~8`v5�,�"ăi�'�2.p&�-��*��?�#*S
\ǠJ*�>�ݕ��1�[t���4 ���-��4�!"s�M�*�\��Z���uC&k�!���gn%��{�|@ ��1��r�9��B�˩#��=�|ݭcrGZ]��zb��j+W�Z��Q�Y"����x�y���d�C�w���D�~S2��b�z�cp�yMz��C�����||�!���H�c�|�� ��5�~����e��L����E�������)�G:qï��(�2R�VA{������5��[|�
�*ʈK,�[��O�֭���7&ݙ 5ͼ�ְ-dv ���~�P�*70m�Tc��Q� t	l���P����f �N�z�<%[��u
fq��s}���t��ȇ-���?V�6� -H�w�ڭz�'�֡`*zsC�CHgnEg����$�렾�`| �.ą������B��*��������<'2����=�`m;����Ϳ�3;��LF�Q
�7��֘�=�K��DH>Cb�V_��A��N��'��V�"� �pu'0�Q(G�.�D�w�%>#-̳��� 	K�����9yY�U�<��D���Év��j�
a��izv��	��/���!�o��h!)v["@���H5C���������8���X>���!����{<�_�4�-����s*��S&U�EA,)���2��h�^\������R��4$8�s8VͲ3J7
�Mi���X�E��w��ɒI�јeH=�,�D���Z�W��cȭ�9��<�u���V���%�B��SŞ��S�C�,?����qF-��2�@<�ڕ��8仧�fET�����HX#���w��nx@0�n�Ana�3
�r!LgȓG�u�_ZC=�*�걉����n6�����j��n�m�$qz˸-���j$����c嬷��LF�p���'
�o�c�,���
���_���#���)���NS(K�4rtf�(ށ�Ha���K�Qw�f�pF��d�vY��X��470���4�ɀ"@%he�yTv�ïY����_���}б4#��(N�wU랠����#֥Z��T��-N�	:�m�e�\�m����}&%�~�d��#yx.����
��\�x匕2��L�-T�b�7��I���Z�O搲8��S�CM�+ub>�p ƞ�"v��(}1 _�>>1����\[�c#ő�k�3G��'�=��[Mɖu���(�V�T蹩r�
*:I&#;xr�t`s�ϛ�F�E����A��9e��U���6�����r���!��ZI�:ڋ`�fh*��p+,t/��K�O䁔h1ŊA��>m������/������o@V՚2�WP�h2�����Ag�����~���U���_���0��9��N�d�6H���,;��~��&�&*p���)ο��QRs}�:��C��.�7"�i�K����ō�R�a���5f33[�o�/�87��qD6_�,-K�u�����͑Z�fT� !� ��I���R^��=����R>�7�">|�E��a�{�.�<w6�PA����&��D�ꍘ���
�Anep�j"_)�2~��RW:[:6�! ��E����!E&.�J���r�=&�^=��$!�ù���N�� 4��b�)����h�5��H+������~��Uf+�s8Bc��#d�%пT��Б�ԑH����_¯ϫ��qsj���]��;�k�[�lify�nZ��\���z ��H�Q�]�v/��Epr���qK��b)/�*�n���/��CxP���M}R�D��t�@�}_�g6�Q�Z��'�·�8w��-�����5v�w��g[��@<惸�jE'V�����b�W�2� E���f����#�4�N�'K�G7�'�����W�W血��7=\;������,�#���$5h��z�c����ur��jA��y��
�͑:~���b$.pƺ
� �(��7��
r�I6�<I��Cɟ�A���j�@�:�<�
��Q�|��1�Gʖ���R3xV����ף���
a ���Z�I^�E�N��pP)�|�aBO�G�.�������r���!ٸ�m�r�l�_��8�t�z̳��d��.�R�[�%S�a���6A%�X#yd�z��A-���l�>������&y8��[�?�������*�tm�˽q��
ڮV��N�O{M��1���2k�zj� �Z��Ud)�8��e���8��c�� ���f�"��cW*[~w���Mʵ�c��J,���C�Y�Z`�ԩQJ|w���Vl4��	��A��E�Q��br�{>r:��ɓ�>�!?�eq[�ѷg�%E� #B3�	�|H1	�J	>�V���b���d �1��Jń�kQ��	��D@E/jOf��AW�Wa,��)]؄ˊo]�?���j��\!�h�*y�w�����P���c���A���g	��A?Z�>
��-߈�7���D��p�`��L,�Ƴ��|}T��)|f
�L�5�`1+H��Eǭ�4��h�vȊ�q~!\�(M��lJ�����{�j�6���KP�bwy��5�%\�e��M�ߠ~�8�I,���?Լ�,���[��ad7@�
�*��ߚ���oo4�����\���acm�U4�����-4�WI(�tma��#��HGE�;��-m����d[�zM	�9/� �WƢ#I�� �l�~"nI�\�P��b[LE�	�u�`��9���}����8�β�!��%S���:mo��x��z �r�� +���3[Kx����Ļ�;-�l����Aх3����ؕ�鷐�3?��{B��3��Fф�#2��?��Ă��}n4��|A�^�I����bh ׻���.H/�J=Ȕ9�ald
_C��m#�/���,*�F���w�i�ƿ �B����={0��:�6)s޹#|�u?�|^�:�f7�^�*W�֌�3���̐ͳ���,�0����Վ���cZvn[/������tu+�x��	繵Ю�[���>z���)���&�7&���DT�"��׆Ti��)����f����%�WɣH�?�;�˘�w��0qEǧY'�"[�NΜY�t��(7 b�k;k*+���AK6��~�]_����K��N����}���O�T����=�r��E��4�]<Χ5�q`P���W$�禼��a�~�i�br�pUzօ��x����{K ��逸��՝>t�̋�m�p�z���Z��dv�4L�_/��m;�����;� ,��)�n6 ȉ�!�;r >4�'���N2�I�"{�3n{����+v# G��nlE%`UG�����4Sj󠘀�x<��MxX�´�ՈW�(O�����G�O`���G:]ˍ���)��� �+�V$BSgM2��7�xp�#��[��v[��U��U�1�s�ڎ���(��iw��>�\��n��[�B����9]p���vgBZ'M�W���DCC��d�C�a����������[,y!c� p?Ll�jmkܷ�$[��u��̐�r�o8�����0�\AYUg��ش�"�+���v7��L.�S#��I����{KJ	��s�FIo�(�� �Kf��g�7-��T����p��k��闱�DF2�Ɔ�Ӳ��D�)հ�E���7��ʯ ������ؖ�F��e%����n%4�NQȜ��v��6֧���,%���ا[sT�a�{�3@������F5U��N�|�Ɲ���H�޺�O`�x�9�^<�������������� |�qSZ�f<�����q�a�7nftĢ����C�K�vIPg�6���1xU�q)KG��,�
�2��lz��$��=r$^&(	�@��� _T�9�%���������l2�<����o���!V��ǝ��Lq�[�w�IOzL�f��˔�Ν���sq��9��)����o]�����Y��;�{���c|�[�l��ӚK�	����a��2�g�M]�t�������z���`��g���!��w+B��w�׺�����?�}CjqL��Y2DJ�E���8-/[�g![���aE��s�L��3M#x��H*y)G��(�Gܖ(�9��!����K��<YF�8^^u�p,.�u������	_�@VU|-�#�L-.�qS�-Qp��)�~-2\;�vQ��t��+Ѱ>�d?��q�=�l�4�����9�;R1��U>�8��Ƀ��$��nzV�Ր���ϻ3t�1z|��7,Q�U��V�c��o�e: �#���)��%�����R�:��"U���A�������Yh�`�ƴ�c������H��;i�k��,�Y�1�*����[�VTr��;r���|�E��>�lnx]rR��&=���*�lV�*�ċ���JZkZ�	Lן���;����tTi��_I}{�&AIF�M$
^����p�z3ۖ�v/��ߑ<X���c�����"ÞHb�Zk��wf l��؏�)��߲�W╼Ks�H _�yK������%�N�P�Y�ߢ�c��p����8��5M��=�"h����ӷ}+s���;K=J�+P�����K޳P!U��2�S�/*L�*�O��gF����{ɴ�bi���@�A�����Y��'������$O��aǹK�Taq4�s�� .@���vE��N�v+~��D��P>�4��R�]?lx{!�����f����PE�=�ΉAB�����/+�j��E0۶�,�(h�8�[<y�Tr�������u�^ '�ho�x�5�=.��jD�����dW��&H3�ZH����=�>������_r"��K�@��������/�ǧ8͙�7Þ�7ˢs�m�O�I���^!�ݺ�(/�RSGz��GP���m4��s"�������L����Le�e|T��9$֢�@=�>R���G���#-8x�gX&�-�	��;ޱ���d*�"��;��*`F��\ :�Ax�dbE@�����s�F�Y�y������ �+qd��ǋdߘ��<w��z	m�,=$��
��=ƿ�v�	��CR���n\Cx�:W�;�5�����*��p2����	����(�zn�
i
�w�R�Gz<�����5p��vf���'�n�:O��]WPp@ ���v��h�p�3tȄh��OW�ό_M�����P�Z��q�mZNM���w���W�Dr��TQω�^ �k�6�+T��$�V-�EE����V�Z��rLjI��yG���#֏B�',�����)�u_�e��@�I"g��%�	��Wh;I����o#�)Q�Y]B��aMJdMK�ןL���w�3�0i{��U�����z�k��DEn����5=)�A�Z�D<y�ar'-��n.��/wf"sd��	��d{+U�D+���
@��p7��ଆ~Ό��lr.�}�NY`�}{�rBe�go�S�Ȼ1]8�>(�D�w:!F�u�:��,(���I�(}��Z������ �Dr��"=�Z6h)Y!Õ�kB���*/7O	���8�����}p�E�U�&�1E�l �e�ꉓg�=dZw�Q�=�{�7�m[�����t�?�5_l����V[�iU)�s���ٴ��\V��=�f�^��X���+����������k�7��`�.�l���C��b����'!/ �|����i�б5����kK�d+���au}2l��� �N㰕:�4���U~�@��.�}�<d0(�Ķ^Xu�g���2o���	u*�w�0ϣ�ah r���"�<8��� ����Ҧ4��G��W�$-ͤ"��3�:b����0>f`#7��"�F��q����CI����Z�k�vy�(0���%K2��EM��s���"���0JQR;o@)���2�d�Z	0?p �b�U$n���l�?�þX��,F��H�Û��$(�߀��478g�s(o��Z�����fgǄ�i�ɽ��x2Ք�/���`ޫ�ϲ̘�nd��q*�M���#R���ܙ�>��V`>xL�J�Ѯ��@�~���˹bN�}3'$��"�?��'*]�MP��ZIO��$tM���dΩ$"ߞ��̕i0[ta֒c�\��]������c���f��8�r�L��{�o���K<x�G�,E�o f�c^��T5�]�,�]�o��?OdN����9�[�f��83��'�%�J?a#�!7�ޝ_S��?=�VW3C��d�S�z*���0>�^�U���o��JA���~�V?yen�t��6OR¿?���2��P���&�����*s�ʦ ���J�B$lᅋ�T�H��Ēz�Ru��v�akg�JԢ�o�����#�)�� �7+�_}�,�!�E��Rݲj��o����c���5�<m�̛ƛz�e�sA�9w+k�쬄vk&�\��������YUG��x(=!��$oWU�Rz��^*���F�I�2E���!pʰ-�Եn�(�4�A���\4�N����%л��Fs@`�dQ/i�����A�YJ�W��_�T�Z�'��"�N<��~�@_�R�gO�9?�j� ~�,8і���>���Z�;����p�R�zОlm�ҿ�,��Y�u/���~*��]6ȱH�ɧ�x��VB���2�/�������'��4,�7��ܴ+��H�M����&�4\W�����B�	�2-r���&�8\�wk�<	HU8$Em�t���ʴ *-}��.GƸ~�b��5�1�j�c��]9�|�iCF#y�4��k���*`����/��!=�E\s���X��r4�#�b�� �?�:�\��m��3�e��B��.|qN���ð���_�b=�U���ݸ����w
���/.���<s�&���{����M�n��}�Pun9%�Ϡt��g.�Պ�y͢0�b�Y}�3E���lz�+�'QKl	8���ܹ�����8N�8WS߱=x�� �%�	X�Le�[�W>Wό�dj�PŨAJjY�n�~�\�`2g/����<b�e�#{�)����t����b/,"���4	B\f
��4+�#�	�_~	�E[f�EeL^gҏ Z%��Մ5���83�v���P�
��,\��T����d�j�|�6���*cr�z�J�V��c2�ӵ%�R��g����C�w	�șW�O=#sZ�_�8Qx�|��s��_�w��	}��b8��&H�I�r۸��P�K�����1��:]�S��z���0���H�����<_p��3������^�����$<JW��+%��L?���.!���
w�{$A��rήр������Մ�~S��KBh�m�����IK���%��yDϛ�闯�/�9qA�ho�Z�DB���r�"�����¸�pwg�}j�O�I�|�"�=�Z�e��e�NbQ�L�\��b	���*�׮�+-�)!()|�������v���0C�h���p+�;�0�_ֵ���៶q�!!�q��Bsj�1�9rG��[��+�͍���+�zV`���D�R��TC����/�b=T6���j��-��ed�z�u�X!� ��6��+m�Yȧ�JYXPXE�x��/�g5������:0( �Pk2�ɧ�Sܗ�(�f���pU�����eSh�E3CO!�̔�����GQ^n��jA�k��ɻ��%' �t4�?�����:R�H��ѓWIw�V���{/���$8u7�S\�	b,]D�Z��"ꏐ�r]��e����I��'��#��&�DMAh����S�oN����̦����|{��a^}���76{��cl!΅�,+��Y�V ���I����%���f#*��"tn��7|��{M2�2 �����] p+D�_pj{s�i�+����E�
�&�"1����,~� Dbߧ�Ǔ��Ը��~-�(�u@O@7&��A&R�I� �>[x�V�Zz/ �cSd����"��x��ﴳ�T��_~�vE�֒3�S�t�P.�����tp�I�&\�e�"�a�7��g�0`�6��������kƕ��7��	l1��6��-Lsv+�06��s u�h����f
�ľ�C� �.ɰ�V�,��7@� _��y!���� �f�R��JG�<q)�,%�~J`� ��f�X���Ľ�����-Aݣ�I.��y�GR��q�e�+�����V.'�f��^y���o�n/6s�Lo.�DfN��X���v�V��ъe%��N��0����~�|���_�����r���:����e3Ϯ��o����l0|�Äj�KM���e{WE��ӺH%���Cd,��������&؊��p\�������&4q�4-@o&1Id@^_��]b��������J�I�IH�8�*�{���%7��_@RG���za9��>�<Ô[޽��D^U��ƥ�����ՅI���L1��v��)u�kNr��jv�xd)w�p��|S}�n��Iq��$��:��|]6d/Q�ڸ8#�����I75x7=(�E�g�� ������˳�����f"'-��sɝ�\�b��w&�L��1�,/8A�ź.$b�B��F��.�EXE�e���Q:���Z��~n!aZ�[�sr���)G���)��e�H�W�
3�T7�+,�ۜaT9E�ϥ�]�hT���h�y��@��cy�;s�U���Y-����/�,�`�7$��K��Ы{��_���+
�f����s=�1V��m���ߚ�V�	+Dgx���/���~���J�M=8π۹̓Z��w�����飜����?SK;`aFqczUd��V�N�݃�{%�(�G����8��xG����G`֠2���l{%3Ӂak�`��t��o������8�?B%Խ�1dR�#2�9|���/}ba�u��d���`M�ʪ �d�#��X�����f[k�� Ѥ�bbr{M�t!#Q>2be���k�s䘭�:$����wi\_�0o��ڸ��� \��՚���u���$�
�S����,��^e/m�0���c
y�%�riZ�mþ�����ɸqI�!S�HF�0*�#�	�����p����	�B& V�v��?�</��>N�<���o��j�hM\e0z�r~����	d�,�4��T�Ec��լ)��� 7��.}*G���Л����S� K�@��PQ m��9sب���T���ny�R�4{H�ͦ�eʸ�8��?�^��N��'$o	yclV��ӡ�0��/�)㷅7̡ �U�ח|J5��'�|p��T����0���G%�]�U��~O^�����(��D/�5���A���Q�1J�q{&�Ul��n���[Q���8v�.}Qs���V��O������$p�s�;\���FrЄ��������:��gYnR7u���^7��e�2�b%,dｩwZ!S{�$j"��ъ�d-y���n_�� }��<��hI����������v���D�v\���;
|Z��C+���$)��¥��[�#@�6��[�wQ<!ؑ���Z2��'��_���L��&N�90�b��<d�O��ٙ�hz���J��l��*��+,����a�Җ,����w��]����G���8
��w�މ��o�����
�08��/r�2��Ə�4����1v�����O&v`��(�	� ����6�R2�va1y�]��*(b�^ ix�����X�nq?M���_�W�U�j���tr�4[�>)�!�1��ˀ�?��
Ej��6�
'5m��AY�pw��+6$!V]3{����%X�;@��'�"���� {)�Ta�4�U�Ƅ�U QH�6����Jw
�.��p�)U&���*wX�������#JH��y-�N[H�h�1����kb%���nEU�e�B�`�t�C�{d}�#�mrCR��M`�j�u��r����ٓ�[��;�ݳ�b �}���~�ޠ���%��LL2�63v:6���F�}g��s>'l�UѤr�L9�?����bTu�Q��ҽe����U�:�����P����]��v�87�h\��6�q5��,�.j�O�x/6GPΓ����#$��`�*\Y'�U��T��3A\{��,�@҇+����PN7k����5��6�JbQ!�zI����"c}3�����Y�� E�%���O��Pʹ���d��yzaN�E�Q∸w��
 �!U[�UR"�6�YܵR
�hw;�L	ٖܺ5����u����n�|[Zh*��]ڸeQ�ڟ�J s�<����lQ�_��5�^Zeځ���I�;ٸ@���=q��6y�*a�"��퐰��xf�E��~�"������_��ĩFh��`jP�*�a�Gl,Z��%��
R4 /��RG���lg�D4��+���D�6���G��k�>�7��\B���D.��۔*��q��װii�&n�0�"�g�?��(r)����s3��5+�8sX�v*���M�7b2��&Mvb5�!k����J>x�&�PX��w�ڀj���DA!Z)����a�9�Hs�R��n�\��ū3��<�v?�(r\j�@!�<��D(�N��FB��ݩ(B��n�6W�x.�����hKc����u�ذ�&dG3�#��)�j���[zi�����@�[%D-�}t:&���G�X	By����ܦ��kq�m���Π�8/�����ސ��Z����vr��^F��J �&B/�аE02�����ėҠ]��5r�=�6K�p��ڿQ��@��G��UMVv��)�k���" a�Z���K]�\�1�x3�f�,=t&eX@ �^�]切P8V��iG��YYX�"$aձ)��(�8j5�}�vXo^����(��s������<q^w��\���6���gՠƑ�,�>$�ި3�Sdb�L\]4H�\�r�5�N.dA���5f����oI��ᲶU0~<���� �� ��3K�!J��19ㆆ��1`���k��-�^'9�<����!x�v1�)ے�C,I��/��Y�=lO��6�l��S��3���NU>�ܷ�&T��kOI �|��7�'�<�T��W�`4(G�5���+V.ȤO�"�<��lPԧ��H����I�Z��n��ʴ@����Ƶ:��P�|cv9���~���q3wnY	r3e���F���>�ʵ�Q�3,��ҍ��� �_@YX$7�	s��ǋ�o�}c 2�wY�EK��sG*��~����4Ҫ2�+mb�+��z�.l�+��@f��IK8�ߴ����9�v��լ|>~[�^���_�l�(�)qg�C�<��9��@]l���˼c�m�5���9ڒU2)�����֤��d;ˈ.E(&J��0�ѕ�b���L�[�A���d�	��R��[H���h[�S���V6�R)��yC�l�l���{����U��Yh)t�p������w�(�̨@�� 4���Y�Tf����� #
�����y��1��
\Zu�۔�r¿&M_&5���ŉȋ�4�����x*�e���c�*�k�c��炝xz�-F��t����V�j�5s�h����O!���,t�(�aU�ǂ	�x�Bx�ߜ�W��+ݖ5bdE&�^� �Sn!:C�.j�'
�AJ:V���f}u׵�"�C��A���Oߓ��a�}�o� �ia��Sl��6�O*�x����sH��4�i/��9�L
9�e���S������|Ք��_O��t,ܣ���1�2$V[��1p"uP��{ʹiGm���Ĕ���i7�>E���p倕�;Qo���z�#��B��-g=-������V�6c���,i�Pd0���c2�E��� �>���$����2�h�4j�$�}������b�I��1��#���v��.y�Zi*��qe�.8i}���4&�5mo[Q	�d�'GVk�!/JD=f�&��`h	�y ���-F��)���s�sH�q	�=�bJ7y�q���6%�\����vM� -]�z��tF�Z2�խ�m>?����W�[Q{{NA�)��I�����uqӉ�P��K褍���O��c�����j�8�u��!�FJӰ�C.�&�#��JA��6Q��A��f2�`xG� �C!�I	8W��w�޴p�F�.����#z����yGs�+��B�?��Y��F��*T'�ZK���+KK�`�.A$������B#�*�3��2��ve�{���c�ؖ��$6���h�/
�z���<	/��`<]6����:�>a�x�x!F9�+��λЌvrDu��s7���gMN��i���2��:�`!7����@4Ԧ�%<�_�,X�äK1A���D���dt��������Zdxh �--�Nd��S�h�t!��t=��%9�D�X�V�f2�6�	b�2�v؜eA�V������Fm泳��Ʈi�����ܜ� Z�y"�,R:3�S�����K�IB��Ê�-XX���&wӵm��0�g�.Ψr�luں�gZݤ0��Q���Q��o6sG	���2���Qr�x�N71}_��yJ��'�D��A�ח�x�^"*�4$��܋A�$����I���s	�䥗�k˙{�e�>&�V'%���EY}>p��|�(��c��vwB"�<͐���8�&�.�!����.<���7�ǅ%[�<1�<��"cdQ1�`m�u�T��O���܋<	 �su�.���@�%Үtja���R��l�Ū��Af�PC��b� �B��8WB�M8:L4wq6Mw�Q�u�J*��۸�p.3�ʋ�I3�C=��R�aLEw~>,�1��օ�?�ɷ��?&xG^�H,.��4	}R� �ћE<��-�`���+��^�9���L�&Dѿ���t�t������;�M�K`5����έ㈚�R?�3���L����F�ߠ�+b����z���G�^�jA��?�*����?�,�Ѥ��b��aZ����L�U��r�	.1�2�//z�/��&�r����:�^��A�����N���&}I"�4�8�o�#:օfhJcKJH�Px&w��&�=c]�CF�*���@��id�$��Ԣ�`��WJ�(����~���� �"���}JSm��QM�d��S �ˉpk'H\�B���Si�`��,!ٗ+����6$���m��"}��8$�%�]��Ԫu ��S0�B�/@Vh���1lP耝� � #<��mp��w,�ر-�!^���e@@8
u"��ln
�R$O�:k=��$���?K�S��o�	��J��M�H��x�"�m�;�C�&��f�U��/���ӳ�t�Է���K�,�s��Y�#�:RS�m����J�e8j7��Q5'B���$p���a�@���� �vי����3�ރO���[,��"[: �V#Ry�0h ��Eo�!O!�3�0���D���Nk&3b@���B�A�^
m��ox��j�~����Q��]$�N�~/Qg�ԫއw�����5���N���AΪѩ�'+w�a���r�]o]�E�Gp}fȡ5����)lTax�����K@�Yb��o![��N��lV��g(&r��RpP��4c��_L��L�3���MI@�D���MB�bD�S�[��w�	�z�>OާT� �L[�ʠik�N[��DIc~\Ⱦ����I.f���F�����y|�<)4!䙅^�������X�_����/�;����$$��!�~���G��r�{��fo<G70u�<��h����������?G�B$	��K����%�6��L�~����4�����./r����V�N �6�o`�3D��D-�F�k�u˯���|fm\Z󭾆bt&;n�+:���	���IP�H/2s�섒���x�������+��=��ǳ��(� ��~7��ϭ�E�
����K-�4w38�\����cL>L�h�j!C��� k[��]'^"|l~���i���)�aK��Me�=��
������l��3��E;�ޗ���1���-�?\�!��y�w���d���m�S����W�aՆ�<
 ��6�_��g�Օ��}��Ks�I�6���7���[�'��M���zR��9�rǸP�Mb6�Ѵ�r�p��W� #���wY06K�m���Ա���PK�|[~6H�|�7x��s܃_3��&�'X9�T(MZ^�?���`���+���*}.fN���������"�ﮞ�+x7Rm��À�r[g�<u�^�L_HЗ1����{rK�\6�bRr���]���M�m�V�Tb��&�Sܧz����RG^I������bU������8��W/�c�x��H�KP����#=�нs�crS��m>�=���{jW��y�P��(�ۻ�!��u�I�g�]�XG$@��{�k��O�g�U��\M]���f�ڵ�\h�,,*o�2a)���xgl�ܻI��X�܅�����T���}�r��r9��@�!�-b����	C�:��E�K\#w��m
�"xl��(����y�����Z��V�#!)���-�� �Ƒ]!�\�-#\ƪJR`�Qrdۘ�k����8 j���ŷ�xH�pt0]9������~�A2�g��r��E�t���&ܚΓ��$��4+�d�P��B�����?�2D��r���P�{w?"�O��_.�ڝ�&�-[��ܥ�ޜ������I����B0�۲��K�k[˙�D���I
�����B�p��Br�$0��f�.�|���s��3��mfiH��u&u����Z5Y.����17�[��E+���*ho�v�sD��j�٫�<�vQY�,B������{����L�����c`�U�����D̚�A���+��~���MI����B�	���דּ*�.���@@� �r�T�*Z ��Rk�8Ǎ�
h6a ��,WLN:6(9��Ǝ7E�(�ntt�fM��#ф��h�i�Weӓ^��_��z�;��@���Tk��u�#���.Ő��mAX���WGMV/f�YA�v��(Ž�W~�`�g�<;Y��2�C̔���+'d���O�3V� 0M\+��t�kD�sm]Pe����� QXb�a�X���'�d�
�������~5�9����&���Xv๪���P	#8̈́x`X���h�ͥ�:O�#��{濽&FL��O��}�y��_�|Iw�ĴYÐךC/c�G����}��h��w��z����7#nӨE�yT�d��J��L�����OVq^v �?}r153��.���	��:�1�g���|�X'�h����gM���'69�%�)��؟����yF��1i�)��V���<�ӕ<�����s�e��G:��izE����[���t�<6.�oH .N"<����p�OLV��MA#<���	����b���oQ�N:��0wr���Z_�S	�-�,�Q�����p��̢&�v,K��&=�����LN#��q����l��.��;a�4�|�=�(' NG¦�^�D�hهq�~�F�;�pv�texm "�h��ǀ��3"y��.8�X��ؿ3T�f�nx�&N�ʿk�E��6 Uc��S�M����􎌜$#ӟX����pk֔M=��|�n
��)n,�%Dg�,8�'�����@��Z��-Ϡ3�oL�����Q��Ԭ)16����������*D�z��-G�
��u\��tT���~��BO�:2	�D���#��s��L�:�=�������Z�$!n�Q�)���F����7*C�&$N�K�D?Ko.>���栝Z+�(�Bg�j��ͨCj6M�: f��!�����"� �8�0��79Ę�Vp�%ey"�}��D��wg2}�*�,��qm��I��?��2��*�6��Y���!�jYǊ�YL�����d1���9"��>\t��� _�������o�{��^��Pd�=�gև��\����Fc1�-�7�d����%��%�m�{JAx�s�18q�[B���z�wh�+�~���Y�{��l|n~��v1%ފ�8�2J��`W��<]��� ������`!S̨R�xG��˥S��⁧��s������u�����/���,�e3��Z�4�׹�6�m�z��3d%z��rAR���������\ds�� D.fT���񰫄P3}��[��8WF�Y"�_�Ɨ�I���F^�!8ڶU�0��m�W�#�X~4���B�/i�.#=ԍ*��=A��s ��)�;]�����H�v���,��$l�J��N ����j��j�e�E=��.�������H����aa����jн�r�e5��Iq`XG�<u�]���@�'��d�$2�f����h�"Ýy(���4#�U��ѿ}@�>�d�� OCw;�?v3�V��L�̈́f��dB��_�g���K�X�=���
���Gmzy���~�.�L`��y�9/ �a�aD�z�j���M�W���A��LՇ
�~��$WRۏ�=�"}��T����ɝL:��.��٘���-����uZ4ӫ�o:R�q����ԽZ�2� }��$XiѺh<0�7D\�cs�/����t���������P3o��
J}3���`i��YR6�BW���Nr���N�؛�q�X�-�i)Β���~Q���:�#n�$�Y����n��9{���$�J�8�H����e��h =��b"�]�߫s�Z�*�s�1ogX�6	~�UZo?�K&v�2��O�� H��Yo��,5��-x����K��}V<�́;t����aQ
�&
m, ���ڹ�G��I�vw��]��s�W��W�gk�Yo8�u@E+腧���eQ'Rᩨ.`��F�����ߝ��N0&�l'_e�+"�{3}�!\�g*>)��0�4����4���u[M	{����-��Dn�sH��{B�Е��#UY�j�3���f5������epJ��
;����N�-LO����sJ��ס���֠ǩ�<ʻQ�,�QC���R��1^�?ͤ>�Y�$��,,�W��]ߛ¢j�z܆oj5�7���Nܮ�L�%��5�5#ʢ���j�]�4�w�ɭ P��I�)Ѐ�����$+L�z����u��|��ֈVV&t�ʓ8���)r�H��DE�rG�Y����6i6���I�ε����W4�:h_�D��&��FM\_:�`�������!Z`"�jћ�]��l�Z��v�ߣ8۵��O���c;�t]���P�R���x:�3��#BO,���!���j��Y���.�H	Q9���ܶB+p�6&�[��d��ی��+!�۫|�]j>q(Y�_Ԯ�<���7{ϳ��R�6��D��ŷ+X]v�6�H��FTIx��5F7f��Nٟ=۩ܓ7����^I��D����]1�iLT9�2Xwg�����ůK@�����re̝��?���\_�s���&�g�5�_&p^�F�-��B;�}���	��� ���y�~zH̻\T�2�$,������xp�
�#h¼aW>�AF!�dL����F�}�D fcụqX�E�SER��\u��"�{�n#H�ǣw��m1ފRE`�E�w�	�ޠ�n��.]Q��� �U�S�# fI줴�;B�������u��Vd�z�F�̳�)+ d��*����?��`8c���2(
��7�SNu������G�,MYm\�Ndm5����&,�m�=�-;U�#s�6�dKyzrrG��E�Eϼѯʍ�a:0��7g�f�O���F3�̾?�t�`H�f�.� �#"���K��-�-2��#�W��c���x�9_"*���J£os�%=I�d�������G2	�G������1�i����߽,���o1��벨TtH�)�ہ9�0�A/CԷw�L�s�ꡟ͠t�Y�<���n�>�?/��o
����2����ˁ���_�7˵Qrck���R���<��`d���^nt���z踫[�9&��s+����	t�`d���p"K��v���	F�
�W��J<��^H��"Ӌ9��f��4���[)�I	7����y��N_�'~B,�u#�8�~zS�v�`��W�D�,����?�?sF�Z]SGD���_u��/�[dc�.��1�#�4kNJ"�QW��D��78?E��'��|���i���S�C���\
	B�s�����x��A;��'��^7(�������@<�`��"�h���0�TwzbkwD>�kd�MD"d���f+��J�������I�䟍�^]4�цC�+���~,����~��JS�W��i�Ii+�kǫI?ss���"��u��� Q��H�,��ʽ�Hz�&a
��jH�xކ��.~'���}�'Nl�O�[<����U��/�7����e�NQK>��=��&^�����q���+#`�s���DaJ����4\(t���E��EdpD9ь��3(ih�q���.�Dm�bev��"t~�ut�]G���Vt6s�Z(�^��iVb�6�8�t�M������.ղ=�U�v	Ua�DU�	��KH��c��Vs��Ry�U��P��a�(���'�ɏ�,��r�/Z	fxl �d��yv�8�_� �N������y���  ȝ�k~���&�.�;"1�q1�R�s�K=3 l�mu{g3m�Ɍvo��-���H+���tA]�����1f�,���0�l���0�4P��MU
qO�:�����}jz�kߚ�EI�M9WQo�Z\��DS��$N��2��v�H�4J! ��H��+�T��v����5F�Y�2��]��~[��$�|�l+�׏c��%��x���~���Vzr���9�Z��V��d8�G\L�r�,yvlaޏE�{a��܊Ǟ_
 �w0��z�4��=�����:����|�s2��k�ʾ{Rb+������|*�K�e�h�l�Qm[���5�}�=O�Lg`{κW�w�S�3O�~)���_���ηp�y��<�Թ��?v�Ց_�e�u/h_��!��Y�1���֦�G?�zIv���/*�A���$��<@��K�$�@+L�S���u�&�u�d�=rn8|h�z��6�7����(�D��?r�KHpqOwCn�����$Kf��t�|^K�D]���I�ˤ��}�ilX�KB���16#���v���e�'������D��� ib���!v�̈�;��Xe����T���\vv�6�E=3��|l���M/��9!$\�	՟~?��$��J���p�4�{2�<�oE��T�,+�!�&+
��IQ㖔�KIk�S�����f���)���5��l�s�04�I�x���{�Uw��ۥp��9�yD^\���l!�sK��}��s��Eԫ��G��s;y*�cd.p��Of5����[�Rn�����HE���M�Zt�HD�Q�H�Hh��5O��]&I]� ��"��4�σ��
R�D���(,��!�Y�<��U@�k�M�F#����Aڣ�5D�'�}��[��U����9[��N���J8�]v���ғUh��z�fL��y��W��K��/��$`���D,;=f~wZ���E�8"ԗ�%yo�RCf��G�:��e/�����UU�%��<A�*}��ʽ�o�ӵ~����j*Vr�kv0�`x��	�8�{��2�BD���w��O��2����Pv��� (��dRm�)M�����b�;�����"�B�b��m�3��LN�4~�M8��/�!��sЄUvMnP(�4��1~WXm��«s#EG7�f����.�,��$o�t���5�����QB1�OJ��d�J��řy���oJ�7��7�)㺕�ZE��l�j��5�W[3����y�����<����j ͔�P���� �R�Q#U��$Y�7��jFc##���hyt�MWx
+��<�'���]N�������Ǣ;\��O		�a1������>�V����2:5;7�@�H�L��������e6���__+[�����GǛ$�fݕ0%��}Ӧ�O�r��A$pCG�da�:���[��rnޙ�ʏ\<��nMs�$���K�K�a �Z��I���)��S�=�z7��k9R���#�T5��OϮ�T��r�?
@(���T^3uBs�E!���l$��� ��څ��R{�2�6h��|-������c���Q��v��[/>#�PT�!�{Q���"D��w�SC�u�O�RD(ɸ_��~��!Y�
9������'Q���]�����͹�7���keg��+S� ��������i~��*���(`V@�V�X���w#Gb���NB�SD�@�?"�E�co�\���͸pr�]u�7x�UQ�0H�h� a[W���H�����G�I�h}C���#��,�U�[��I����JP@���G�!�cc�����y��l%��u�>����mD��DO�N�ԅ��>�h�@;���LyQ_굨2��:�"�o�a�|�b�e���c3���0N��[TŬx�Gj���U^�ֿ=�N���Bc�����K�SzgL�lL]�:s�<G�O/��M���W���UD���+s��N"�?���q������Xj�����yA^��WD�rv5�jow��Sb�lY��ڹt{оl�� �b��mIzWKo[!ǪC��:k��7�`U2��q� *k�����v��(�����c���`�<̲ށ���d]�=�Т�N/@T�`q�#�ȹz��2j�B��5�~��.�n��f|�'�����@�<,UG��E���O�2�l8Z3R�q��[Y��p) ���͡��_*f<�xXO=��$���%r*O�m���t�B�����`R#��@���E�0t��>���Ż��2�ӜŖ��݃���=+*����)�S�*L
7!V@xK$C,P��
+�~�.ts�$��m6&�{)gq�+P�ky��n2g��;�=Z}J��g����\x��r���Z�lT.U#�f�C����)�
yn���j�	����T*Jk���5�Z�6M�Hh8��Coɿ�~��-2]��}��5�Rs)9�2����9;r��"��a4\N\�)�a6Db��N:�1@�X��+�����ٙX�o%��:�/��)�ťl���pېc�LvW��s�Z�^�J	p� 3{te���� �"��O���_�a�x�HW�a��~��g�����r�>j�3"� �}Gɔ��j�Hs*��0=��P�wD��ԯ[�(�������ֆ���l����iPc�̥}Xg7fA�k���$e��\ h�Y
F�����?�J��w�#�O���~�l��IA��>�6����|.���E��C�].Բ}O]�"���8��ʶJ���h�>�\uު�q��n2�6�^��f�Js��G�q��k"Y�qQ���
�bh��9[��(�F0�b��7*W���_&o���]�����$�m��	��x��;�{��B��D��Q�uT��s�U��Z����A��� �o#��0�ZD��\T�I��
�EDB�*�_�L���w?W�i�aI{2m�D�P�.��>�6NU�N?�U$j@M��_<�!���V�R�O�}-ȡ{$Pdj�d|ZipY��y:PO�E'�>|�rt�����A��Y�H3B�!o�`*�Ta����K�~�BC��ŹC��P���&V�^���pX����H��$uGD��hC>y�J��2�U�J���V��[��k�l��w�1�	�q�Rۓ�S2
,*zW����~J鞼�ʝ��Б�d�gɄ���sŊ1t]	�-.���:9�4�ȵ��ƌM��M�%��R�{&k�z�9��	�E@��m�K��P��Α_�%aFi>�e�:dg�
�3:�j�aW`�|ڰ���2��ֳU��G���i�����P�w��H�޿�YzR�Z�/�C���N|��"�_1�dD �&��𫡱F8g7��FǪ�w����}�Z�$6�Nc݅�^��:&c�tI�{��%~i��ج���7�R��*t�2FX�?z�5�u��iV�����\��L%w��K +.�[��擽Zub�o�M ��{p��&��"9��X��UW�&I�>97�)�\M�}��	�j�h�q��ueBL�c���2k�|q�X{��5<�	�� ^��HV�W��ws�(R"ߋ�(7�!���Fh�C�.w� -i���v�O��AI�B�����Z���D2���f��������z��H���%����h)�)����� �E���N#'��M�Ώ����Q��S�E9@�	a�s˯�j��j���<�I*OMl�(Y�����=NFI9p᫺DJ�Ć��v�Gj��G�����k�˦�ŗ���%�䌘S��_Z� M�E�"�6�@���h��-�g	��R���f�&�.�OXƁ��1�2���!vB
9�S��u�<3�2c
���߽����@�~�Q�|�W�n����	��=>j�p�8�y�ȸ�R]���K ���z���	�[�OI���_a�<	�f�|�M��ו-,mk32V"�7�^��"�iZ���{�������n+-B}�ڙ��Lu��a���m[�fZ��S�����7�k��qэgm����+C��ߵ5�p�y?���d|�a���y����ȑD ޮ� �6h��g��!���{�.�o ��}SJFhzHz(P��Ǆ���h(M�y�:u�7z�@ף��
�	�psl #�AvJ�y�����|3�!My�v�$��e�� 9>�p����>/������Yun"��[Db΀�R�ĥ��cFük��n�~;�i�Y=�E���M�췓,}�0x�kR0� k�na�����{��������
6=���y)�g����R?(Yۿ�V�S\�&{��0XE�SN��eX��\��RO��j��h�[~��S�Ḳ���Ԡlh3*=��+A�5��O4���P�Ath�� pZ�n�m�;��X=|w�	���N���%�zX6�!�G�7v'mv�Mf���9x.�8闸��e|Ie4P0�� u��˺ȟ���8%=��d���ۂ4��7!>��ueO����B^W� �Y����P(���=�*���Y[�(TI>�mTJ���6+ڱ�1S��q�>sg)A(A?�G���C��׸W}eN�l���ah�kn��z��8��~;d��}�84�P�9�h4]Gf�[h9�XY��R��\��*��"����9�Pc,$�"��LP}���y��y��Spx�f�NY�*�Q���S�r��Fo�GL[I�`�y�zW�X|Sum�^V{�Z�q
]��Yg�x?%6s��Ҙ��.��C��\��O��BE9sT)��O�.�C4���p��K{�m�%��ʺ�@�&͋q�9�H��Z!�����N6:���쩍��<�G���y\�g�qmK�m��j���n7{Q���i$Ш�m��y$���q���i�OU9L�±�ao����|_��F�^?�v��ɂJ�����A�h�b����-b��g1���f���iT#�2��}�fԬ�Ã��� ���&�#�`=@R�>6��d��	@����-�.X�xcqo�ՌD��
Xu�.l����ڦ�.��O>zr�T��ó� ܰx���p�QV��dqf�6�>]�#�쐹s<$+K=qdQ\�jz�J�nv)�2V��'���Oo�q�L��� wk���$��h`P�~�@3�dw�;YnG׆��G��	��8[o3�ڛV��U�z>���'��uV�YV";�<��Qad��D�I��/���[�6����n�:����[I�5g�#-��+AߵE��9�!۔��$7#�!��/����,�^bi���t�W:ȝ������sޝ"��w�ӨXKz�|�!�ᠥ�.�A�g�'�O�K $�/=֕T+W�"`��UuuR�{��L*�]�t�KK���US�$��?,3�s�:rqqm�)�SE�X��y��(4G�v�S���YH�T��(w��Z��DW&�I�
S'{m�օ��\0�ܸ�EIL\�_)R��뒝\Em�y�X�j�Fnht�x!��ɂ>+�C�f��-Xh�d�P��㳯Z�	5�	��Yb�B?a�z�w�&0������I���)^8Q��� l�g���)�g�f�w�+���ۓD`VYUu_@n�wX?�z�`-=w{
Yy3�fbm�c���vӆ4�������Ez�vv��]�c��.�@[n[���>r箙0��dsA�����0S#N7�42F_㩕'��N�,v��o���2�a3u���Z������Si��q�9��+nM�C$4�JLI$=!��׌m�B)��BIn�z"_�nl$��	S���Dc���n.Z
�'s^<���BɆv�+zy���*Ԍ pw˧�@_.ɨˌw�3�>���a���!�J���NOgp�rUZAn~%�����:�y���u�^
7'K8,ਛ��1�l�N�W
��r ��l��&cb�}4�0��_�ĵ��������E ��;��~���`3���Ř��D_W� �QJ���t��/�޷$}4���u��~�R��� 㫞�{`&��F�#���`>���_�a:,�B�e�XyW:K�WppЄ��9��	���s�9�,X|�L@C��XD��� �Yb��08��u;���v@�F�,]^= ���p�k��#kl��d[� ��=�� ��)G6��@�I��$Y��w�T���Z�P	��]/+$)�A�q(�/}�x�^9�X�'\.!�J���Z����vt�,s����Sb�oV�轶��G{Px�l�0 D~���P�=;[��?_�T���F��Jh��Y#�;eIT��$S�����c�����b��`'�řւĢ��:j�X��X��oK��o���*�iީ�Q#�T�0��ǈ�tF�V���V�@���,9� sr���o��tn�,+����#� �0��(�=�3��Į��k�lȷ�M�qwҢ��=���ҼSO?<��ݹ\��|AorI2�T0�ݮ�w�l����(-'��&���e�E�#��J�,��A���2�ճ�(�1�����ʧ��Y��uL�]�%��h2�r�LC{�>A&9 o�{e���D��JPO��P�-����78Pa�|�A�� ?d����ѽq���;��*�Jշ42�t�
;��h}0��H��Y�kl���L3��֧v��0=.�2|���yz7��Z����~:ا/�&�D"������.���V����
Ir94��R?�\�S���4�r�G�	��$7|
6������T+L�]nU�#�JA����W��d�b�n��D�DEE}��6.YZ��T�ǌӲ�K�oɩ������4P>��L��EQa#/d1�� )d3L�NK�*�����^ױN��dE�Zl�v=a�Y�~���/R��F��Dr]g���>7٪��9<���ƂXXx,:9F|���@gO�J"����ۢw��쨰�c�D�DZ%9�`�G���|<0���8���j8�`�؏'��5s�L�iC�t8*��]Iq�_T�JWá�:=W�����~Q�s�7�<��B�,�bE��p3nh���D�:A3m�ke�nw2�J;�	.\�	���^H�gdUჄ��ڠ�{��[�L������3
2���Dt��]"��O���jCb�Y���P}}iR>��ɘ�x*&�<(��w��:+��)���RjC#��恝���Y��9����<�M_��b������u~��0
p�� �X<�-��ٚA4P�6��,��K�~��!���$����j�LF�6.�b����9�V�I�k�?.(�v�l�9p�B5>V�M��>8DO�ϻ$$��q�5/�)��DfY�X�$&�/�����؜A����sZb61�Ff�����,m��DhíM�݌����zQnP���Jmt��v�jq�`�d��퐙
�4۩�k���]��A�h%U.�*S�3�̅��FF���⿦�x�n�4�Ǥ�/���09I=$�-���ot4Nh�Z!�%�	�䄧s�V�9pb�s�(OT/�^
�ѪzH�hY�{)#Ҝ&f��r�E�E�>Ň�fqM0�a�/��۶j4\�]��yb�| �wX�?W��r$.���z_�/ե��>��VT���-\��+��)� �szx���C�Om6�<F����,d�8>�$u�]�)�R0�d�ǯ�70�5Þ
�_N���ٗY���p�Our��,8˒V)A
螯p'�g��ܺ�]31j�ń�&��;�Rl8�:8��a:��)�_;#����N�9��f��A)�
a��y�޻���i�'�2���['@xE�[�� b/���j�M��!K�Fc�g�M##��17�W���c��fD�xc�
�ѧ&7ƽt�ϛЬn��fċ�{���"��Hg@�,&�{�z7$S$��Te�j�C~^�Eu�Od����02������G��e��uZ�-m2�}����3`"�@f���d�e�nf��Έ�#�$^/R�^�O3˟���' �tέu�	��.g	�4�)�5c|U���~����mh2u�8��\P��W��h��_�D��rJ��C�ʕ����q���i�*��nְ�
1�}E�|��B�Þ�
!S����cC��L+p�Pqq�g4@V�����T/p���9Iϴ������\�u`d��W�6$�n.��4�V|s��+2��o�\e|�7�G�ų��;x�J\�$� o(���#�G�!P��B�N��C- �|<[�J�Z���<�ҡn%���Ҽ���-�:�=[)�~�Ѧ�c���S��}��~�H2�Xs�����ʠ�"��0]�OrG&ٚ#�[��\��Gݪ)�����[y��$�����>Es7�9�:Ñ:�$��r�N�f*ff7<b�΃L!
���A�N�����G$h��a�,A3��6Xf�,����fC]�n){7�[�Ҏ ��	0��L��d��Cj$��R���KXMl�
���
�"%m���y�u�Z����p�Ȓ�43}O�T$�x��+E�c/��\�>��H�i+�P�$��S=i[���臠vWr�Z��T��� ����y��rNC����{���γ�\����%�k�������pfO��̒wSq����0�K�}y� a��g�C������Tr�%�0/�bd�ztT/X�Q�X#�|�>%^�G��J)�ME�p���x��=*k��U��ö��S��}0��p�%���8͂����=-;�ݾrt%��E��QP���ٞch�Y���K��<(oT��,�����J2�A��`?�ņ�h�ܑթde���Y��LW��q@6��	�/l.?���!L�p"ە�у��
�/�g�|)~�+L?�W�G��eQ���p4Ix�L��ݘ[ݪ��ң�Q+˧�
�`ԃ>�4N���ZK���������i�۬o��r������ϯ�qr������r�[k  g���Y�sf���W�>U����Mc��^f�ͻZ#{+�1>��T����7m��;��Zֲɍ���#��Jʲ��Y��8f��S���9	h;4�e��C�Vl�*N$� �� ��s�w�_N�	��'ԷI��FTk*�g�sP�1r�q�x��^M�:"д��l�<��I� _%����V�cFS	Uo�����&܊�avlv�W��?I�f7>,�A���_�p��NQ��C��xa$d�C�XJ���A��&�įB%``a���=jH�y�n
<J��a��A=��y��H0Ľ��j{%d�3�e����Q���h�4u� xH������5��H8rF��&�-TԺ�Ϸ��k�cM��y����"g�X�xN��L0P�(�ɣD��������w��`��-�����kOM�c^�O�jQԇs���;Ӗ6�9�@y�(��99m4v�[��F~|���i��,�T��9�Y�;ҴX��.���6m*�%��:u2�KN�h�泯r�$�8��˗��<Z��(��>.xӔ����k׻�!�D���˓@�%v��F��f�"2Ǘ��sc�A��`�����b��F	�zS[�l�*#���W9C�YA|1񅖝�/+�+�e���N{�p6����3�1�W�f]���곥t�Ҍ��J'F��@�8tT��_��Tw�g�8~j��v6��U��lo�1|��k��Τ_������˘f��LY���κZ��A�976��Y��G��:%��q���.��'w���� =��kQ}�jjB�3����'�P?5����H�����0�'<=£����Fa���gΐ�fi������ޱ��H���%�`�d|��	������R�����t\����xU ^�����Ј����ʼ8��M�MY�azwFi-b'?��$sk[L�3h��a�2�WgP}�e+2�8���_��jMBTQ�'m٣<��ԢOp��k]�=#�&�.�.��|�#�X�Suـ46F݌	
4٧� 5�G�y��i@�tn��y�)�GO*�}UaƘ`��&�EЇ���t��&f�t5�<���zi���\��N1_a{~	\����(�p�*;9F�����1���f"ǡ'������<���?#��p�����}n�:��г���OSZ�"	�;>e��D�~�#��D���ر� �ʛXᤏ�On�9��\M�}L�C��J,���?�񽃘�J�͍�����>�������w�?՞�po�q��p��4��cߤ5�p����']�K����Q:�6�޹���A޾1Y���V�P]�iB�21J6i��}*��~K�B��z�z<>t����`o�krzfT�w��MN|��P�<�&��[
��- ��M�p�ׯ3��}�A���ꇷ�**"[�K�h>"�O�Pk|�K�_�,�Z����'�N�퓡y�����i��BW��9Ґ�#���I�;:�9Ex��5~�æ���3z�$d?��(��`mia!mSδ��q�L��CC��Y��l����U���έ��+��x��N�=��~@�K�X9Kh����e�����q>�2%��9�/����������L�������O�W���7{{�p�S���Du��w^��SSW�mey~��az�tx������9",:(7j4����>���R�ZXA�N�vlx�����V��Ĉz&�5q?#X�����nS���ô����48���[�� ү���'jS�=C��A��N�<h�љ^z�Ŝ�z'Z�-G�H�8U��p�	ܢJ�
���%��i@���4�2�|>���qx���b#7�Յн�ԑ�o=F��i�}��&O@������py�HP�0���@�UX�#�'fЕ����L��.���ϲ��܊�\K��kn��	.�
��!�N����.����<�)^|�0<�Ⱥ�ױ���ln	-����V��"�H�FYq+�}��a�0%Y�jJ��U��C�A�tA�t5��}7��b[Q���	��@�N�����l�Ģ��wթ4j���x�pU}C�꣸��ŋ6���_z��$כ;�Q��/&E
�d���? c+���ȫ·��6�ƮkC�K�_9~����!���@]�i����]����V3=D�����h��#��/J�q�k��`��f>��	�e��̮lBO����y�ogԆd��0/���u+�u�@�j$&B'�>"����a��r�2���E��kyB�eJdi�xvO��u}�Y�'��+�/}ׅ���:%w1
it�rD��B�Ž�U�!�������i��ޤ,����UZ#�DuS�ߜ�S�	D2O	��'����F�����~z(�=Q�����w�=v7�%=�X
�Ju�E�a+@�'2;lT��������������9�C���3R�K[X��.}1����0����wǷ� Ʋ���^ &��͚��K�d�!ґi�1��IgX�J͂)�ڹ��RG`�s��P���D
}5T��=�dN��菧qmN�^w�u3/:5O�3�;�B�rc�Ok�/�Ku�ʵ������K���NFpF��-;��!/��tղv�6}��{}D}\#��_uL0���Vlu)��RN��\��
Ui��j
�<���*���Z8��i�J{�*{B֓dt5j:zf�2�A,�g��(خ��K����t�*"�)�[���u���z�O$�۶_#�vPj⎩� I��y���/��O]=��{�o.���k��W%IF�idy���Z�G��F*'U�S���'DY��HzX=��z��7��5�+�UI��d���������n81VS����]u��I�ؔ'1�\a�B-��1���⁡$�������5wM���վ�&Ӗ�b�F�B�����0������?k��F~[���̀�����x�����yX��.�B1)?_�q���z��B�������X�D/�~����>X���4��8ͽh���y�����&g}��6k����+f��*�2_�XL��8�
zHG�chȢ~���%��ݙ1f���i�	F���7�JO�ǎ���|�M��mhm��N��᫜�3�z�)օo:=�(���)B�P�R?�w�њy��!���f�r3~���6��T��`v-F�� �T/�t2�e����Ú��ܚ	]Rl�r��"�q�#���
������Iim�3��w.>���#@2&&��{	�#�\�7�k�sc�Y���6�,a�	����B���j������o�'N�<݅�[����s/F����g+! C���8<N�.tE�g�}�*������bܾ��_wf?�4�P���� d�I(rsҊ:O{��,Vf�m�1�5�r3o`f>��ip���sna�"|��._��)H�%XA���zJ[�̕��#��Ҹ��9!�UV�9��噦�i�"Oz��OHˊ�Z���NS�;Oj��e�F�,N���
Nb[�F��֫�L��F>�x����Xd�J]�8�\ިk��j�*Vz�����R<{WL{�ZF9��u�ɢ
��"��B]�]��8Ǔ6�r�����3��5�B�qoN�	�}DN�ĘZ�u>�=�&�S��.�T�3�s�Ty���/zmI�˸�hi@� ��0�AR�ql��?-w��o\�o��Ac��wm�!bθ4(3���M	��4�3ť�5�m-T�^� ����̉C	҂�|p��$J���q�Β�
?�a\��6�g2��(6$sH'�| �9t�'f+a�MH����S�e��@��gk�C ����K�����e��jewh2��~�c �.�>�l��|p�nZ�����֟Sf�|u܀��Cb�ߍ��I�nQ1���C�n���*�[��f%�l	i׎.9V*���%K�����I�J��*G�6J��5.*2^?�-ֳ(ڒH�B�/h�.��#Q �8��q��ԦoaO�c�~=nA�0ؙѳ��.5p�,��7�D���OD����9b���ՠ�-���@ԙw'-�ܯ�Ϟ�����S�46�Z#�"9��à�8���V��2�3�Lj�m��`�m{J>�v���d�O;T#�y���5�"ZԿ��]�%O���f���}�qC�v3<��p����F븖�\�l �-)�ᆿ��
�ܭ���̕"��.i?�GRD���&�E����g�r�>�����m}��
����ȏЕ��Y���LiX��8�m'�� ʙ��,K k?�|S����V�o�t*�W�R͒�8Dn�����M!�!wUv�8%��2?@Yڻ����o���jD"��a�-T=nk��?��@CǇ����"$;(�!��\��^D�KK����5Ζ���N��*�m���Ғa��[�O����J��9�ۋQmϲ��H��Wr>E�W���$�o�G#�/�6LŔd�7���D�m�炻��~�Ӭv� -����^�Ϧ�W�\�G���o�WV:'A ~����6<m��� Zc?�gc�JԖu"p���|���$p�un��̬f���)-�h7���e��/��83C�Ep[�H���0Z&IVlo��� ����2;@��`)]�;\k��e$x4R�.��s����Q��@�G�'���a.�����X��ЋH�a�틩1@�!�Zk� ����{d.\�aAV�`3aT(3v���~&�0���3'��uM�5[���B{(^�r%�5E�Z�����h����]�0U�A�2��Q���#|���h�~\�1Ex>m�m���?�����hG�����y�8|���X4��tl��3P�Ɵ�����a��m.F��I�����Fi�t�� ��A-ۮ�2b
ђ���7�}rD�Z�-���
<ͺD�X�Co�8Ĉ�.-Z�'�����' ��"��)�iY$ҧ��x�B��#�N{�%)NƓ������SND|k�n%er)Wr����or!���T@�K݃����ʞy�d�'N�/V�@g��;����$Ԧ �#CKrab��%�����`[r+���>ܮB�����.T8�{$dl�.iC��ǩ=��}����Mb>�Y�dG.���(��v�+�ı��G�[+��kf�)�y֕Vt��]�滽q�x8���`-/��;��$3�K���"Ù��4�$Z���Xs*���?���I�7@�qV�&�����H�$��R�����lQ�KrB&[��Jg��IW
9���nKs�ˁ`I�~��8�S���l4�������b��䍕�c�U}�ԋ	���E4�%zi���}�����@>Ck̔���rm���k>b��,~Oi��M�o���cy1�gG��g�E�(>-G���˓�P� �nP��X��G+��s�A,�p��4�D��UU-"�jt*� *V��љ�N�^0��c��%���/L��C�M����oB��J�@E�� �m�T0�&ԥ�ip,y��I��u7�~?�=MJ/�jý��-�pߤ�=��HL/�{������7��(1mN������a�;7�Tt��a�joƸ݁�!�dA�\��o�z��?zG�p��� �i6����K�B\?'SIK���P��wf�+f��yLS� ZP���kT��T� F)-�=���_ɾ���w�>1,M�m���z��������B�B~&�:#�cM+G��?�������@��1-�t���aYć�=�������ό�����R�ʤ��e^C���6�"���aEDF:��%�}�p��X��ȜAly�I��3`9����n=�2vjr�m��Ƴ֬y�b[���)M�ؗe"��Փ�#^��^�����%��K��6�Tp�Z�Fʄ�4u��i��Kc�������FB��-�S��ݤ���	Hta�'Y7L��U�r�^��S�b�G`����sEѕ'�TK0^��9�$ƌ�����?5fB7�co8у '>�}c�"��QTnv�w�����](UZ�7��&���1ZR����A�{Q��5���vג9��q�Ux2)aZӂ/ ��{,z�@ۨ
����X��$�;J��"
=
2���1���P����\���X��2�nV��\��X�jxFfl��O0�]��hH(�T�<2}j�nQ�u��Y�F�v��
��� �r�n�h�U;�v�go�q�|��z�p4y����@�p�8#,D�������p�ꮙK���=�>���RNu����>�
tW�^�N����I=wz���BU5ODܰ�IOV�a	���UgD�;67S�#�5k*eK��(%�� GǶb��mFL�A��G�#Z���V*kr%Mh��$� �>T4��D���w.��O��x����:7=��=i�k�i�f-c>+;n?�v8��V�=�=��B��Y0�<�GCSF���A��5��"ܶo�W�@۲'���칖h������*[6�1�AGm�Y$ݳBb� ��h���Ќ�~�uk�"W���Hʒ0���z��Ns���,_�3wG���Kc��BS ���p3MU�*-�pɜ�-1�ې�E3�Șz�W��]�K��/@���T�
E��{��2�dL;ӕ�^�ܠ^���gA�Q�¯���f`��	o���V��}+�ɡ>�U~��M�&:��.fփ�F�l�Q������}F�o<A�RRW��5&q�.�����CE�N�I��y���tb�Q{������<��C$�&���p,q�������<���q����}8�=��Q0� �D�\ɶ	!�1�$}�OSQ?��J���85=���C��T�=��b�|����XE9�QH�C����=m_*Q�u��{)�*s�C��%��^[��{`I8?c����9�,��:78䕆R�;�Y��"=�{W��� t��{⟚\Y���q��ƨ�G�~�I��"'G�p�{|Ւ��i��{��F��7g�� �uV���JBa���4��čy]uvx��I8vd6�gч:���2}�L��e6HdJ@��Q�!ARD�1�d���`����D�
�3�#��m���<1="�e]�r^�뜻zD�
VK���=m�;�2�A[�έ(3���陖\�Z�3�-���b��>rM��9}�rz3�]��`ߜ��;7]�N����Q�>����<�-�4f˪ZO�F4nr2N�ˮ�~f�����Zi8�-�P�[�P�V^���ʯm�7��&��� ۜ�+ �w9\\_<k�.��^���x{-c���v�پn�������PZBM�f"
�?$�@���6���0H?zD���˖*EF��Mb?qJ��(ȥ��ޓr��9�a������b��n��X�1��0kI��9�%��_W*�7.�&ݾ�W�,�\����qa
���CCr�y�}�>�UL��Q�g ��.���<1pY���M'����8�F �K��\%J:E�h���]߸��s��!�Y�B��_W�-����5'�M $��i�>�Q��!���Q+������$��쓸��XQ���wU����ҁN��I���+�������U��N�?���r�� ��SP>Fg3<%����_���}�(�ggH3J#.B�Y�HJ��P�PP91�?I�t<�To<�T�l��k:W݀���Y��) �+��z�옔�/>�n���"�dә�Sw$��A=�=�@[rL˰Q�D.�?�ę^9�=�e�+��M�Q��� �8��/�6 i1H(���Pv�S'��\��{�0�sY�Tt���)f$i�>/�]�7d���и�����a1���]Y�i��-���s_ƬS$��)]�B?���fs�B�o��1��|t �P��K�Cjg<�ŧG��s�K�d��ڒ� gW��b�켏!
Ť[㜤q�]�����8� ��n��Lr��} yԊ�q�Ǒ�qM����+����k?�95l�/n"p�~�]�ji���!���'=�<>��Л��ho6ω�2�j���W+J�����ٿ������%|!� J���	o����j���fh�%U��[ N&8��k�^�
Df�y��M�e�=G/T@::F�Xw9OCg=O���R�������υ�j:m��kt�Tm�_�A: �8:��Z��H�Q�ŵ�5:���GK�]_j�'���t���a�j��=첀�cW�pQSm�9x	a�jN��胠3@�1��'�f-�D���ke�]�n�ٿB���פ��한;���/�+B7�z埈ߚ�9�;�
ؿW>1u3-2����C�� �S���C�b.y��B���F�S~sC��0\�q,�b�ٚ�:s�}�q����V,	�4Ai� 1���ꜜ���,t&P����U uWaI�EK҂��2C�9帄\q�t��ʌ�C��\g.��D'Nń�m|G�Hʞ�8G�߯�W��̖�h����Et�����3�1���C����tl�,x�̜�V��0��~�^�d�>0��ұbD�{���>�19h�����~�K�K������a��]����`u���ž�yi�uJ�ߑ��7u�|�FE? ���7�mj�3�ᑝXҒ$;�L�w騬a�&�Kf�Xf˝�r�kK��5����^����b�����<�!�+�^��&�c6�+��%C�Q[����>Jσãҙz7��o�~��N/8@P(��ZŬ#��'���B��E��<Xr�H�<��U1gc�<H,8w`ҁeoH(�%
9ϑA��E?��d���9Xv�Gq-��nHv�q�n�C�.��M���O��>��m@��l/Ű^���M�\LMA�)��Jf���&a�;��y���X�3\!�Su����Q�8	j.m+ZQ=��.++�}����D�E����'�߾���F[����_$�����U ���?a7�e�Ҵs�(���s2'h�uw�D^�:�)A��U{6��e�.�	�<��=3b�k'�G��M����$z0b����ʬo$�[�6���/:3T�E6<�o��VoA�7�[V�
�2 _�_��ZP߬@ l��$�aP%���Np
{9��VV.�TD��M���<�]�6��v�fqg�����W�-7�C���w(��k4C����&)����k�p�X�i�Gh�,c�x�q�����Fʔн ����\5�zr�AԔX�.��s8!�g!3Lg��Qf��I��@
#]�L����a�&/r/ᨙ���y�-NgZrbo&%���^q#�LW�ol+M�X�э��G�N�A��?FN��^g\�f���A��
������7ڣ�x�7?*O����*4ڽR6�-"t ��N;<a�W���nsq$f:��?~��>�<R��2̤��O���9�C����A�z�!KBIY�D@>ϟ��tb��-o�*���F(*��~�:O�,	�OQ�M�acge/�^��BMH���+ؿ�C��TH� ���7j�=Mlj4���k��gw4v��Ꮂ�@j%�>��Q���980Yv��zV�
��`���\;���<�z�_K\^;�"^ߗc�� �B��6�N�N��� EŢg�g�tݔ�X���G�]�U����Ox���q��u�G�+�k�?@�fz��s�ݐy)� c��O��H7�dP���Bq��:?�<��J=#�E��P�,4���ٽ�]ߏ��_J��A���?����9-�o��<��tBY̵f�;�#s�k��2x%�C����	z$j_�E�S�K�*1;J	�wї�K>
R��Vp��H�������1�B�B$��{g�ԇ���&����iQvSF>>��j��������ڐ�'�k������`=�fU����υ}A{;�6��������|��w��
O@�"���?�UE�I�����Q��PP/ܬ+��,�qN�yTL�|���jI�j���Pݻ�����-�k��-:��s�W���w�<�qqL��O�B�<tm1���$D�,.v]o�M�����s\Y�I�J�&�*�y��k����P?"o�i���F'Sޘ�Vt&;�����>�i�4o�*g�j��	�84�3��#����Pb�c�7�3�����iL���G�ZiZiӌ���a/7��w\�eaQ��~O��Jv����e\U�G���Hh�S�z�����T����G�S��B�-�'����^rۺ�<�2pZ���s��~�h��Y]7g/+:�8,��a�z��b�v�^?mA|c�d���1����c�����1?�,uAS"�n��fO��h�^�AO�cMTX��9pNY��� ���MI�'<�n�[��~ZC��J�u���t9H�Z��=��9�1Q��H	��C;cQ������=�0��hU��G��|Zկ�bK�.m�SM>ᆲ�1^�¶d7��~�[�Ɩc�ɗH�IZr����{tWBR�/����#�_J�N�<K;��Tt����.d?��﫺W���ύ6:���?L28\}��Ջ~�~�m�0���{
�{S����œ�l|�R��Yӯ���[v�j�U��"ch�L�}
͉��������u`����2m'F��s����6.Ϟ�[Yh�Ş�}QZ�{��5���4=W��8���8����
4���Y�3GC��9��r&�{�7��<{@��8�q*��F�H�!*J�D��Z� �;6U6ɭ����X�0�v���������W|6���I۽��r�'x;��!8;�����Zي�bg�[�J*����䀧���;��l|�Gэ����Or�A UE�,)A��p� �Ѽ#�0�Q�)�n.���h?�#W�Zw���S#�
D!I
�t�9�k��+�L��@y��ީ6xR�d���Zz�+�b��Hf�p�Y�N+�H6���#I{X��3!i�uȎy���VO������B�}�����"��Q *.7V&�>��Q®$/��$���}�V]x��V���LB��;�����Q	n!J��anܙFNAű1�9�?��I���4��J�a���3�����z|Z�ǮWK6L����=��oò�ă���b)���Yn�����nXF�9q�Kyf��8�Ǒ��k�B��_b(%�РXWA��w��d�6�J:4$�,i��僳�=m��W_j����*��N3Sp�U{Ň�_��E	<��^�J��C�`��{3y�t�ۓ�[��D bŪ�3��;S����ޣ*o���B"��`�.ß��`��r?r�)��R��Aۛ�}:�J`��&�@�t��ib�<���z�3Fy'	��"������m`3��.Q�^r��t��Z3�sݢ���s�&L�ϧ�UF,^�����n:��T���@Њ�b�[맠�ဪ]���\2��.���7�
�Ըm�n�]3�y�[���u#U*�ٷ歛�kSz��=8��0��0x��M�|KB�-$�ϸx�WO�p�hzO��x��O��$3|�,>�h������,�����ذ�b�L�c4�i�K������D[�m{�Nf��SOru[_#npQ��/	�|ٙ*k7����-~1�;����g��k��1�Wt����n�2A��;}���wWJ��61�">�:�M7e��Z|,�@~��ң��S��^�:(0�C�	�}yBC��k]��-;s! ook{@ �?�yc��:H��V�r�K�w<�$�G9'0֛.��zٞ��P�<jQX�;g0Gz��BFi7�m=G标�/��,?��!�ؐ��v��Ӡ�6G����V!h_4Z.��rO��>"2{`u�$�l�W�kЕ���<�"�(�wM$=�����ݭƊ�@��+������%��4�=U��c`���T?NO�~YxP�s�9w���SO���k$5>u{����;�i��&��b�����J!�Fe��EBӪ�����,}g��ac�=��^�5��J0���)(Gf4`O=���.o'��[�<)���Z�`f� kØ�G�*v����<�2�m�P�/���I������ЁeQ��In�[�p�]��<��e<#"��������*Út�����8u)><��'3J"^_�9t����Kw⁒~���&C�{�2�R�ѵ�.�!2�P��	h�f�B����nYָٽ=~nH��C�̃���A��+�x���	��)I���t�q:7H��f�S/NB�Q����B�ջ��nд8(^s03�e���I�w��!��Ha�V����W��=û@9���_&2�0�־�S͡ɑ	�!p��7��F�C����� ���Ҳ��J�
-��?x�u%���C�|a������/�J�Eczo�q����3�����{inK����Y\���߀�ľd6�g]5W�cM<5�R���N܉|6*�J�,RN�-���Ԩ�0������yF*��ly����m��Ǹ�J}ڧw�M;G�r�E44	ry��*�u��#��Nzc�W�*�*A�A��lf�d"�Lr�I�`�h����"���V�������~rev~xԸ�,Dmd�;����=��?ٰo$�2d0��H�e#�b�n��ɍ7l�M�Na��j��Z>��_�+v�c��P�Ql9Y)�B$��%��FT<���_)�����R��V�l��&���<�߮���6QK�%݇N��I���gQh��� ;-G���pIE�딪�i�k
��~���,p���-I��ށ��zh�c�����m>��]FnZx�Kܗ�!~m��K����H"{SM�[����*�W;m����I��i���*L��U8���/c��0[������L�% ��vٰ�]��]���m�GG�q��l^��;(%��1F��-;�3IQ������	q���5+��:u�����ϫ��T�� ���g ���\���=������x�4�2}�z�u;�|�՟�1�NL�.�E�O]8�!��8�H���K[�[ B�z�h	Q��Y�yE�L�H�/��B"7מx{1�O�r����?����L_�I?��G�Cr3��}	����Q>v$w�%�Q[ILU����E�*��p��sM�e?�{K|И.%B�	U�v���&c1�Q�߈�$b��ت�������M�?�o�cqo��u�c�g`�W�Ȱ�G�f�h���F�Z �E9&{�4n�g�Z�w��\8}�~�d�sMn�!��v��P��o"W����3���%�����Bv}�c��*��a6�a׌O���
\n.��hP:bz�	��K<g��ƹy7K�#�.R����"Ӯym\�y^Q�*��;l���v��5a��>�[Ԉ�x��Io�+WU�T��h���#o��,~��M-[���Ѝ���E�2�$�z���hY�z�Z�U����o���_�)GJ�����N�'�-l�j����ݬJ��Y�*� */mmぇ�SpHHT����Ȭ�4>��=��:;��՗��YĨ�.i0������EH�ٹ圠	�_��Ym�ro1���Bh�*��h�
_�]���A
A� ��c&~���e�(�;-����}pTt�<؄���i������^��a#ݿ�i_�x���b�q?��[�^��kW��il��M����YAt*r�燓q7<|�i%Ahrqסl'nvT�ɣPd2R�<.��M"RP��{®s�䈬��"���/Ջ�X����1�%�pC�t�Jdf�h�a!L�Z�'����9؜�Y�Y+��ܺ�o�����7ql�5��f�eiS��9����z{�7=��韴x�s�(��=Mg�B�������N YU���R�u�;'� ��f�WY�'r͞V/B�N�񕗸L��m���=4|��Y^�N2"��Ɋ�����ߍ��ob®ӟ��:k���Z�g�-#ʅp	�ד���o"���Q��:?.b}-�suҗ�BѢ'����-C7.R�]�� ˀ��pV���u������=�X����8�\��@����[���A�&�^�\4���!��  `BMMZ�K����oN?��G09����zn�OA߭�i��l��r;�ؑ���F��*������Y�YK����M�TU���ў�T��;q��`a;s���h�iȂ���%uL��W�&&�v�VC�[�a`G2���xQ�[��'P~n��Q	t�(�<��M���X:�09t�0m���iu�Z��6A�8��b��]b�����7i��Ӫ���+'��A�ua�H���ya���K��&���-?�	pf�I�ٺ�A���T��0�N�2k����-�:�F��v�/Vh���X�����s�<����ӓ?�`��@��ƈ��Uh��}$��AME��X4���,���/ϒĀ�	@U|��lf�1��*s(�o
�ʨϺ��f�N�����nv��̂����+k8�z��o��9���Ȟ���EE�^:�l�ϩ%9��Su��->w�%;s��j��[��Z��i_�-}��&��Qh�ܔ<���x��RjȖ��(5E��~���$i�;TP�z.U Qal�ܖ]���&p��]��zOL$^������ o\3`�^CXu_e)��Zei����̴?#qY�����&u�3A峐w�h[�~U{�F�O� ��0%ɡ㛚�Č�U�����&�Q������/�z''$��	�H�U��5�>K>Зo�W���`9�S�s�D�-�r�I[��Wۺ|�I��4���L��Z��,����\J�/G��U�wx$T`Ԉ�B&���d�-I�F��B*E�i�3{��">��Ph�\�ze� g0��%�w��L�'� �^��<�e�rk�??*x���@�M��ϔ<��+���
�ɲrT��5�P��@��l���"�f�P��T5#��@�S {w4�����i���|V��n
yy���N�$�\P]tFK-��d.oLʂ������K���'�f�W����;��\���w�&9R��eێ+�f����kp�w����F��$3ᩨ^�ۥesH�aW!R���� 6uߠ�����e�v��\>ZJ�������H��#ŵ3�~&�T���6E� AFA��z<�Y@~(���8$(��7�Uu7� ���׾Cy��@�ر�r& \?w7���F���k��x�O*���NRl|���W�żǓ�0Ə�C����t�\��]NA�q�#�B�zLEĎϑ
�%�5q��E��-D�T���4�; #N5̎8p=)2�/��a��H�1���6󗌿X������-����:�;�b��W��a�˾"��SO۽��c&׻~����$5ۚM}���π?��߳�����^H�#��RqW��У-���(��y��%̫���CE�9�>+e�_ ���=� �]m�g� ��Bה��pa:�=�T����Hx���@H��`帀7��ۅ3��,�h�o}�,��uܪ�����1ý�0�-B�]��<�QC�7#��v�'o�բ�n�)�����o+ֶP��]�<���B�K��9�{�W����o���x�%+��[8�\$��=@�����g%��1�%�k���aЬ��=����U�{-2����m��$�.`��q3��A��-Q�"�n-�p��|�,!��,�&}f{׈�*kP:Ϡ�� ��@"�=U����EK�M�'�饛=��ܜ�E%(=�����&h�M-�j���E[.H,�w�7���������@|��8��Q>x|����Q;�;��j<�7�OB'��ӆu�B�UG��;aǘ�'�P0*�D��\�*`�KI*��}�Ģ�ӺjS(���,$�,�ɥ޲��MR�J{��b����Γv���^G]2�0�u���Bw�Z�M���a�d��b�fז�\��5n�_1���MA�z��+� zsn�5��wx�{4]��*ȑ�խ��U�ҿd?����D������.1z4��yԭ�5� 9SSB��O9�5Q$�������)٬i0OH���TR��$_�ޥ�<��~�e��)�l���o�g:��YQ�$G�`oH��i����K]��*Yo����mh��A���u�����[|睴��<a(=�u��P�̰�ᄡV7��,��n�9_?�dd��:8\��� �"àZZT�-�"��������������͕�o�d�ez����嘎����tи�E)�e��J����}`����R��s�MOє�ֈv��4O�eA]�Ʈ{K�o̰��<!E"��f��	u����W�L^{��@܅Lέ`��&t{��~����1���=��TR���i~J�^F�O7Gn��2�����ZLǗ��X�|a��<���L$��k�V�%O�VntEyB<k�B��������ay%���M�P� :FЗ�fJM|���<�C�?6�;���]�9:�j ?����9���3�\ɰ��ŷ�vs�h� Q������*@ox�g���;�q.!���{�=
��ǩ��\�o�����Xcʑ&քx��AHG���	��5yT���~���r;����!FE�K��{���������KV�:ÛN_���(�2�؜��*RU:�U���˸%���b��q�r<cN["�=��������� ���Ōp���_����=�+�)Ⱥ�Z��K�����ky��$W�ڶyɝ�_�8c�+S�0��J��1t��'D�C�u����J��jde��}��$�f]�:8��&��r;����-�)����2 �wK�C]*�Z�o ��2����,t	}X,񼛻	r�\�c!H��v#��\�n���C��Z��"�!_�5��ۨ�� NDc&Y���z��}0�)�%�q���f�5�j}�\$z�j�?g����9L����F*��`�ns:z�m2���Tw�ϐ��L�2����#�!�*�ӄ'!�"Q��S2��������Wn!P����k�yd#'b�]E�XљR�6����(�5@�Q�+y��[�,�Dk�TF��K*���S�����I��(�Ɏg�?lD�[�H�6��%�\q4�D�0���hŖ�,p�V�d T��0ʵ2��o��a�"���!&��g�&"3�zҩh�$��og�|�vB��f�a�+VO)�Ɨ�*�� �תC
 Ȯ�N�M�#�k0���:�+�Q���.��|֦���bzB�D��ւ=)���RO?�[�#���6�ը�] ���K/��R�b-������w
��&<h�ey}�Z��}�l�c��W�{�z�zJ��a�ϵ�Sp��B���V)cbt�΢_�(��N�����؁�X�?�Y~��>|�^O���׭k� ��<p�x�(�%��u���>�㞩��_�f��g����I�.8�D�E�6�4,��;u���(z�UY	]|94�i���>��Ή�LS���)��M�S�M�[�+,ǖ��в��І�"^®��ak[��x��K7�dn������xd&	8��/se\������5�	��蘒 ���Z7�8z]鉲�����`k�B���s�8X�`*Iz[W2������6e/��{2͏Z"�C��/�_]%0�]��R�ي�7FF��]u�R�u��72�X�P���g4x vҨ&��"T�E��Z��D��@��%���a�W^�L�~(����%�lc�T!{���0��s+��Ss����%.f%)�l'��5'�y/�P̍�ķ*��)������9��m_���
d��yG���}��#�$��:x|�j�6U�Z<zItǧ�I	GY<���ެ�����d$Z5@va�K4���E��Fd�T")�C�Up�xc{q�z��io5�����3.�o�n5�����}"Tv����� �O�ˣ�-
�#�`�gVޫ|S���N�V;�I�s!c<ᄼ���s��(I�?��������Ę��
�\�d��{m�]�6$�>�*�0,��K���<AWF�J�{Qr��ZT �x��!���JEF>����^K��Ƨ�pa"[�^-�v6=]yD]����U��"�W��`Y=�p
J����y�fDY�-ř�K�$�"��r��/P�4�7��
��(~`�L,� c���x�E-4)�Em	�C��s�4�o�m�r��z���y���qua1��`Ƨ�74/T�΢ ��{q�<�Y_1��~��iWM���Jb�O;���i$��I�5��Jn	O����Q����J����U��v*h?fw_g�{e��qf�C�͌��w7ta�Y� ?���H0�ź��v�]%��]ӻى����Ⱦ���e<�Du�[��I������f�nt��ZA�*˻�w�Z����o��e�
 uw�u�	OAM���!����}qЕ�|�P��*-_������8���A���*��&͏!�Н��~�'��h��ίg����3|�p4>��� G�`��5�'zˤ��=��rh<�$6a�ٚ%��
�(��ܼ�TF��w���3�x�&[r�xޔo~��uӄ$w����z\ n�L!�ͺ�^M����m��a��;e�}�����[+`�I�G�����A5v=�;��Y�#���Ƕ�5Мz��$k]ȡu�*Zmn�-<��U�'TW�w:���4�"lZ��-�}<Pd�!�R�B���H�0Z�l�'C���o�,�?1$)�>Tt? �{��b�=�� ��-JT�'�P���b���3]O��{�d�
pSBl���� &����
��tbi�.pzv$w+��#fy>�tw	�Q���k�䫫&��YR4�� XR����C�,�ZF��g�K˲W*�Q�s�o	Y�,��R&� �%R��oG$g?�'.G ��"խ����`Trζ�IO��R�,������x S <>I�	�W��Ĥ�8����FK�ݾ�����.��5�����f�فз�-V�˽m�DH�eުx���$P����#�]FKOE.���G�[
Rf@gjB5vZ��j����Xc��?)�{�e�'���`o!9Ph���"���K�h�濋@��=�Yg�V�r '��t!c{�� h(�#ZZ ޟC���Pц��\@h[�לn|�{w#D+Y��+G�d�U�*�B���U���aY�t�M&lfy\�G���~
6z1~�,՝פ�f�����^�Q�`FRK��6�N2U�Z���\�8h!:#�y���+F�b���Ϫ)��K�%R�l�4�<�R��U�$H���a>��j��<`&S����&"���=:W�T�GGB����Np
ƌ6�g���t�:<�W~�O�Y�́�C��'��ЂV�2'�����UPh�8��&���G$]���I���Ғxf6�
���&���߁��e�!�M�7���IK�j�̛(9>�����L�iݘV��+B^���+|N��:��8���g�� �2���`�9���k��۝\�NtJV4t�O�3��%�f�w)AO⯎}�!w&������.JIph������$�֬1}@.����~b��a�)Q0PLc �=��R��u���O&>�eZ�h�	V\�ŗ��1R��ɰ!��Ɠ��uD���I;�)H�@�R�~o���QE��$�&���w���v�ݖZc�E��+޳�:�.�Ɖ�6��!�T�b�c��$.K(9��c���=����_|Z�|&"���dJ�.�}[q����6�a�$������,M�z���xX=F����	�߿����KޘS0Ν@֑/ �?S����D�o��| �l�G-�y>��#���,�\P��1�h��&�d�o���r�+����Տ��+����e=�����-�7^��Tރ�=�C�74���9���O�+I#�:qHU��V�SĜ<ݓ"[݂%���Bd�R��R+e"S�8$�w���U�Ǜ��`k�7�a��I
�'O�:<�se���}�_�5�����@�mz�;�f5��P�_�󕒺�sCw;Y�vM^<�)�|bm��`��p���}��',F���zѫn.�E0L-�Hp܇�N�f��m �����>����?�/��������轌ڐ�%��Csh���>���=E�8����Ъ��_�["�W��Ć��8�K��ab��v΍�M���D_c������+���t�Q�{�)!7���0
�a�<�����{�e�]�Ak�u�3��HE�oH��S�a������Op'�b�9/�I>M��t�'PE�]�l��C-���yz$�Wǘ����:ͬSh��s /ia��w��C�z����P���io��ĺ���}+�� �F�A?|��J�EiUچkZ��)<u��N#�k�O�8��i����M\@ɯ�10�f٠�\d������"#�+��op��|�+)F��a�,�MOҳ�
�U�Kx�Fj8ނ��WB�2T:Z{`���U	�Au}�F,�����So�d�!{}ਨ�M��s�V�ց��(ȃs�6r��.�?2���Jg
�q���Õi�bU��:E=r1B�t�JQ��B�:S���+��Yӎ��pIۤ4���C��%��)���V�t��{(�;��/>���M��%��J�>#���Z��o8@�FwWT4X�G׃0}�߂Բ����[���K��n���u
u��X��r���
��<���<�M��F��q2p}_e#�;2�Z��ߨU��_HA��?�k��?�P| ��[�ve�Ed&Ue��sE��;ci���r�\���X!dI*u���Rٖ�o����O?�n�����d~Bh�����,������m�la�A�q���w���AzfFW���^���!ie�\Īk���'����;�7X���9M�W�_��~=�5}k4��ŏ���;�m��+��g��-x��O�A�j���	#Gh3;���6��K���ȯ���oOx�^>|�Y�S�� bjF��
�<iɤ��ˌ��I+]e ���W�gJ.����0}RQ8m��Iʵ�)�f:�$yiTѺu�0�}��#�tE����j���A@��0�� �����PU��|OTYA�0������#��������ԄfI(�s3���\f���T-�!�P��(ߓ�V������ɀ�~F��-��W:mr��BsH���o�Y��G&/���3�����AH\�������8A��_��7.����C�r&C�,Y�D��{rEbRq@��0�n-Rz�����͝O�H���ETg��~HD��Q�AI�m�/9ʤ���ewЍ=ʈ���y|��[���Y�Xܦ	5Og��S="�)i�$�U�N�.���8zÑn���@�!�������`��!���|{я���� �~��-�ȱ/�}��h��!��p8�t�GR3!l'����.]H�Vs��gXX�����ş��Z☴�H>>���-�C����ً!��?H>Y�aF�a�A��%S�������i�Y�x$x�/��M�����e�� wV
4�$bˑ/�C���Q���i�{6�Rq(�T<�J�o+��շ%&������Dځ1�%~�\��}��<����x?�P�i8�r����&�8�8���
�j��b����;��eZ���m#�~���!s�}���Fa�!�xȡD��U^y����:NgD�eL0'��/x�J)s#�����j�-���P�l��p��Jɹ���%��.%�d�r��ؙ����^�0Υ�!��4��Tu[���$�p?(�P5��9�����,{�jl����<�Z%��al�梹|x�OYP{��8NⓏ�I��CUX K! �=p��hИ���@2�� �˃<�r-�_�U���(�g�V�����S���ѭ������٪Eo��3��u� �g�()$��;��f���H0*&�������VS�<7�Tu�������u�.��ʖ0o����G���Md�*~��0�%� {@%�M���@�����AEɘ��B�|a�z󌉽j�ڲ gK�R:�,�W�[�u~��*�i�^n�;!}A���O�Cn��oX���u������X�K!��4-EyzѴ�.Ǯ������8�؇�@�-/���]��um%�%\��j\K��2"��[b�.I��wp�M�{<��n�$&�����1�6~B��+R0s��x ��fK��/Ō�{d�ї���r� ?v�i֞g2�4i�tPT'���Q�|�+!�����Sf+�ü����0�Ԏvkx���C�v�AI,��*�׆ML�R�<���o� |�� �B�\��M#e� ��,R�<���EA׀T��Bv�x!}��)B�>ۖr�(�/�U?�w���:��+�;�B`�s���,(�&!�A��[��m%�m��M:���:Q��/q�xBv�R�|�b��?z�ku�,
!@Y�SZ�n�E����=�+9]Q��|��F�����kC��Ҳn��O���vV�k9�+;9N�폢n���$帵�'S�"��z��:���kKv��1��T|�Uy�R��]�mE;�����?�0]��������&���e�\�Φ("4Fngb��7��?�����n��,H/u���<~�I\)���=���dalY��I;e���h���J=���� ��/7a�mu�lH��I42ha!Ax����jc�Y~u������x?�_`���逮@�&{��l��ZR��/�����/#{ƣ`;O�}z���޴�ׄ~|���j�}�V���H������B���3	��`YZ,�RLĨ�s��m��7�o
�w�?� |�R�N��;i������$@@���>I��7 X�4h��)c���������֘k4 �@��/36���My&� oκ}���%�vY�b2�E�aYh�������n�$�MA�.Lf���kz^�J��ܷ5������֫�{P�J+��K����t�H�c����{�jm[�����@��/Q�Hϟ���#�ٷ�SqG��ۡJp�!��h�7�A��s:٭���1�u��0��B�bv�ψ�<
7Ǘ�A[�'�A�y"tl��f�^��ԝQs��ǯ_~c��S_O��bPB�;��!�����y��]���Gi�mww���Gٵ�U�M��T�ﱤ�+.�9���ԡ^�hF�<�b4�jg���|��F�lN����1T��;f�'�ѳ&�\�$�=��źD�7�;Ň�%�[��$�-f�Z#ص\T�$*�Q��
�s�y_gY)�Rd�<��hO�P_4Z��\tMG��ſ�.�Mh�����DL�E{K$�M���j��uή���Q�O��O/�I�#(���W�{P�p����A�y���Ĩ��_������\�Z�і[��$�ؔ�DI9�`����s+{fYI��N�\d|�L���O�lr��1���%[Z�۩��U�B���rn�Q';&�ҭ�[�u�Y�<�=�k 	���FC%�&mc!-�m�-S������.=bP���%Q=�[�V�E�_I�~a��vY4�8�3��b�`G@���{��A@]�be����b?q�����)��:�@����i�`[bP�;��[��s���F�Q#�� ����j
Ny���N]�G@UTa<!�󌿳���a�1�.#����p�3]�*�x#�~eSnE,��������[�n�P�u%�+g;�6IC����h�%H����9[fǓ2����~�$����	��ǶNկM��������*��B��=%�Gxu���G���䮰 ���O�T����K6�y�i�o����=��\'J[����
R�3�if�^��린~��7#�.��a]h�K�hA$myč���0L&m}��a#L>��u����wDE�� ���(�[M�Ѥ^+��5���iO�7iP���i����5����vn������;���N?vYt�X��v`�G���n�X�<>~��%����;��/:�$�>R!m�M��������9�o ����+@AL��m�{z�Z�8B�Z���Z��9l֔r����fKܧ��QojWB��댋���߷'�W����p�$1N\�F��1j���C�J��I?��1�"���i����䎸Ő6�H����N��i_5J%+����2��Fr��3?��~g�mk,Z�j�p��(�y<��ԧ�m��b���Y�L�K
�HKu
h]__����r��ԟ�v!uPS�t-)h�nJ8���gk?�l�Ir�[vaޫ��{΀���{F���R1��"��G�9Oô�JBy^
VRg�]Re/���k-��J�ɏ~֦P��GY��m������<�s�gO�<v�s�!rg�˔�Ӌυُ��}�Vv�U��u��%��M��1]x%K����0��
�*�x���/���41�$�q�C�5}��k�UƓD�=M�'(��gM�NJY�z�@�خ�f�
)l[�n��e��$�nUr��������
!]�N�"P[�X ��2�*<�y%K�*�m�(���U}�a���g
nr�<a�������(2�6�y���d�1�.k֡I�9�cPR���N5ƻ�
�ӟ�d쨅��B��-`Q�]aAG��q.U�J�����׀�F��)�0�ՍٳX���g�ؘg8�N�qO�Ǫ��`VE��'*�8Y�z��5u���0���/�U߶?�:n1U���O+l�P7t����G--�5��q<�	[o{Uܲ]HT���l��%�ҵu�C�n��S>a�c:�j~-E<�.�ވ���^�`�6c$L�`�tr!��Nk �jZ��)�%����[�3H��nH�۰+%8-��~*>�e'��;���(P��o>�7��JY�q�&�q��i�gg�d]3!�#F��k۳.}̚����8��5f�ۜW���x"s��\��|�d�ݱ�T��BuU�"���P�U#�;�1h��אD<�L>��J���d0�>"�ā:I��ԝ���vh[&�\(��}��1 �s��E�O��xͪL%IIl:������G��ܡ�ЛB�%D��ks,�Ġ��J��#--�N� �cF�$���$��hE
j?-�ߣ��~�����9�r��g�H��!�i!�{[�l�N�Z?�;�F6<#����/������ j��	���L)��NM�7с��l��>�����#��6�/kѣ�>�Q@��[cG��0�(+�t1�l����c~�$O�ԷvrʬxՄ�]� _���G)GjpS�M_R�������,Kb�̭�ȏrbE� �]��b���A��l'I�m�1�����>��_)�M��f-�	�lG֗X 0|�5:�P�*[���W�6���u��>��ꃔ��Ҋ ��(�C���Ƌ$N��h�ooQ,J��=h{���<�l�>�� 7�^u�d���=G��&��>{��2�����j�z�{�D�P��M �翽�D�,�hF�g�D���E �('�0��f��X�'�T0��}�q�|C��G�m�|�E��U
���ZE�����栭(�ͦ�� ����xgE�`W�`ش.�-��}���M��p$XA�6���̀��DD���\�Rig,��Iİ��K��<�,/Pݛ�߿�m�����A�uq�P���mK}�=h�-f�����*��	gUj��@;�#7�X�%\�\��|��O�Q��;C
D�f_	������:4r�ž���Hշk�\�5J���}�ֳxK�VgO2;��N���2\Ur⪕����m��x���X���o�Wcuw�S�^��'o��=�F�* ��+�O��0�&"�q�A���@�l1~�V�޶g_�dw?NK��n(�.+Ca+��t�>��{�z�-;�j���ǥ�E�_#{CA�-tmʹ������Y��q���3Ě|sLM��$�\u���ЛZȶ 
#�����ro����Þ��ɼexV��ߙX�����W�|9�O��ڊ{A\b��;׬ [�5 <�8o蝟,qMWK��J����>��u8��@E�h������N6Q�G��ќ�Di�Z�؞O�an��Mw)S.{P� Rz%-�[*����Ӳ�w.H^�����t��*���Of¾�[�mӰ��]2�U�.�~���J>�	�z�:������cz�)��g�sT�����8�uh�h�5���9�����������d��0�Nqj�L��VQ��l>��ȎʁP�k�.H�+p�J.-WS�c#ȝq����z8~O��y;S�{�m?��sі ��7�w,K5��g��Z\��>�A�cB�����Oo��e=>l,\)\F$=��}#��N\j6o�H��X�G�$8���+cY�� h���H�f��	�����a7����`����3D�ז�6{��tDBb&����LîW/��;-��a=�g6��U����~&
�q)ebՓ&�K�0��ɻC�dI�3����	D����r�ڽ�����җ��4�����4]�wQ��"Ī꿨|�"U�n�ly��.H�M.��5�l��E����u.$�/�~�YK��6hi�p��^�=�aE�2�k�"gg���ê��+Do��%<qT�p�A�e�i����r7��6B� ���\��&�?�^!����1�=ĉ�T�i��t��ˡ�Ξ���eE��n舃{gS���#'�?�I9ӦO��.�D+l��B����+�����0���L����e.������6,�ѝ��|�9�2�6ʉw��+t�6D�}�!d��`����X�^}���'	B��z�y%'{��j�Z�
�<���w��������>l�G�|�)	��U�u�!��u�* ��0/.��5��S���f��l@^V��o�VQ�uW����Z������5�P*L��K;j�`50�%u/�e6�&[hM��R��" ��M�@o6�ޮ��ӟ���
��W��ts��䒦��y��ͣ7�:�����/Ċn���"���,*��:�[j��R`Uw�B��::}H8��@�Y�y��>YL�cD����Mk�s�lD��h��<εqL����։��U�o-���̮f8��7�ps&���*2���8z�Qe��a��(���A(WK���i�O�`y}�7=�^ 1���p�4��C�n�z� d2ʾ��ź��&3�8�!�#�'����!�}��8�� �j��Ato:�E�G	Wiv����JwU7�D�8�̥	B
��~� �Q�-��U$�Wopd(�����?�X@.į��q�����V���f�s�\.���L�eY��i~���A��~׀��[��hUlF�l'P�(�{�z.l�.���i	�)L)֥L��`�@��H��=�)Q��R ��z��!��.+5�����`�`t�Mڻ����Y2Ne�.�~q;u���~� �_����d9�~d�X{J��3��||U��}}YX+7rn���,���H�[����&89\�DL���<�S�XD�L[��D���9��y�=`6��E��9�&2�hE��%s?Jv�	a��� �L�=���Y��_WK=v�S�<~�FP��P�~�6����Q��m�z�_�&3_Ԝk�;,a	�x��H���B�S�Yw�sL�!ˇVD�i���Z3r�^ۆ�E		Ŷ���T
����p��5�m{�e�Nב*K���f�x\(��D�߿xM�*��;��ZS9x,�D��k�bҿ��V�=|����t�*IP"z,�{<w�ݿ:�J�x��\���@Xci��(���%���rPO�R?:�^���S6
�2��Z�"����-7��U�6w 
ԝ��Qw-b�r������dW��!�MD��H=�� ��%��F��)���ܔ��ZD�,���1��Vƾ�<)�$�l�;�`��">&�'�r_�px
��S���	{���"�A���͐�>���[��L���
���(���qZP�3(�lsՈn�/���|QМ�j�NԽՍ;�#���v������ᒛ.P�Q�܍�u��>r�,�Z��r��� $�rZ94�L�Y�\p�][�H'��A���T��"V'	s�l�r�
��&P�i7��-	d�ĳI����Ꝼ�ر���/>��0"2Ƃ";����d��%C�����@<��3�:�i8K�^oc�	�1��)Cs5TһІGm(�ع��?6���w���1O���Z���?�������yr�:�i[�׶�+#�����T���y�ek�扂��#����?����f��}�6�P`6�RB��8��<He�6[Ł�I5�sj���M�"�{��L_�ړS1+F��>�)��e�jQcry/[�3��gMy�_)[�95��79�v+r0����i�\��7N_͎��t���ā47G������<� N�pNᬨq,�J�Br�i��eyqW8p1�p]�8����W�N����*�"�9�s(p��$*�g��9�Jl�B������Ĉ��h��4`e21�}3��d�8�j�ԇ{�����U����n��äOzg�E.��9[��T���(�n.�DlA�ni�%Ò��/%�U�o@:��
B�֦8������ehѭ��r"�4�?,�ౙ����j��	�J?���)��fL�[�� 8����06ꔎ�'��N�����|�(Sdr��ë��ⴚ�.Fl7iqڗp0u�E�S��z����c�K�N� ��� ?}�JL�"@��1���)z<��ɭ������;/�Qx�ꫀ��#a��P�E}>��)�I|�������`��n��+0VI�}]U��Bka�ǑR���g�[I�?3qթ�ٚ�{���Iw��ػ��F��hX�x_)/���"O�ys�V�&��[e���}<��/Y�2�ՙ���l����%{ZMٴ��+���9�I�V�f�ⴠ�,^�Z!ʚ��QnY�oK?L:K<uH���"Ԋ�v�!/lI7!z�ቛ~l�A���x�|N<h��� %���S����QOz%{�ð#�I�l�%����س�r��y-;�z! ��*�b�k	�	}�\�n�~𨿋qx��"�w��$��iBbs*�9���I(�LV�8��2���лE��Ig��F��W[�F�-�����l�j>ڄN+�u�D���܋X���
{�pTDU3�Z������.�	��YC�̧='j�����|�����	�!M�c�Hԁxc�z7`�V=,�ƛ
&#����	2���9E�������c���R�s��ZN6��,L��GF�j}*B�{�ݜ�
)�r
Y�����]f���j��/�mop��Bol)���:,�ݳO�������+{A���nJ[p榥/;	��y$������r�@�դ��>;P:p�܍�s��as2���A����9]�y����Şߪh�#'q��J���#���hv�P�	�`:��b���=�}��@���IS
yS�>e����P�]{�UP�fm��<�~��v<N�TB>�K+F�؋s|�����hpu	A��$�;P�7+k !~a�L\R@P�J��tr�# V�}L���n�FB�`;�H��0��c��W������BČ<۸�$�]�(}��W.;�zjn�j��
���Lg�_a6P����~{����K]?)	�g�ϕƎ�����i]K��p�quO	�2��gG�L&����އ�:�?���4ۚ�w3��*O��x�;��|f�=��A"Z�����$�9\-���wŌ�����Ťt{��⦨�y5�a�lFѲ
x��`�["��)J�t�*ل{)���F<w'��(0�a��Ġjy��#�h|
���ƻ��h����)�~Wr�����'@��e�#@��o�.������H���s�@��D��j�rUNܿ�Q(	�z�C�&��m��A�����^`�0����x���+@��&,3"�XU���W���B�@xq�X��Dc�I�;>������6����^��!E1� C�5�X��L����}�_�H�&v�D�g��K�ශ"�/��D	�t�o=�:�B@hFg�����v�Eo;�ׇQ�ѡ�(��˼M�A��L��i�E�"*),PE��(�CW��p����������i%�)xn���ߺn��S��ʩ�LAef��>B j�g���DNp^���dhe��*I�<��d��k7�brS�5j�1�M�$'kz)l��(|����b+��O>f-p��/�$�'0�)�m�*R�D��U�wQ��E��7���3��O���,�u�a}%|7��a��#[ڰ������.��������E���@d���_#߁�J+E�%PDW�y�eǃ<�,{_i����+��cP�p#��1W�I�����B�����.���c�qTj>|��!���|W�oI��-a׎R���s���mԵ�6������,Q��|��s/�����ƔM))-�V�5p�#n̾��w�偷���|o8�=p�>Ca3���v��x�/䫘���<A��ّ̇=����y{�8�6�%��Y���������5���^;QV�ڥ;��)��t�S�������'�?�˹i���QdA�H��`h�7`��7����K�<�r͒�?@r9�a�-�8آB
a�%������?g2@Հ5�P�z�*ALVMEy�'��
̎��{��#[h��׆�!W�hE��5��G���l&Vԩ�?_�*�'G5($�6��
�{FA���>O� �����hG��a�'��~�`�v��&��o�3їvik��"B8F��l��|\\�>D���U �Y� �[��ySzd*��9��f���C�m�Q�2�N��Z>$��s��%��( ����extw ��)�x�F&y��Hχ��Y!^�}*&����z"��P��r��w%D�傔Oq�k��{d�IMv2��'IF⏪t�QB���kq�������(�;��t��)gU7�������$�`�2�`�����qB2=ޱl��Z͖�a�Xc���{}<u?l�O��I��~S�#��Q���ߥ(�C"n���_�B�P��`|�c�Rg�|S����i��	���
�kC�����|�vI���]��O�d�7�QS�*��r�Z�<�x���4\��+��Ψ;�*:�Lu�D7�@B��x����>cq�W����Xo>�EZ�ܲ�.z>/ۼ����<�ު�4�\����P#?sv74I���|+�e�΅�H?�M�jm �h[�:A��o��wiO�3t�ל�V��i3#����JɪO�����rN�� q��^f1����ټ���c�(�ޘ�c4FL�?�K,u�%{��i)�� �|uq{��B����[��	�
Z��7�Nv�����cXߌV$�7b�ܴkp\|o�lY�ː���ΛwK+�����B��8S:<[����T7��e��`;�]�6\s��A�8E���^t8(2�ڵ��p�MŮD�oz��Z�Pz��#�%�P0B<m�1�����y��xɈ�z�\oj*���f����j��9���?�1��"�6f���8tp�1���p.(���`�f�ԌO�!
ˇ��,2(�:��n.A����*�cB�x~ۓ	O$\� ���?���#�v_�/WՃ��@9Wd����B1�D��hV;��4	<9�?p��B��d��l�}B"��>n�$8��t�r%3t��%\b�.2ݮ�!B�ȩ��N͎YH���\�Q��<s�bmF����/g����H���N ��Yy�?�.�9������g:�=	ŋy�pT�^����XD���ж���nJ��9���7<��nƝ��;}|�W����4� ��?;�4�z��5{��)*q�G��(1�!��&��Ki'�-Lt�ć�h駄���[�|(����Lae�8�͇ �V��,�ǒh��5럫�#ߕv4v��Ke��Z�-��S̞�{'�t4�M� �����x����(�U�~�.fĞP�X���B4�W�{�H���͕�*kOlFP�I��U��U�WZr6��FE��eox��C�M"�N����4�O#
G�)ؼ`wj��8j/4j�b/�b�gd@F���2�D�I�oߵɠޏ�+Kb�=��v��=��mS��)�Һ���sz3
	����\�����$p��c���䌸s9&�M��aIjd�c%�\3��,�������-93���f@�U~�%(�Zq��(�����#jJݝt�8���r~3�%����"���p�K�5�Q��F�X�\[r����V,q��4�W�$�ю�>A��x�&V��S�d�����$�;�b�F����c`'k���]K�ݭ�\��,cF�j�l9�e`lqE?�6�MP�_ή��f�u.3a5���DV�3V<������@��1^�_`-uo4<*��QJ���]�X5y��;�G�f������#O(�����e���0�oDCf;-�&�-�wg�9�5��S������8�%M4���j�vy�X�$�!�����)݁1��u(�N��$���V6k�S�Y�:��T�)�CoO^����k=Do<��r.���w�ɠ�3��D�.C�}�Y���lPuR���������՜'��X+v��<�{�QFʠ�y���r��U�P�+B����.)Ӹ�@�3>N��nA�a8ﰯn��Z�u��{̥�-'@Ee~A�aAAIjU��{�7����B�"��-C�H	__[��1S����y�PE��"H�f[[�'T"�����r�\̀�S�*Zȷ�����k�dR�C��vF4�*V4�|"M��/�Q��U�NǪ�\zy7}�L�҄a8m[�>��=] $�a �l��͂��>�FR�T6Hq�b@4F:1T�&Z�|��1�=N4SX���Y��Mr�(��lf�\��r���P�`�
��7p맠��Y������ꞗ�d@��9��8�4<O��,���>Y��cX��k�o˨���F���e5�[��m��b�����[(�d��ې�� � ֚_	z����������Ag[ьh���;H�2��g��!@�fN	�?��8�.�A֣Ք�w��X�\bTH�/4�9��Dp���,���lu���]pqY��Iz�5jv�����m���l�%VT+w
�"fë)3^�%d(�h��	B� ԰ߧ�+i��u��L+�(��<:���K���[H(f<��D���,5i�Cj�����ȁ�Z�"�	EQV�DZ��	�d�[K��ݿ Ž rh#LT��E�����l.�m���$_�`��`j�v����{���Ru�{M��������859��дQ�ҙ���ź��q�3�'��M&X���ܾ����`U	��7��=��7�W��cl�sAv���n�hk�:�e�ɧ�&���Ε������r�k�Ƽ����&d֗&̗h�x��]���3U2����(��+�~Q�i��7�x揘 �T�%�ޅ?�_-��J����Af�z'��+&� ���p�����eK��g���P��7.U3T��m�4Ǭ��4eE{�B��{/<�!�_�����8��,�%��1+ �>s���y�6������.�o�������[E_axMf��w:Sz:��|�,�Լ:���&�x�a�;�P�$���B>�-����Ä���sT���P˼�*څ7%��X���Տ��#�v�9��?2B�<�I[��"S�)	{9�k~%*�;4PV�	��y~8�:���n�����&������@�ۿtn�*z��'1�#k�wBFA��'Y��`��).W��ܨ���r-��f_��,ܲD	U��K��U�	���3�c"���c��M�x��oB�&�4#V�x?@��K'�R�)`����٢皣��g�^�� uрa�9|�k�io8�+��~7��ŀ'���Φ��>.R��;-�#�y�I	]�ԢV�QM�2����jӷM��dsA�Nvf<�%;ØȰ�sf0E:+�ޕ��x
��]]�R�N7}�|u�G］ÿ��v��zǳQn�����HUڅ.F�NM�$Xw���\Q ���D��~Z��ݳ��[ݚ|��-������'�wǶ�d��;D���	����$��x�,�7�K.��;��/��q�v�k� �Q���*�����2=s+�"W.�E�Kb\6����5*�����&�������G���1��7�����i�rEr`|����+ d�AiB#(�^�!�Y�
�2,.�QIp�gJ�����o�鰜nD�b����M��ڳ]�����x7̜����x=��F]�`�g�zNd�����v�
��5�7��r8���B`@Ϳ���9�����W)!�5�����K�~��	�D��F�Er��Whf"M2��6K?+��k>�{?x���=L�;�#:�D��j��>���L�h���*e<L�!�}��*��~�v�(��|S�`L��r5C�n�4���b��0��Ǐ;�m�𧍱f:����O@�ڂ.���.���2ޝ�ƍ�A. ��FnH.^$�t�%Xv�i���d�n*����Կ���6xz���(+����e��
�l�W�t%+�F"v���,IRu�~�{��DȎ-;P	�#b��_9*�)6!�����$�Lu�6���(��W��(N��@�� �5�6�A�4����Y�E'���PC�e�S����͂�K�u(7x�q��~\J0��>���2���J�~k/��a+����I�]}�-c�2�Q�Ybq�����,�G3�7�Ek(�$��֊2�r˫B
���^���	=��$��˲�0�mWO1T[ڄ���d 
@}X�c����3�x0t�u����;�Y�o��Hh�A4}
���*�/�^_�93�$V&��X�tTO���9�6��4�)���Q��	�+X���8ఱ�0�V�]#QPG�#m�T���a���Εy3~�׊��1퉇�����68�����^ET���	��F-�vGE����M#������2!-�I�!� �����\�w/_���a)Q1�����2��z���U�ԭ��Mۅݪ��[�)�9�����*��#�����w��Z�"\��`��ұ���a��I����5��揨��%"_��K�Y��fa�$vWu�k( ��;D��g�����F�	W�����}˯��j�x�w�Z�沶ʜE��,��������3@�}��UK�ciu� C.���(=J�C���a�![є"���&����ʃ]�@�0[c�7r(׿C:f+�	m��L�ԩ�f]/���]��^b���$��"4m��~��^T�����5���mϮd�ɀ[��W��V更ٙ�y��W�:x��|�w�W�~^�*d��|�1�s�ڸFM�M���z_�/7���i�wW)�7)7aΨ�2��u���ؓF�k���t�\��R�bSC{v޻hsY����,݄s��%�}�VR�L��!�#��eWT:?#�z��Z�xE�.*p�ӭP�M&@=m;�q�(�Բ��D��8Svw�?b��s<���g��O6� �=4_xi�
U`0" �ӡ����p�!8bJ�����DJ�����3���K-����12M���a���iS�p���P.x�,�{�|�))�-h�&�&J4��vTwt��_��5�(�T?`�`���x�]�I0+�|\��$C��j�z 5	��%X��i7���M���P^�<���# F<�ӹ2~���߲�N`�IS��I�gPQU���n	oP?���Y�X��GE�J�5�dLC��d�m�D���X�0��O+$��Fٴ���]�=ｆ$�]�%&�����9���e�8J��k��D���'�L�w�I4R��`��Zf��#���w�D
�p Ȗ�A����,��#ɯY�M5��IW�_Cc �4ҊH\�x D4�a��<1EVô�n��B�' �2���Y���/l�Ϙx@�^�/!�-�9hB�_Y��s�M�[�eDn ����x�M p�~G���4aqጬ�W���d&Q�c�o�R�p�S��Qf,�������2Y�ˑb����k��s.�>�Xw�S8��_d�4o_��m�D�uΐ$�B����E2�G
3���Z5,�7��U	;�+�����$���I�G�P?.�jY$5=��f�\��Քvv+x)�|�C��T��ѡ��s�C��`t��~edŌռY�f�V��b@^ǖ���v>��Ǣu�A�=s]��5N�����`F�.mi3�@e������1�<\��d�߀�o{�����9�A�W�F�� (<�h+l遮�f�j=6~k�y��u)X�0^���A�,��'��v��]l�-����sv9���\�B���rxiA���U\�.��K6�����w�S��a�&��� WII��ϥ�j��q�:|�i�G�6��$�e-E�N ��8ߞ 8�-�j=�arY�;{��?ݑl��'$t���l�̷�v���S	T7�Y�:�ݠS�VTC~sp`�j�w�>��a/vw��j�h0��[1�??}&�h�y�=�Ӗd�ZE\�p�چk[0�L�]��0��)�f\�_���*��;We,,�Quc�#���I��[H��+��& $�4ѽ�A^�����'0fH�=f?�@������.�0� ̙0J �pe 2�u�<�\0� !�깠������p&%�ۋ��r�/kT4XD!�+R�c0�i������OὨ���8ϲ���An���ZFp�K�.̠��,8�r��˂�4oC8)Ce�`]Q��yX7��j�徦����`� Vh)pg)��bl�C%kP�5E�f+��H�ۺ�cQ�D��-����2 ��-������?	#,�d�jFɏ��?ccDoH�2X��ӹ�B��^�sʀ0P��_	\ϔ|td��,��~�Јs����P�[����A~��v��s��[�)��֒5�0�'�c�,m�u-���~y����J(����B<R�>�)�߻q���;�7ǟ/y� �����4!_�����a�ͷw���G�y��__��V}NHӴ.�_��[�z(����ά��b��H�C�=�s@߾���m�(�<��*�Vv�n!���?�?�n]���:�����t!ŝ?��W �[�Y�ˑ.�zf���2(UO��p1,�O�7�SA�y]�Y|�	��8��C�qv��)��nIN�KB�b%L�r����)y���[�!=�������H�~��i�?�ߑ?�@�5k�bW�,)5�Z\��Y@W� K�5��Uє�:�;��L+�v�Ἧ�#���F������]/��pN��Â�%��=ڄ'Պ�,��O��J��c�4ŵ�~�Ql�P�jhD�<�u��ข���/:�V�H������,S�N
�(!�W
�R�ɑm��9C����B9����2>�����l�D����}���a"˒3��A_8-`��`LdC�O�	�"���Ѡ�bu�6̠�V^�
r8�^<}��{�:�̀�9��b��d�־�N@�5��.
�+H!�[:�l�Y}�j��a�m�r�5¬�_�e�9����m�u�Ø/�%��|)R��,���ИE�T�O=7� Y����!�w^)�A�����>������=i��S�H��L���Sڧ������ F�1���.O��kt�����.9��/�,�D��	��t�;V8<o��/�G�c��q#ɹ<r��_$#(x�p�o��>!~��7���a�ޚ��z.qf�|�)\�y@I]�n��]�äŕuDVI�ZU�6=�^MO�
߾�	t����y
uwD�$��Rr$q�8qεJ��x��k����\�V�Mx�޲�󭺛B��9^߉�e��YfrE�jl�*��>O�|kX�cP�al���s��l�ը�ŨWE�-�7��i,jÌ�u�"�ԡ�Q�E~5�f�[��\���.��=BUV1)>z����VQ��?�2y�ރ�h�i� !s�XmI]!KO�]8V˵�z���_�k/�V:|f��KqP �ޏT�]P�M#��kpQ���SYu ��@\��P�]�^T�axAÁ�����[?
~ �2Dn��X��������49�13�j�̏K��T�g�2��WĪ��P�5C�B727��~jh�ⶬj[�xx�C��g��#ČB��';<$Dv�]�Og',cX"^�����k��c��y�A
W�=d`��L ���o�]�ئ�R���w��N�TI�aoi	' ���]N�,/>AU���WͰ�H�L�Ͷ�����,uK5�����$�\/��t�0j�\�U�+Ϟ+�hj�ҷr�o}F�0�.��ܹb/F��(w�{{đ�L��7��`�*gq"��N<��Fn�ױ̶ut��^��H�T�6iI��[��π������̳Xy��筮ڻ2���G�04�t����~j^D��2�N�|�ͦ�F�.V0�5#�M��ϴ�h���J�]A�0�g�/F!&w���@�Ⱥ�0�I��"����h�Uvn�f)�w�a�8�N7�7�$4�����_<����}���Zf�Y7Ŀy3_�l�˥}��2.�k��z8}?���s���Ix�0�R�zZ*NeD˭�J/:���`�933�Ľ�P˫]15qR�X�7�~^:��_R�H��B����=(ܗ���u!�7�f�L¼��+~��(]��w�Iw�sޜ&�o���;����В̈́���DW���@LXCA�"P
%��80�H+.�]%���ݦ�h����#�.�f�/1,`�כ�&�v��s�	cU!=������3"ϵ�$$�����(�pz��
 �΀�)�O�̇&����v��c�l��mm�Qg=9�%biTL0w�i�3�����d���u5O���H���%bF������W��ۏ�.��sPJ��@"�孹Y��'h���#2�����9S�~:�~R���	�U�ʭL0��3�3��Mb%?�}�.hh����1�>w��]g��(+�����.�[ٮ|2]�/�B;���7Ce�阔�o>��!��+���>����)�	���6�Zا�������nN=8~�|£wH�Ƅi5i/ ̓�H4�g�|)a�+^��Tw�T��ð����F�\��P�����MYN��(p9���a§6������g�o�
���
�iM��i���CB�Q��zB/���r���S��C�
{�f�,�Q��3$zR��,��	�S2_A��n���?�b�_~���]e���%l���w�3��b,@X�W���=�V����Y�ݳ>ȃ��k�e�<Ӌ$�(�F[�A��zO;��n&���c_�A��ɵ�|���m�U�	��Z �����k���� `���_���"�"���0Dh��VAk8���|e�6FBm��O��"�%�al�)�U��h�ӡ���LY*��d�\��'BF��ȶ�����o��z��I� &JY�ʶ�����&*���E:+"F(P�<"�4���`Ox� ɳ��-Iʌkjm��i�����d:�Sw��prI��`�b��0؆h��ZQ�uX��J��3&�3�݋���F$Z����]NJ���l�q�5��͆O�i����A�����#k����vo��	��M<��j�~�Hr����V�s�|�}6�PŚ���;�mW��|��Ǵ���Br��w��k�,���P���}���-O����hP�+AD�������c���UyB$�5��]�*-��	.� ��Wx�M�Q�����s�M�P�+eQ�+��]����"�h,�(�����FM>��j�����5��`�]u��MA3�������2s��vX��xX�G2r�]���$�:,�N������;*Y�mP��|���wo�&q��PSFWc9�$j��~��,�邱VGGb{IV�qq y�����0oi��ZU����UV�jp�W��Aj ���	���-�̌S\����nV8���_P������*��ܝ�s00������{?Q��X�uC���
��4�s�Y�U��:�|(����?(u<��v!`~��I�xx� p�ְA��.~�;g�I���l�{[=�\��+o3򆲶�ͽ�#>Ar'���JC�el�;Q���3	`��73�v��%�|b���KPMv�zG��PrK�©�TJ�7���]���/{�N�8�zRn8�{Q�:S����Ү{�DY�JQQ3��~����mP�C2�����Hb��kL�g%�qY�U�a�mn`S����<�U��o����� V��u�A�Tw���K#�A�麼S�v�%���}�:�B�;�?�?�I�x\�����7���}�|�yL�{�rb�H�Y�,_��*CB'Fi�{��9��Mƙ?�3�Ȗ�0!Ye������L���M�5u	Y�^b���Xh�5��cm2��ӎԳ�ބb���/ԏz��gL�}�m�j���&sE���ӽ'����`�U
"j暴�M���15bdь�\�گ�+Œ+L�	\Aiʪ~�s5@7	��I�0��yUۧ�X�͔s!��!�_J�	��~\��j�j�����1�ۼk�/�^��2}��
�!@�3����atCt�׃��o��J0�0\ZWi�Q���[|i9�R��6�6�����]�� V}��u�a�]=O�.�ȲЊ�(y2<I�9�$�(�E��|��|�w2�j0��q��?��'��]�M��ּ��n��s�6�|��C�󲤇���e����Q'�����{:�8o��!�ʿ��vlkd7�AI�5��pU=z%)��Y���l�9����y�{1��j���$.�mC"���+\!����ǫ����8�T���r���H�d���"�ֹt�	Q�%*|="�%�M�0��D�i�>V��f�=H4`<�σ��K+ ��$�'�ٗ�&�/�9k�]!)��vT	�34�n�=�S�ri�PB}��1���I�~�B�� �y�a�tN�}�t`I��ˆ7�3z�5m4�q���-f���{�Qd�c��X��a"n?��@ǈs`�u#B���uJa��!=�Z��Q���C�)�i�[�����xV���.��Y�դwlт�?�\��TƤ����1���]�#5o����Xj�YR��I��F��= C�K!�v��@���ve�����&�tw�P�;w�ݬ�Y��Ұ�>��9\(���Vf�.��E����R�6��$+���pjxo%�m�f��ݼ��v���jt5����7nx`�(�H�X�R��[,'�Y,��ۆ̊{X�ڣg�}���p��_��X;�>BU�p5/������u�֦EhVn���|9�5�J�L�O����#&�j�eg�:Ӂ��	UF:d�gK!��$/�����J(�5ak,�E��9$���{�E���_w���:��u���a�_�&��UMiߔ�^^ˋ�k�@�v�r����̙���n�T�s�+�דa˟G�zQ��@ʨ\����s�kK����~VY�/���r	a���iJ�҃̎!𔯂��K~�;���+���]|w��+d[fmK"�(��fGJ��
��*�I�E?MsJ���5,Ҵ#�O�y�)�Gj��E��:� +�}�j�!����4����c/\��D���I����H9��c$jpb��,��̔%5�?��c�e���>��
M1[-�u�-�ޒwby官};n���e<�d	6HX������B��j����?jH�=h7P��2�zp*<��n�fA�
��&�W��z��5U�+�>Q�[kh�=Z��M�n� K�UT��6�*�1�l��>bRO3T�P����2����[���ʄT��	ا��� ��*���3��8\��=&�˥�������J���d��~en��2^W܃x��>���)��fi��h}ϖ�'�������=Z��u=���9� �&r�F�#����RwR#Z���Ӌ�����Ҳ����[YԈ>u��Tnрh��|����,�џ����ݒ�Gn!k��n������>��T�g�veLhl-��y
?�;�J7�i�
	{+K��@�ȷ�T؋E��P�1�:�ז@[����Ë�J*z��:��,Q7u�>ag��c�B�RW����ã��q��dPb��REJ���\l:(1d�JMi��U���~	=>�Oӿ!�5����S���zA�M��2т���{d�,���3��@�(A��&���7�)/c�Q?I 8�}yoVb@
�iH�|��t=�סPe�ԙ�+U^j���TN,*?�';�&Ć�	����x�v7%�&��׌���?[��Dg]��ofy�����)�Z��J\6R�й3fu��2P�_�����\�w e2W�zGs�`�D���z� �3:���VbK�B�?݇ �N��y�=QT=#�($��O0��^�f�N�"a�4l9��~<�M�g"ɺ���īU�^��i@�r*�nE��ᢵ�u����%cD�ذ�M�����S��_�y����p��b��-��._Z�yEo_UuG�ϝ͞�3JtS\1$»G BqYe��9��nTʠ'A�t��Qb�EϜ��a��i��
%���_�v�F`��y�i�@iw�?� ��
�������%^=�$D�������B��q`�?���o��#���y��Z�y���&�몷��N�tJ7�#�57�(�|
@�(6�LH��s��s��R+���Q�d���|�Jd�CG���6J����Q�u}���$G�+U	������fID>�!s�L��$}�$�c8u��'�&�@�H��'43����T8M��v����/�����|2��J�b��c������x#���#���x�IЩ�Xq#�НPE��"J�:N�9-��+�|!�a#J�w�_�����3%��%]����0���I�z+V'�w8+�2�r|��s��Ӹ^MS�Nu+�]D	��s���d+]B��Κ���Q�z��L����]�y�fb�m��`�+5J��=����0v���l�n�W�&�NK4�Gt'��w?�v�Ӛ�;/�ʂٸm��a&���g������[��.� �1���(�%pe�@V�n����8ٞ�_�m��>�w�+�U�x(^��z_	�C-����}�;�%s�G-k�Y'�$�a�s&|�O�O��>��5�`���_���;<)�LHA"|����+��X}K(�S�T
Pజ���h
�4WL�[ջ��bw��Y�~�������l�d3u1���%0����������hg`-9.�_�vqӎTA��?�X�=^_�L��&��{���r Q^{�y�Yu"�+e� �PБ�ؑ��+�7��d���r|��?#CR^.W�9<��0�\�v[�s���E�Fն����ב1�3!7����m��p*D��ş(��C��<�X�"������T��ŸJ^O��Ol�&a�-��.��-=�fʖq�3W�~L���QA2W��͙�����v@���e�N�ʆ��I����wȲ��"�RD:c�e>�N�?"����51S�1��<Ո�tߟt�`�)�M��ז����b��C"2��a�a�CX��[��O���>P{�G�:�+x*GL1����?O�6��	�q:��u�wM�Q0���J.ԧ���2��揺=�(�=��q�<�Y���W�SY*���=E#$���ֻ�,�����۝ᬼ3�Ml�2��e�FUx��D���D���<U緸v���� 7��Lý�G��u�	���Nn�"�s�@�I���>�g �����e�i#9F��Jp'�j��GLC���Z'%�a'>���FC]��s��;-�(�ٛ��r�~��_3.?�Z��i�!�a0Sk%*'ac��;a��} U��}}QҊ92�s,��ׯ(���;8Y5M�,�}Ѱ�L�H�����N�\ ��kzd�̣���Ž5�����qq&��LaW���]�YZV�#U��?�u���;ONG�B����������IN^0���[�1�΀f�c����"ۀw�tE�4:j�^�n^ݟE�¿K�1W��uoi��.?B��gt���,��7�N]S��H'x�Ϗ2����dW����?���<*�\ۿ�lj�>�vIE�.O�{M�J?z�"�D��?�|t{���4��+�\Jr��3����ɚ�	����g±e��k��S73��ir�Pڑ�8����K��y_�qQ��I��m�T�T�hA�W|�d@��8)��)�z���M}�%�H�$���ŉ��%p}UZ�]U�rKVԪ5�=�| �#=���,�}���f��M���&��r��Nۮ��\����?b�$�;�t*��	�c����%s�O�ؕMY�.�l�k[$�Fu���Ȥ�S���D��|�{a�YgP8d����N|RR���3�b��B���{�v�M���r0�m�a��R _�i*���V/k ��t>znuϳˍ8�;�y��Kk�3��W�x����<�Ti�名��ʖ���U$QՉ�0Y�=^���ؿ��p;Eax�,�����	&�C���v=�9|�͒���E�>��˅��2c��F��뿗�T_����u�@/,��5Q�:&<�kEj0��8o��ȸw���l�_#N�K�DT��%�+4^B���<�!4�J%�G��ih!�������4�5kp�d�б�~;7p���\9bX|ӜCw�����a�46���j�9���]���H@�6�n�+f�@c�l��Hiz���R����d�[ɔ����OD��sထ.�����}f�@g:ѣ�k�,�S�;J��M��n9-�{kԺv�^�w�ո4	�����%�TQ~Ʊ�M���������'�"`oL���x����:@2�H�N�mO����{���~���*�{�5jc7����8TE~Pz���L�D����陘4���$�t���9�ydW���?�Z��xO������%�bB�(YW�R{<������3�? ��&B!?�W� S��n�_١�n��9�^�����@xpo����[�~�%���ۯ���[ci�aX�aI�X�>E
�͛��(͇gC�k�?�����.�	�����������6�K�)i?����A���3 <S%����	����Fߡ�6�鯆w����@|]2c�\%8�����"5�ֈ2�,��^���7��g��q��g�$��`��Bc�q���s��Ӣ�������+�A���x�х�`�6�~/�vF
pK��[���A�`�2���`Q� 4�78W2�t�2Ʋ��Ss^���R�K��!��C-�p�;�{��g��x<I�i�p��v���&2dۣ�ь���)���v�qE�.ȭ% ؐ����Wx�@V6�^#7�~X��g�Y?�d��c���c�3J� z�y��������${�!'n܎�3:$��x׹����d��2�I�P�6�,� �`��ͣ7��Bja�<�L���wJA��P6%��~%zi�	,&�� �:LV���BU�ȩ��C-�Y�D�c]�׌"�#��Fŀ,â�8A��gͱ?g��F�_�����C;����_�IMTHX���Eu�����[�O�A�5 m�`��迪Ȥ��t2/s`h�[|�}���H����`��J�Xs�s��-nI���
Y���i�G֖R��K��]^��'<�u߆��H���cRJ×��А�'��H)�H�a{�K"�΄Do�r/�":d�qoL�V��q���β�M����&���&z��oD�)�sн�b���zh��'�����5����a��Ʈ�Z`����͙��X��o�R<W0}�+8���H2�"�J�أ_���\��i�7f�#��8�:F���"��O�*���I�'��`��;h���)%e+_S��t�C;�>�*�ξu��������;�D3�
�K*[�h0�����<�����D��πI�򶒄�t��V��w���o�X��]�\�$s�ilCvL�|�1v^?��|�fn��'h�k�Ѭ�]�('�N�;�P�=�sF��pSg���}!�p����+)�����k���V�{@�o�f���*;�!S��$:��%���d&	P�j�ң #d�4�i*��Y���v����"Yc�X�ȅ^GC{"��T!������G�{�hy�:�ⵆަ�zvkAc�O�b@�#�ó�}�<����!��(f����m������J�Q��괇��������Dr�9F��4Պ)JB�s���(ĮIq�wV�8��d�ߒ�P&��O���!���8�y�60�o���B��VQBl��R���tZ��5�JNJ�c
��pOx�����Ux���]��!�n�s�S7��6UW"����TR�lݗ��![UV�Ľ��X~%�Kj����*�I�<��؏"b�~���t�O%^��ߡ�3���*^�B��P�|����8��˵$+�+$�p	���`Q�������"��LY��]�O��΍�Ц�I�φ��]�y�����7p%eSM#��ڗa�o�X#�B��Զfd����z^���ax��@R���v��y[���h>��n^��J ۲�@�ʌ��c��Rz�Ѩ��:�v�X�\S0�A�8�R�S~�����[
�^}���"�rNd�@ [��R �8��6a���8~����ݥ�6�����j�c�j��+힫�i�K4�FU��1�qCE��G������.�m|��.v%���������dkZ
�ΰ�)Bۚ�|��|�W�-�:�� ������`�G��|����f�*׶P�����M7�5�u��kv%n>J`�4 �"�Ƹ�D�Ru�NJm�[��ߟ[��ݛxa)���b����|��4L��A�)��y0�h���"z|�����`���=�;����P��g���X��B-���1�Y��{Il��`�8G����v�9�]�,7�z�\U�UO6��\��[�<W��((�i���4aH�ߛ��x܍`>���, ����w+M���AIi;�Q��)%;8���G\z���<Z`��M���t��+�Y@[�̟
��"��,@����� {ߛ�b�)Kʦ��1}���"M�.?dr�>�]#P13���jZ#��+:!����y�Y1���h�/�Й�j��O�C�A&�L�w�"/�����2��6\�'_m�!�B44+�l
�ex� �_�����#_`�Vϯj�B|�?G�\=�(��z���c*7h�rq@�L^�Uݟ3Б� �2"�%ٱ>�e	)�x�v��`x��� \���/l)H�>����3+S3��~Y��V��x���G�-�bJ��r����"�M|=V`��v��E7&����`ԁ�A�p�^w�7ː6$
K����r3���Z�n6
��<����Wa� ��O�`�h�k^O��-�_���a��~J�B;E]537�/*Cw2�~XI�t��F�G��C�5��&����Bj��*�1jp��i�ݮ���|^�S��=Ч;�ȿzf�}�C��R�D/N��jbC�4<�@�8)��_���I��pϠ�^ֳF�)��`.��p�o	�a��8E�6���4�h=�]�`��T;j:D��ga��d��_0�q"����v\�]�MA�?!&���eTa���!���R	�����Ⓝ�X�g`����T$]Ҟ��j��]��񳅥�b��w��,�����۠q���L�(q�)"l�d�%
c]�@��������~Eى�5]<&[T�/��0ɷ�����^9С��,ǋ�$w>$#�eP a=kI�[p�1$�%�v��Ń���aK�I���#M]��1#`@$۟��"'�g�m#D�"U�c��ҟfl��"����{ �HR(�\*��6E��17Y�P���M��L�0��"�K��U�Z�#\5W�>d�=�F)�$��O�,c̦ 3?�IT�P�����	t�M�����~`��e��s��H�ʑ"�q�W���8H���]���� ���|9�2+�1X���A����V*Ay�i�b�#��p�\����+��۶k�-_�@���i��.��^��ٗ�Qx����9�Jg��M�:s��w�X���ġ�W���3#�QY�?�M����������5#tM��C� w��"T�����`D�އ=�#v���r{�>B�O��%8��!��N`G@V�8ߢiBv��԰�Pߞ��7�� ����� ���(����U���۶ZBS-��TG+�`����q��Pw"��a�t=h��Q�Nӭ���T���|Q�=%,�1u{0��j�N�6#8x�s����!�1�[w��,d�M$˼J�1�i�~����1�1�=!H�U��jo�n�F��!ԉm�*�T��C�
�����}"��(d<i���B�R�ǝ�$N#}�W��H �UiҔ6��v�c:��-�����BH.f���Qڽgq�(���G�$�wMq0�j!�u��ῐ��辄��Wj<��PZ�v{��)P��!�eΊ��إ�X�s����$�zkn�����ϏF�>�g%�`�(�,S�,Ѝ�2�%�=���k�D���L���`�N�CE_�_�c�b��U  �{�V�Ũ5��)~�ok���X��t��᳌������D��m/]�ك^��#瑾�@�~��'8��9��)J��8��*=�#+q�Ƚ?f[:�nҲ��Ar7m�{�"U[C��Na�?��Ʀ���D��rL7{c'��ʂ&���+m6���nKJo�G�=R~
J��K�_oE�~�/DN�j��_��:��h�0��:�LΈ��	��n�*t:"dr���ȫ�"S|�g�^���qz���Y��b�*���
Fn��Ȅ��}E:Ŋ:��/��	�ݴ��m���Yغ��9$�h���H	j�>�qni-�Lqn�,K���$˓�L��6"y�I^�ԁ�Z &�m!�u�\V��/u���_sU� 4�82t��$@�z�o` >O��`A�X��7��'F>��yfb��cӥ�f<�^E/m��Q\}��qvg�ae�����/�����(1r�-TA������K��%v��8]rf����'?-�mZVg$�>g�3(}W�B ]�3�P}A�X�[*��8��Z��B=蕁_I�F��EV��kċgX�������.�,�0"�R������5q��a�h��A��Ģ�\*U�̹��B����f�+�&ʗ$Y�#X��W߭�1�y�������&��t�s�Bm�)E�TK����Bc��f�VG2�����Ś�M�݅Q{�ܤ��64(�F��/Kc��?�5���ф�RLu 4wié����wEІ"���g�P�#L���3hU�\�D�qE�/c��T57�����,S�8�
����Pk!� f���4�f�YsL�(_��m=c��t�a&�੏*H�������o2�Fw�u��X�ǿ��Ay��؛�ݩ���Rh80A�č�<jH�Z��Z�p��M)���|�M[ �9��n`'�p���դ.0�Ė��df�b�;�1���5��$��q�x��Wh�h�q�ښ�5t�mx�\�i�A�&]��iw�n����I��/�@C�=kk�璢�"�Y���g7X�J�4�_R +(�O-�f��R��)���צ)����~�|��>��8��kV� w��#9��0�	�،y��l��n���h9�f�ʌ��w���UR����V�}�êb�����I?\���8�T&��߲�bd0%�y���n�p��Z��VE-���WȠ�>�t1�����p,yA����x��^������� �9�´����s*� �i9U[�B7���U������"�L_�EX��w�L �v�8 rKՉ�ZQ,%�GZZ��1�L����v�V��Ƣ��?T�<�&g�"3�%�y�s1��߲�n�R��~�b_��Dy!�܇GlB�%RB�{u�Z�jF����(Z}�T�{p,��9������|=�\�j�o��x�EI��mlq���~����Η��NUj�_-�GS	�T9��1v��<�~�[�c�5��{�U��)^@�$:�����©R����J�K�	����ߑ�'������"k�{�$y�~����o%�Ȩ�:Z���+H�U�(��D�K�!@��$�4���5��Z�Y8�å�=��ӱ�ִ3�G���EI�<�?M�_��	'����Q�U09���P�iC��AJ�W=�y5�l�X�mwq��'J�"!GS����'��������M��W<�V�_���9����`�je�=>�ؒ�vD@N��-�/��Ʌ�$���}�����9�%���JNܣ��m{r�rU)��̕���b�d6���E�g1]^��7��lq�/�.D�G6�?�)�����t?.nX1��ܱ�Y�A�gz���*R�� T%�M=��y[�l3\?�(��Q�j�����b���ι����9�$�詉 f����䟭�f�����~i0iu��������6x.lޱ,A5>�ͩ=@�v��B̺ ���2�;��5��ɖ:eC\����]'k�&oF@����%���NZ8�
�:��e|=�5-���x!LS�3Ii/��xXtF{-��'8wW)>yB-m���Ș��J#�zMt��k�IsP��$	���+��u�2��x�)�]��A���5E݀�x�W[�W�p���%�c+5�E3g��_�m�%kae}/9�����!�	�P0w�K?���4��y�E>�kݸ���]¦�����=+J�zxJ���<~�<�������VX$.Z~%V#�}��l#3�$ȥ���n(�$�n��������������y��"��Z�ߚ6y���	��񔣃O{	o�[��Mښ<"�,��`7+�$�a�wvŠq��t�9X��� r�`�z
��:|G93LO{$��U�Z�8�g�#�>�0z�s��*oR��o����c��	�T�o����Uɠ�~7��5X�ȥt:C�r�!�{��%��˻��6�z1#��[1I�)�)��
��q(V�V�s���XNcA�7[��$�vSN������N+!Kha1F4w��m�7�����`>��܌���_��߅��҃�he���N{�����R� ��<VVL��ۋ��ո�m�nq�C��9!�����}��>�L ���^+�Z..#�Ў��l�w/3�T���#5�(�����u-�̝TN��0Ó�]׸t��͒p��l���d�%��Wg�uP �0ը2����e�r��c�*Q7��':�-�����!�{0�(1�1ƴE֜J�����aT��B�v,�4����������vZ~#��T��F��T�V���ty^6����g�!��<�Ȁ3�|>��jf5o���(g�`����U���xF�ں��ye�)�)�DU��!�ҰS��*0O����(�QISg303����gQ;5z�U��} ��g��*oQ=,��"�o�jb5�N�B�摻'%ם�y�9���':�1��!���b,�m��x��e~��A�G�E�&���&�%�\�a�4�:Ǡ�&��� �M����\�22D���� �5��Ar�*c=^�7����$�oJ���y�v���m*-si��W��J�>`���ހ>zK���9��|A�;1]?:�vruF�(p����ƶ�W����jWE��{_���C}����0��Œ�����I��<������I�Y��\ʃ�J	ԗ�������O���P�ы�ϕP����iG��v�D����}e�dz5{)���N�о�^L����RVE,덄��?x,mnΈ�������]}���}!�����xHB�;�ӣW|�A9��M��`'�so疯5EG�9��}p�a��!ڬav�	�=��upqJk�UI	���"����Аi�6	�F�CW�~�6�zΚG�]w_�jP�鷮`޶���E�ZքX�ߩā`�6@���!�VbP`[�0�Kf��yG�ש����~.% E�ʃ.vA��$P�Ģ�&�p�̧�Kg�����苚�,�YyIu�S�B�o��}[�e��Iϗ�β�:
�"�n�tp�|Hb���(��Je�XQ#��OG÷?L�V4_oЦ��!Q���L�CpШ �[���X�a�L����Ǜ��]��t{��wp�!	��G�d?@d�K�yi6Nq���yF�4&A��oZ�>A�����N���*3QRǂX 	<l��z�R���@K�^���7�-�u�s{g�c��rV�خ�I�̰���S)=Q�V�Z$�����NJ+j*iN6C�z�9�����'���WJ8�L�:�A �*�A���J�����I%���2��?�q��a���<��zvB�	�3���$�F<�w~ ��Ѵ��19�?���%M�r����y��Q.|�w�8�i���[ٟc�lj����\��q8�&�I���amC�f	�����1�qz�N^a�w�_\NH�C�=.(=�U侂��G�17q�˴	�-���g*�=��y^^��^x�uh�xN)�d'i�@2�{�Z�1��!֟H�����<��&	�_-m���\�Y���~�`OglrK#R8�C���lަW���F��:�.Ww��J�L�M	|��c��'��ZGtQ�|*�f1c��ΞA�虙{�JB�,><�-\1���#�$ֱ�4/�9�;��lD��M³�@ ���B�G0�T��#�az`5d�N���[t�ƅq�|}��@}���o�AE����&�g���gs��@\>�/��$��!��Is�0
'F�H2�Ӕ L×��~��U�*����T�o�h�1�~=d���f����oo8���Lx���H��P�(�F���D����(�0�&���~9�Ԃ,�7)��l�`��m~����E��_�/٠��f��F���ySǠ6z��ߌ!D���]Ir��t*ת�5i�:��*,�:�h�E �ԓ�f�6�\�(X��2�ps3��%������hmC� }o;��e��24M��-��pr���mP��ҡ_�@����	Ę�F��;+yg�9��$~x<��歛Y�����-���+�|�iP�p�^����j&�6����(�R�墛�d�^a
ϛ��gS��%a���%+qi��㚥��
*��b�@o���zI��V��v�:�u\��	���J��ţ��\���� !��~���⧻��ۺ����he�{Nd��4C��i��ff�g���'��v��5Se��@y�cvk�~����/�-=�dpa2��˖�E_���
����<'`Q�&���FT�3<��&��Z]�%�&]��H	��H`&{qb?���c.���̃Pû�j����a##�!��L�5<��=��R�ǵ��D�n�(�Sb�]L`b���)yFn �*tsJ!T�'~������O�8|A�t�Xs���k��Z;�5��i=�-K���u5���%̮V�4�� ��Z�-C&e�?�l)��V�s���*��"t�*8�:섇�ȸAA0_��q�؊�"2E���/ڃ�bⲴ��,	]�[�FME�kY��aA�M�) @�
��V�p���'�7���]~/�͠�x���o���u�$���$���R;�]}������	ÔD��I�\K�R�]�Cf,}���O
��BzKm�<�TA�zᣡ�az��)�
��q��:v�Ӧҭ?�Q���ud8τ��ƞ�ʽG��q�f#�	��qJ?����qX.�e�^K��_��f�lX|:���i�ؾ"�j�!!�wz,�[YY�2
��߫��>�����,�ח�#��Sf�+\ܶՈmy]��|���Zi8$R�4��t� h<��;B���)5�71y�(]���ۤgZ2v"@rgx�^K���%u\dP�����p{0YSU|�gD��Ӫ��2UJ�w}gV� u;��V��b�e��@x�h���V�<8J��Q�P?*Iq��1|�2�;n���y_1�@@E��
�C���$�t�c=��L��+�Ԭ;nz��P����r����:�'>E#f�< 
x�g|�4�b�	"��[�[|�&������HDr�U Q�vv]hH�=oӳ�-�<���>{�b/��%]�4ڎ��'��h�!}���1P��X���u?&j6<f�/������Q6.'Ri�6����Bw^c���ʤL�K����*��M33���։�qԈh뒯e�$��Y���NB\��J�����w>ΤY���ّ/��eh����%�&��ah��pT�|�%n�ܲ���3�g�bO���kis���>��m� &L�\�x��y�*=�2���B�	Ds���5Nݤ�������@U��aF� ��7��"�n9�bd6�H���	�r��!V���l��=e6*�j+��J��)���H!4_�&_��%����L�^����L~g�s��v7��<�k�Q2]ɜ�pC����S²�
c��Q9:���٨��+1W\�JI�hM�2����((ك^4�
�<�>Z����a`:�DuPuZ.C��:p�<au�v�#GPz�:&�ɍCa𹜈�XP?DZrU	O�]���NfI�*�Qtyq����bS
��z�t�'P�.&;�����y� �e��7�EL����o�d%+�$�83��;����w�g�(�7��(9����;�^�X��.��e�0�������d�v�1E"Ly�Pѣ��W	�&9��h��-��^ܽs�u���tGO�����c���FGX
p�U�=��E���̿}O�7��d��>Q�9� ���6ԡ�vh��v���m�Mŏ��l�1�&��V�t���?JR�,�_��}W��x��͏�١�z���R�$�tڀ�X��i���@ h���!�.�y���kV������|��6ᕂ<A���h����uͷjc�'9]Z�U+<>|H?ʙ�@
z���ѣ�³.'��y�L(Aut�{��'���J1G����`�'��к�A���J���!��������W�:t���w�w�o[�|e�2fa
�����z��;�V{˩ތ�aW�*50���mA�޹�[���%Q�HX=�W�Y�R�۾-����R@yW�Xn��y=U�8�����(����ے>��K��v��ooV�G�;�ӸjM�&�u�rs$�~����؅^��zu�B�5���f�z U����o������W���#�7]��.�;�_��]2p6����l��*����L���$�8�O7�y�/���k��������UP�+ZH�����aW6 �x���Vz�X�9#E�M��Hp}��,H�̰n;��ٌ�,5�8��l�״�.��4M�u������ �r,&�bC�9-E��m�w�}_�$Xd5*Ʃ�\�P.L�:���P�D2��Ng\4^���y9, <���� �����)?u�FQd�ʁ�`r%��w�>�.
=�(��X=J�o��W��w�@yǋN��y�s��}l�}YT
^���Ns���Dy�J�p������B�;d� 8Ab�_��h�fn������"���8u�'P6�{�ZT ���:7ºi<��e�ϻԙS�FQ|e��)�|�Ԫ�d?E_y��o�`q.�T}�~�x�iq�4k�X?Ĝ���i���ً�*�-{����	k�?)����5��4@5E������P�?��U%�fN��T���.ض�����VO�o��"*�L�@C�)��48�9��>n8��1�\=��_����]W1�)�x���j�o��!ܹ��R��Z�QB��	���k�Rj�C�����G��5�����(L��C��M�o@Ch�$��U�Չ۸I�
��l.�d�g��<��r���emk<��X�*fpF�Z��z�9�!�-�l֟A�6�P�� O�r�+��KQ��!����+�=�� ��o����v!�U��c�t�|�M��Hǂx���\�4�qv��e�\-�|���hJ��-�N�D,�ˮ�}���刢	�����4�Å���ۏ����-S��} �M������_I�deA�pi_��c������q�Z�_�qq�
=�DZ��9i�}�2�x���"_�ɸ|��u���z���`�M��M�7᪁��R��K��i��������n�>zj?�����m��S�&�U�ֲbX��X���� �)S+"u;}\���Y���玧�$��Q4E%|1�v�U�ygQ��Y�p�ƮM���|�!�L��լnw]��1%�n�H�"o���YS�蝺��XݤWt6��]�0Z�)�,�hd;i4��o�Q��'���;{DkMQ�6��>z�:�0�q��ȳXs����>'�7�_���^AN��
�`[�!�6�4��Q�c�r
 �-��B���u��k�J�4^�bđY��٩6�O��T�;Y��G�$pˁ}���R�����M��H�ILi��C��P^�%��<�.5-d���ӧf��i|�#uN�ia|߻�
f�˪�����vс蔇�������z̞A���iټ��h�����Zg�&�\x?��m������0=é�ݟB� ��)瘀�5�~�@k�E���D4{�i5��w����i&z��咘l�]/�f�r����� NM�?�l*�������
��8��<�LO�,	R����������2�>:+����y�a��^M�i ����M�y�C(D9��߳���� ���s<iI��Ee�H�w-;Ӵ�?�D��o$����[3�u��ٕ���F���T�����LVy��b-͍�bU���W,�\�2w*�k�7�,�y�E���W�T}��e���I
F��rQV��|}នHE�X�Q͢:���N���9}�6x�Mb5�r�P�,����d��.`��_.u��s�Vu~��>�>�W�!&[dj���8&v�8���"~'m�ZO��J.���Q����ғ��k��o���������mE��B���&�_�^�i?���{/;h�̃��38�0����&E�*�LZ�Q00��W�1�;M�8�dҊ�tM9�  ���[Lơ��r�a��W��TJ��P��hb�+lrY\�(A��v���f���)U���tfI�~y�����?�xt\d�C���Z腏�������J����C�]�9�����A�ocT����gy���Y����6~ �K[gX�@�wfak��QAXFk>$�e�D���������Dٛ��F?��r�gs%�rW�ŤKy"�Y�ո������s01��ɘ�g�?;0(��p;/�����=�3鸚���Y��a^mj&���p�?b��2��Ǩ>A�i�Ȉ�-.�&�֯��^H�MU��,kJ�ϊ�糝�[KK#���z���鵀�6�Tv�H�z��~qr<���cm�jY�(�ξ=D��ҫ�7C��f����?�pQ\���.���;�2����N�B�Y�BΆ̳_�L����;u�E�9T#�-$��:���ā��Ɛ�Ed^'KA ;[�'��ӆh�Ŵ&��6�HĿ�Ӭ�@|c�C �IÔ:�c(�3�7����[:G%�
���U/�h��'�⧈�R70-����d��:^E�!T���@�,hU�x(�����~H  0��7�SBl��2k�z�r��Jej 9,V�i�f��xK�!0�ɋ�b?_7$?���i�=8��E�q��?�-Br��)� 5��Z�)N�A��H�Y[u�xd�}	sva�Z-����U�k-w�I2�o�u�l�R�m(ӫ6"2N?�9��:�A��T���b@hp$�y
JMW�fΈ�IGШ���� ��c�����n����d'�ǢpQ�xD�T�����?�X�uпof}D��L��Η��vY}������vZ���)�����D2F<w�n����#N�_�m.�q��U4�d��"j���3�3�"^�	��֦N��hs���_#+jwE��_�Q���GN�q�\
,�+V��4c$�0��~{!4V'�v�̭��8���$@b�Я)��ķцh=������-.( UE'�X�e����C~C�Si�Pn��˧r��1{@�[1&���;�S�c���R�l�'`lX���F�Mz�{��0�\���~�M�o޹�e��F�t"��K1�딢�!�.@��сf��!+~jR�%��ʁg�V/��k[�������;�wQ���}Xx·F0</8P����Xb�K��vzT]z�v�	�5�д+(�$�˃r��/l!Sݥ��W/���l]HӟH���gd��O�� ��s�}���	Vh0�]������<>��eӠ]mi/��W��n�2��>�!q���$�z���ln+��iܼ����΅�|y m��#�\g �ƃ�g�E+�LvV,����T=�ｪ�W�a����)��b�� F+!�����v�9m'R[�����!�\ޢ}��9���'��\�(�6�O`�G�S��B���cF�S�֌�TgFM�/UǇ�"k
%(���2�|�����-j�l�4q�$_�N����,�Z�U.�3ߜ?БT��u�d��X�6sMN�,�\;�@�x���!�Z�����ğ��'1Ȃj�O��.ڵʊ�V�0��F�K����ɭ*<��n��/�mľ�޹IѢo'^�90�L�Oky%�?�?F�5��^U�$%i�(,�U>r��bC�>jD���Q��Nx��`����ܨ~�Zzұ]��Y�/2�7n�k�ȭQ�q0�_1�,S7-Oh���p�Q�S���G� xZn�%,x#sF~ �P<#O.�k����l�n�|4_r�y����Y���&#��_��;��dnT��'���GZe�	���ѸX�9�O2TrM�gԜ@Ԥl	=ƃ�K��tJ� ��0�f*I�'x�:[��R�E�q&�+���g��JN;H����#����$���V���X:Bl�sf�(���)7�v;�ӻ?�Qh�yaJ�]��Ѿ��̈�$�&'�oe����?�X�Ij�ۥA:�1!|�Ǐ��J{�qi%~]��C��.�пd�as��^�B�#9�! .�R�5���U��ʉ��$��q)��<��}h.�>�|������	�Hغ�u=�q�Ξ
V�0E�#��Q��-`?�gޚknA#���/:�r�Tl�O��<�N`��2�؍u2�L�:�fÈ^����tBg�=�6)f(t׽C�(���<@jP�^W%ӽo�>��!2����8���"18�B	;+��N�B���f7y��� wU�*�*�s�߅���YeJ+�آ��iׇ߸�RX���^u�X�z'a��7�R����2v��3Uf7��!��	�A��Hyj�BnO#������K}�>�c�>�lA[���#��p&=�=�~�sT���B@B��Y~D4��w#�&l�3��{�JM��4�� $$�{Vs{��7K��!����0�-ǉ�L�iJ}�v��?�*gb�+o� O��%�I7M,�Q�\#a�����[ã�*���)NK4�3��c����2W��׏��l��9̊�) Ub����fb���w��n�eä��h�]]�اS���\����[	�����"o���S)(�^.i���S�	�dϨ�!+�)>ԙ�ݏb�iɴpJ9���kp���|�8p��{^ ��YgCQ�p:���G�O�2�jC]Y/z�@֣mn҆o�@C��ɐD��)23�P�@�����!�a,�Ϟ��֤�+���7�w4�'���7o�-D�&�y�r�ӌ��?�ԗ�;�yha��)���WD����)D�
��N����k�H-�;���z�<c8��Ңة�Fߋ����t�P�d �X}�I�%���S�!��%/�O�y���9p� `7濮�{��O�d"EY���Soy�M�0۽��CDA��H�Y��'�{@~��"���o�*�Oڡ��s�J69b\H߼4є�A����&#hv�n�?ǧE3�.���3{��˱�,�	��TM�'�vKC`"�
�E��aK�.J�o�d2m�F�� �$J�_Y�?D�C�4�Ꭳ��20�U�x��I%���5�8T�Fr{~���E<�|��T��3�$�;�0g�ViTXs����|�n Q�Lb�c,�a�ד#�{v�3 �S��p��ֿb|�8:���i׏��픬�_����ޮEQW�B���n~V����ٻ
p9>�� �,SK1�f�
���(ᄓY�+�&�F����\�Dk�5���AF�I�7�⥧�`nl�n����2֠���g�I��@F�@�*��0�C	���[XuC
k~����Ў�ȥp`�T	��`y%�ffMx��\婒\����9�����M��W�-MS�d�U�/dY/n�� ��³�`�BC��zdp�=Ě1`�%�i�|N�Z+���I7��{o����i��$(8?V�>C�	d_�-���t"tbgU^�<���ؕ�DKMwڬ��^�f��L��BD����9J���$��C��gSL9G2n���L8�u,a:�7u�'� Z/�K���w���� k~W鑳�M���N�%������˴��K&}��=�/����.�$�Hò���9�n83��.�JC=���zq�]m�Z-u��#n
�̿n8�mZ�#���dz���l'r�߅��x��x97�55{�^)�Z3@R�g~VFd�Ep��u�ݭ>��n����,�^[�D������i0Ы�n,m�.�Eb����G�D>u�ǃ����_�"K�����dǀ@�����ђ�+�ѴeY��z�S|�C��6:f[*RE��{�c]�����I]fC�{\
>���m��ZXF['{Y�,C��:˙�IiM�G4�f͠�Y0��W�d�H�j֬f�p���E���^��C���r��QЕ�N�R��ycJ�I�5�7�jK�{Ixr����A2��Z�E3�aݷw�d~���U;v�k��+W��RF�'���6!����ق��B��e��v�P��k�B��f�&��Y@{���kC;���������qN0NM�>�I�z�MC�4UL�|�e��F�����"u![�Ϙ��o��l][�@<��x:��^�������M-��m��И��-9�����	�-m�ݝ�N���+c��z{L���n�����7���Z[����W\c�z&�����7ԟv	d�ȫ��m��#���bO��io
����7"3��~v���[i�"�������V����oU��0rxڙ�dk<�H��X�O��ɿw{����."��p�v ��l��<��!�]�38�K�e�>��āyo]�Й~��o�u�����/�F�G��/<Y�S����
��M�o���$�6ٌ���[Zhz�@}j��I����6�G)��c��?���"w��i������.c̷8��;)�,(G��V���[����\���Y�p}�Ԅ�&���:�G4�|�Wi���"��E5r~�)����K-��Q�8fp���j���t������$?<M�S�dE��o�떝<5*BT��	z	k�)�av�Sݦ�N��`��0�����'�[5��3e��iu�6X��$�C|:��p�4p��EY��˱5�.*�6�U7�T��u=�>��;��c�'@y5�;K�s�o0;��z��*�G��7���z"u���\yx����m�6:�#ݹ�i�	��9z��A�`N�7�ﶲ� �F����J�Tk����3O�?�H��3��1>�x����Ww�;��t�Z��LA��bA����k8h!G_$�Mr�iw���ӌ�78��l����L3�}���y��6u��� ��u��e�d��_�c��],N�(6��N�v�FF,Ȧ�^t�ŭ57�1���Z��u2���Ŭӛ��q� b��1 ��<�ᬼ�5����Sg܋n$�^ίA�:����
�K�r}&��ɷ���2jL8��ّ���8,�;.���H<�'x�9�@O?'�-(��xQ*�0Գ��V�j\|Q����b{o+u^��;�����p�=8��C91��E���%\%�&�Y"vݓ��0"n��xJ�Ѳ��G! ����$�Q�}a�����BüQ�5�맖�{�~,��B�#;������O���@r5�iu��SQ�u��Ru� ���Kp�z�[aX-�K]dV���{C�uM� 5ȶZ?������xe�9���9�DN���H���o[`�W�[`I�M/��먦��Y���hܔol�Hy{���ﬞZp�B$^c��Z3�1����bxT�VsjA�w�OS���N�+F雕�������5�>���"��#d���<��GB�N=�}��gN.5�Znb�9��W���;��̀��s���b�D��@o�Tꉶ��T�Q�!cBx��awTτ	br@Mbe�W$WN�&f(�-�0J�5�x@�r�(eo{�%�|
O#���E��	��{7��GB����������af��qtsv:���Y�O���@\�0�#��-��N�]�g�c��'|Ģ�;�r~3�@	A��W�d0_+E`HW�� e�O�D���z4�L^b��F%S{v�G���oL:"���W�[U%l�{ѫ��/p�@��V~!a/r�=�d�#���Ov�:~�L0&P���ݤ��lxArD0����NTLU��a��o�7�����v��������ɐ�u��A%YsH�6{�b>C�hS��x��]��^��5����D%��I�e
G��[�yߘؼ�����`��J(�)�@tdfĖ�K%]{w3}�n�4X�\]�: ���7�7���9Bq���VHc�@3O2|� �`�?�#�Un���m��m�	j}j���'F��pWz��(������y�jf����E_A;~73T�NE>' ��ROH��I;��c�S��׍�������s��&_��d�C:h�-䂿�����}n	�s"�sޖ}�7�����eݾ�GA�R��H��u��B�[x	oyyr�����f�?[�}�-�y#e�����}Gs�jl)�T>_�Hi�"��>��C����f���\}���v@�H��<��*��a7�,�h��Jt0�&Fa����?�����0=x(��mީ������{Yhc�]������Ǡ�.bC��P�d������2�GhF�����;��ϑ9)��<�����3풢�w��sɵ�C>��4?��v��N��=���էPI!��c�"�q�z�	:��	?���2�S����cN?�٠����
�P�T���~OR�NY/JЇ "�f�%A�i�;3}��e��3�Z�ɗ��h�qǿ����ȀPU�Z�b�a�����h��ʷϞuD�>�y���������[P˱��C���&=��يP��h��k9E˵R ���V�=' ���?��1V�[G�z&�R��1=FJ1�n\�*�wݕ��B��|�
�3�p|Q<5`Ƈ�)Q��o��#�`$\O�OU4��9���K����Hd�%��5g@�_��6���q	�SI���bl%g�m��h��An�Z���uⷒp�n�LH��yp�ƫ�n���wq4��6H��:F�~�:%\62��nL۩t�2�����uI��$���@T��J4雌p��;X��b����)�X�棻b��[6��Z__߳s}�i�u�	O���u�� crq���W.���|c��*���ָ{T�� /8S�+�9�F���f��N:�pAb)c����	�|~ܠ��gt��D�ߋ�n�[�~�h�('b׺�Z<9uOo㴻ى�c�r�M�3M��� �$��zi[�w�؝6��8�%�/v�ȩD�1���N-,7�6���~�����
&OրJU	(�}FA�8��8qۮ���S��Ӻ	�� ŧ��L΅��N�;�9i��(�3�M��t�N,?J��I�y���!qIaq��N7����u�#���?8y�����d�k'I�!��Pw�y��/�9�"fm�d_���/���聑a3�[�lX�쨵�B�r��
Z4�vZ_���C��upM�Cj����첚�2��������p=WMW?Ge|3��H*����+��7~��m�&C��{�6#{�iab�8Wq���	>�X��V4����ϔ6I^�Y-��!@U�ᔏ�$CRO��5�t�.l�!?3�k�u��N�??$X���]'DBlz����9�[�}�-�N�Q�,�vA���0A�n�Ɇ�-m������f���FJe������6e��K��J��z�����HV+ר;�K ����w�ڢ�ÈSj�kG�7�α��E����Ǝ1^Ŀ����}��k�B��p�� ��������H$��=B����P7.��J�B!�L���[?8i6@;�_�$��{�N�Q�+���TXz�:���Y�W0aܽ����H�����K�!s����چf
�P��'����� �f˥�><��A7m{#�&\,/�}����)\��SQ�NN���sА��]g/�G`�9�ll�pT^��������g��>'��z����jR�0<��G� ��;���?�?�Ҕ�"�Y�b,����?F
G�$�_ˡS ���<�\���� 3�P��0K]RI���7N��!ߩ��#���n���m�ŌY�EV%�߲�x��8����C%�b��]��|�����Ԋ�Q(7옐���Q���١���_�6��& "H����ׇ���9�Wqu�T�D��(�೼�R��=uk�e�0�e�P�C��gn
�E�������nc����T���t��~*������*�?!�0{E��-B����'E�v�B��W�T5`�o�7��b�~�Ec�����������&:��B�x3����C:N�8I�p����P+Iɟ Omy�)�ke�#P'/�����p�R�H�̀f��d*P�8i�,�s���gM�2�t��DĲ[� t=�-�[�'��~G�S�8M��]a�앾k�d��O�<��F�XyG�H�f�/�>>=*bv�^�x"oDW+��<I�LЬGt�����JF�*�b��ǳ�����fa5z�Y5��ʎep��^�z�	@�:�N�
s�F���q���B�rpB���E >m�Iy����-:��K�?1v�}h���i��mU(�1�XM�,�V���Ԙ�s�[���1[��V�i0��m��[Yф����n)C�yL�&�+IK���W���\?1��uʒ4��l��+QzcT�j7������!���~�E]�����~�j8�()�n�a�XB�a��c�nh���s0n�D'�>j'�h�x���"{e"�5ۺ�2���g0rb�q,5-��# �v���\ϱ,2�׬)��Υ����{bn��찝�0,��G������yQ����%�%Վ'�����:���0�AB&��=�����Ǉ�+�x���jԆҕ�YQ�0�������dZ bqܲ����b��YC5�8f��sS���C;V�&UO:��ÄIj�.�Qs��]�$�9ްX��zs�k������.D��Y��"��*
��[��SC7#����n�B�we$�&W]��_`E�7��~�_*���z �ۜ�����}����i��IF\�����G�� �b��(!{K�Zڇ��g2Hd_��"R&X�R��)�^i����'/l%9���b�l������_�́sO� �VƇ�[�;�:�p`F9��?��QiR�ͪR[�K`�'#��V��CN�Cnd��_�%�4qG��֙��lĪn�\K�Q�}�.�CS���`/sJ~��m2V��[Mo�0��N;ʡ����u��O�D�+�`�f�<~�c����(��K��p�	���ME�;p��N{F��܋c��8����k�>�Q}���Ǖ���q��w�/
�@k�X��6�3	W;�A�\o�ci�����(f�j��diɠH�W�(� ��G3��}rH���O�hQm��g`�1���	8��6 ����}h"��4/lW���8t
�@e�M ��^��bЂ��B����}(oY�n'Z��l��L3E�
#'�Q�pP�׬3�j+�v�Y�$��\bߔzm]7�;T������R��F���M�.X=Nj��K��wD�����j
�,�'��]q�d{^�]mG�,�ȃ#�H��[��I�]��=}`ⰅH���h���gc��3L�p�W��m�=�\+óצ3M �A��x����r��a��a�%Mf����8c.���Pe���P}��_��,4a����"�"�F�N�z[��r�E �!�3֢_���hz�n�4UP�	�DD�#�|���0fx���h��g�^Ą�(�7����-�^�$�'̖S1$���w)����FF���;/UMtF9����~SO^����n���S�eZ7f�[�$�pk�_x��G�kŌ�S;^�n8pI��
l;&]E�3�<I[�E��F6� $�T��dѨW]�7_dB�É��jT�X�5s�E����Qؗ�ULB��s�s�!=&����X���4�=��M&�.�UG^%��Z?d)5)[�+�����+�hl����r�� N��"�åy�id��Z��~B\�<q0G�g��|��1��˃�6:3.�;��i㼀	���>��a֣��V�6����;y;i*9�ɖŅ \�G�iL�*�Qm �f��v6�l�X��� ��嫽�<�]?I�4Q���z��s�YTDm�LK����_=gJ+��[�]˯s�Ƀ��1sUf��4��FY S�E�a؝i�	�߲I�:���ft��� �/pi5UF텶�Y�\��Z*%��D9KT♘����{4㸮��n<e��Y
M`m��Q������Y�g�v���i�����ʚ�	�-|O���@f��#�'��\b���_�9�v�`�a����|,Ǯ�X��q�m�!����Q���&�Z�
�����aE�)#��ϰ!�"����q��AHyr'f���5�8sH������rK�%-!y��
P��{���;?����֛wX���.�ry����g�??*6 �$��|�e{5����^"�ZE������ܼ���B��ڐ�p�������)=S�j#9W��!,	Lx��C��C�m�����	I�#�Q�6)Ibz���,�r�4��c��j�wh�pp3��KSqU �]j��E�7BI�^˩��,���!LX��+��)LI�u3��4Хr~��߂�9rMh�P���ǏT����oT�.Ӕ�m�F��qG1ۨ�[WҞ�U��Fﺂe�z��9c���]�*k��j����5^'bY=<�O���HT�(�Y	#�{iv�M��]2O_��j��7�&��QB�&�$s�����9A���x錀�$ϭ�Z��G�ҥS�n3�8%�{�[SoЦ��Qb7���T�̯W%��ڂ���|�.�>� �h�J͂����09�=��4�-�߭�K��M��J{�����j;����6G����*7�h�.���n�+Iw.%�n5ş�5���<{�op�A�;�}�j�Ca��)�m�rG��zvxw�Y���;�@>��'=�\ϻ��0Û6i~��=tH�	k|�I�����dۘy��G��dS�i҆)��6
?�;_�)�H����*+��$��A�)�U�Ϊ�[���;pS���wu�X���5��c��`��^+p�
�o�9n��W����lzܽ���ߪY7��-��+���{��ǆ���� |����;�U*��,l���Q��ހ���W��cl�o&d���@�h�C$��E]��U����I~�qs5C2�z�)����k�}US	��h��jb�.d˖��6��@N9�k�~�^��%0�[j�(*2�~u�^��w����C�τf�P}��YXh(A�",���z8zx�E�4`p�z-�`Ա��VəGZ�"�7�����,��rh	�zcͤ��ģ����+'�K����0�乎�(�����&�Q�>����ڟ�+/�sZ@�y���4O��	��%@S�8��ӱ:������t�蓬�,�3�_#�e+��ި�#�|� o�٪a3I�=5I��Lؾ�_�x�)�4����(�U@�H�P��]f�t��Q�>���у�x��r^����Xh	SO�0��49;�`=��K�~ij?V���'%_%dH���cǎ�pt�i��A�ݑ�+� O���Tqy<sB	��AN�/|���k�!C c}�&D㦈�2�=�yev%@�N��,��3֍:���mQX`9�y�Ι����{_������H+�;c�ǒ����ߪQ3u�܉�z�˧qO�#�����6.(/K��_��Φu�+�"�S�s��O�ȟ�OR4Ȕ�7��IC;��9"j ��}����4rz�Y���%�I�K��Y�ܭ����O�:'�/��b��b�9�dp?���$����I�SjK����Sf]Q'�T�Y���{ͺ	�\�t�b���S躻2�~�v��8��9��n`:�8������}������R�xX���R��F�Y��WL_�w���qqe����5�$`*�[-0eu��������a����1J&�%_�ޡ�S��M�Y��t�4���d��lfFsĭU����)���  �CT�=���=��`0k.������9�\}�1\K��Aѱ��]�>]I�) pI��v�Q����2�d�.��
ϳ�,R��ˋ,1`�q�8JV�<5���PT �>����'�o'�`ֲ�E���-��0j; !+�j%*�K�d�������Y�S�����н�w���N%6��I��Bz��r�3�U�>��F�8�a`�3p���Hr; ��bij����D��*��P��I@q��(U��ߦ�
���=ĝ�Zڌи
��O5�K�mFL��o+���A��%�~��B���᝚I��{R6�������ӛ�,&C=k�FHx ��p*���B"Ӣ��7���n�HO x�0Y�ܭI�ʀ��9���硛akKex� ����}����F:^��8�ǂhb".���˫�y���N��S��]�S�8�Q ���&��'x�|��?Ԋ��$V�P]+=�����*���r[�}t��w^o|�%�92.Y�:n!��č� 5����:Gox�������a�/���>��Fɒ�D�(s��䰋N�G��۰t�Z���U���$=���q-�6��q��0���
�����Ԩ�R޿ժ���M��,DC�`��Mq<ԣ���:���ҽbe���~G_��o&1$[26L�%�p��@A[ٱqk���^�G���z��ڈy�٨&��|�&�K�&��uހ���7����q
�m�o���b�:�i�z�0�J�}F�qE���Z�D�*PD�� �8�R#A)���'���B�匣z�y���d>E��,���C͌j���ʶ�=�X����TQ�nP�P�����p{�,��0=wa�b�Ԟť$�~��t%n�e����0��
�p[kW�`d+8���	������D��x��V�w������� ���H7��8U��g���������L�^��X�8F��.~4�mK�a���Ѝ)��Z��z���v[�����o����iȭ�,)�Q:��no����\sQ!zEk�����m������)�gsIoa'�syx��p?���n��`�(�ِ-���2�a� ������9���>�W�8���ڗ�M������F����o���l�ڴ�R��}�X����G���Ubk�BC��KH-�:#�� �;��I�z���UF�EfT(�(p���6 �7�ި��s��Iq6������ֽ�]|L
�j\G�Wٕ$�F<��n��[f��y=tף"�C�6�	�m��.�oc4ڍ5������"̫��\NL�:�w����bo�c���R-	��["�����#M���<�u@�m�y�&l�F����Э7Rb��8���T3s�q�s���`j8T·.-nA���C{ɒٰHN�mA�U�>���Tu/��O���F$�Q�G(�Uv&㩅#���G҃�Y�< rx6�{��|lC��!�)Z�y�2o=��=�7LpB�PP����
��H�k13�����$��֊�D`�Y��I5�b��+�nC��x&����8E��a��)��5�ȺC�%:��9���u��P���ѫ=��sZ��㎘oM�2e��\v�}�O���'�E�Tů���t3xk��7 �ȶ�0f+��csQ���XIe"7����U77H���{��Om��Ԑ��h#���ڝ�`��[-|7݄󮰬�(QY=��֙ ��3���^�J��:����~߈�n\�&h��5�U�P&�_,�9ժ@
S�������&����c��a������/��9Z_�%�l.Gjk3�u� ���t������B?��ی��,j����r����U[���SԳ��Ž=��F}?|�(p��;�b����]*|�T��������T=Q�?��C���r3�gR|l 1�_�y�0�%��5���`���G��H�PH^.9xDpߊ�G6V;�4u�h{J�dN���1C����DH<{�*tb�_�M$D.�=�65a{�d?
MXӷ-1	m�§��ʯJS�΂��������6�_j��/SY,������ڛ���&��W�23M'���R�S����؄�U��dB�KF�X"<ȟɒj��\��}c�*TC� �gIU4ۤG�$��~9b�g5M�^�Fr��x��0{N� �g?զ��]�!X:*��D�����mI���"*�焛#���p�9����-�8XUH�|�G�]�h�!.N�]q��f�6�R�ؾC�!
���{����فz�4
hHpaٽ��Jm%��^�G�H0�+�X5�����G����'�Db�	a��赸-Ͼ��X��r�����#��T������󍟯��[�^vt�Ƨ�$_6���N�#�~�7[���a��ңD3s.kPR������7�>��,�}��8iv\��^�ヹ���Q�6��^���I$,B��(ZRO�|qB�~�3�ʒ�_�Aj+dK��$Y{o\X~`�7���|�ٓ�3��
�=�[��+�gJ![���x�%��k���&OX�FH� ��:��2d�I�=Z��P����:��0-Y����y��{0���ޓ���3ݵ?��1D�xY�)ҍ���R���3���1���-D&�{n-}a�|coq�A��َ�Hy�Rvf�ZѥN�1�|�ɯ�B���� ��I��wk�Ons����}���n)�?�$^%GۧWY��Y��^�[r��]��Zi���ɡi��y"R�I-'>�
J[M��F�õ6����s��d�,��sh꛰�{TC�_`��K'�(s�ОJ49���<�_�����	��w�.�9���-�7M�Pf�y�,����zr�Q����?XjuP�w�%M��S�3�4!�Xx�������a�Y�3f�llq���R,�1	�=������?y*��*ʥF"�`X����)�hZc�=���	x��Q�&K����Ɨ��"X�{jKO͒J��zmg���pJ�2���V�ԸD���=��H/��"~�X�j�	�X	+|��%7�Y���T�t�
a4�~å��=�/ﻮ��tJ�'��Ph�U*//�!��o�#es�ӳ#�GF���톨P�_� ��:@Мs�C��	��=�[`��9�Y����������Ahe�O��\�Ktk�߿L�����o4�¦�����=� m��eP�W�[�	�r�	.�B�=��@�e_Y}��x�Ks��Wz�v\�0,Ƶ@���A+]���)�T~���x����Wl�Ճ@Mkډ�J��Ҽ��O�d[-��� ��	�dnG��0a[0�=`�.)��b�7,�y"��PA��V�{�ą���P�S���&���<I������/��j�ݸ�ڂf(�:���e��6�L��0��y�h^���'��A��섽o�w:+�F����x2z���JSf��,\,�F���&+������?���$T �Հ�[��xo�.��:�M���М���6�S�9p6v��*�6���f�bIMe��0�CKښ��G-L�oS�t�2�0m=T+}%����H���éDK�ʽjj(��+�U����iaɊOk;��o/�������O6�)��!��?���ЀB�ܦ�&�>̟��T�T��'�g0�nw[����\O{#�-1L��9�L�����c�E3�l�i~�VC'�#[g���G�1w;��?�u(wT[��w@ATW�F#*O>�֨A�u���g��4)���YF�������>'�Pt��]���� !ܼNN\XIB�tx���m�%.s�m$��������3w��j7,�g��$DN�b-�.�{D�3��0&� �E6q�T�r��ՓY��qp�Y�ھr2������m��y�^��udӿ3��u�`�D6ݤV�U/����� ���f2���ȴ/�~�_B�YE
�>w�T��5Ҽ���dj }�\�F�*��Q;�aJ�FS;������U?CZm�%ՠ��-;�)��\�8b,�V1��ã�U�j�Ĉ�!�.�����N�	��R�.�E�
S���*�4�^j�]�ʕ�8��:�F�t�����
ʌ72�����YʵW�./�H�2���הz�:�u?�q�,�D~�Ġc���yk�%1��#�)���lt��_]YDc����s��O�g�c)*t4#��$W�}��gN&���k�tܔ>8�0�E�bx��"+�Ȅ|,`w�n�4�2:�O�a�ʹK�2�j��	"�R3�j��4��q��$���x7'�Z~��^��!�WE��A�.]������~"�kNKX��Ι�
�xPa�<ÓA�F����I�]�A/���c�U��Yݠow�磃H��j��c��L-s=���CG��	��:9��
�"����mdw�CU���݀^1��ʍf?ē)@7<��6��Zqa���{K��(���m�L񝩫���w���"�ڃ�Ũ�+�|{����]��S��Nt�N	�����x�1c�Bsj�Ƚp!���� 4�4� E3��n\4@w � �N3Wk;]��j�%��e�]@4S���?<\a|>h��1��F_����%�DvHbEy��@f|ًl�=H�L�H��M�+V��Zz	�S.:�]���惉���
^R���L�O�W�'Ŀ�X�ʎ��rD(��'9��`�N�%�bZo��<���S�3�z�Q�֨R)��?c�6ġJ������,�x~D��$�F����[��i����-�^g��TD!Yb��ó�fd�btk���xU�M��J�_j��9�"�*_/q�?�MnB�`,s1{�o��j�U�k/�l�P�|+�d���GY�	��]���I�m,��^R���:���J#_�L����}hK�J���ൂ� ��ҫ��iq��Hc��2�S���׋Cq!j
�;�'�Q絵o�L90h�'���SN��(�(>�86�ѝ�����}����i-�?<��+�"6��y��;g�y&�{��6�^���N�I>�D�Q�]���&9�
n��Hu����-~B�Z/pْ�x#c�3�r<?��os�Q�
��3�?�[�r�.�����F�^���*����ZKO�D�b��l➐b�K-�7���������JͦDy�,W��$��B�7��w^\F�?��>��Y"���ȬB���B�:W�X���?iM�^��3\�'�@�M[�cD�2چ���V�.���17']�s����ڨ�tI���:^�s�{��6�bH+4>)Ə@�	�gj"�����ة���f3!m�YZ���y��bA����s0+V�B�I�AA�m�ѷ�4��YAF]���?�c�v�"(u�c���	H��tD�o=���%��VH���&�+���I�=��ŮSu_9Op�mǰ�M;��8#�3=�~~���#��f�XZ�|O'Ԛ�d��qY�o�lg�B�(	��F��n��6��	�D-����H Rszq

@#`��4h.)���E/�>���;��E�>�)�t)J@����R�Â;ְE,>y�$6�|���(6�Ϝ�����d�&��)q�G�M��eIJG����i^"=w��)��&Z��y��q� ��7���~>����>��mE�J���Y1�Mŧ�V*����1�h4YH_���w�s"����&{b��f���=쒾/��i����Pt����V���&ȴ4���]� �-HH��k��ۗ^"k�uP�9����CS����?����|w�
�jT[�ew����)�	��{��p����%�z$��K��f"￳ %Y�6�4Q���jY���4��-1ߢߨu�ME�H�f��4d�l�jֿ��#�l�OCx��_��;>c~
��-03�E���L+El���U��}.\�\�Hk�Z`+��L�rc�E�hc	���P���En,��x�<Ү�F�z��L�q���B�*��þU��iO7C���;��G�Y����k�啢�焯�JG:�`�y�pV��f�Nlx6L��u�f���_��9���a�~.Sר����"��}�D����v��C��A%f���a����@ӺSQ�9�&�.�!-�v	�ܐE��bILޫR�������|f[��]�����R��6L1@ws|u	"��A�P�tebO����?(p���O�c�!�v��\I���~`�1$��P�-�.iG�8.�|3F�ȟr�� ���ӄ2�,�l3JX�^T��L���ο�&�������*xN����R뭙#�l�H�y��L�6�ؑIU�8�/s���	}��m���@0$��QY7@d���dG�g�:��y��}Pm��֙�S�I���X�]Ƿ[BN#6@�A�K �q�[�R7���
��U�x�35y� I*�mXm�d+g���R1��gÒ�j�45_c|R�E�mĲm!r�;s	�����g��U��s���5�/<v�4/�Jvb�ώ(ap2�o}]I���ӶM�
�x���?�1+o[�Ď���T^�� Y�H����H�Ȝ��w��W�� ���1��t�K��E)Ab.=[�<E�lH� ��������S���^���7���Yu��ك���.�`��yӏ����[զ1@i�c��͹�Kg2��� �O�*)�|�q���]�b�2+kZ��c�|��N�� ��_5��V��4�B�Kt��«SZ�"�k"aK�:�;QB�vr�Ѧ���\BeZ���v�����'>�Y6[>M��;�U���l�� -h�\�,�_�F�0v����j�s��%'Ϲ'��5P^��),4Ɇ�)�2qZQ�%�=ыq�2��ٟ���CE� �$X_�29����jod�y���-:û�$�P�`ٯ��V��K�c=b�V�ā١��^>C��*����5�x$4���#g�2�v\��,6�V��'�%O֢/3-��j���������T�m<�����צ�:X-y>{��\&��#� l;:S�9�{�
�=Ig��4 �a3�� ՖK�u;�gr��{r�Sn�MW���T�T̻.�!?b�F�խ��'�K=8��7��'G[W�S`� �#����B@���kdbr����_�U�KyKw+�Y��8�c*52�4r\��LD�{1&'[���q��e���-ayVC��얖x˥f�̪�b�Z�^a��<̊ U�'z� A�T��$oA�?�3����G{ϵ|�l�.�EኡP� V�i1��K��.Q� A��0��_�dB�nv��d*���c��QX~ʏ9��)4X�F��+9X�Z&��)�������i��:���I���)��aZ-�c�ߚ�}L�
����0n����m�mC(�����C���~�xt��N�JBlW���t !�=q��p� �Qo���r&H��\�����1��ұܘ��|kV3eY�B{�-��a�7�4k?�b��k[,7j,�������u7���oE0=j�������{�.)v,�''���92�L���ԕ���m��[ʨ�էl"��� ����49Ujeʦ`J�P+~����)�c���1;�k��E�hesQ�"� �|)$�D��'�#Z��}X���-�~ޑ5�ـ-�k�]Ī��EǏ��.%*�U̾@��D#����h�����T֧N�]h6��B� c�����CR��L9G	,��8�z̻7�o�� jV����	 g��e�Pߞ6�B�2�jR��S\�,� �b�'�jc��ݞ�˗�w�.�#�X�v�]bt� /�,)./���a�<}I��)\	�_q�=!�����[�)����-�.�
��L���(�R�X%�nZ�j9eQ�M	ǽC��
׮O�i�We�Z����c!�ڕ���8�b(�'���g��]`���L�gwN�!#߻�`��~�#]�'hz
�6����Ѵ�;;���F���cK��箣��	M�#r>;���|׏��B�W��o_k�~j	��`O�D��)��)qC�`���J�8��1#�WR��KMS�̹���Mn�Ӡ�1�j�����f��)`2��4�Ѩ���o��S�
�S���.���K���U��Pq�v3:��	A�;A2FH�3�{� �U��<K�;�o ��^�D��,L��gU%�se�͓�����D��׋��&/6�Z�Q�?E��eX="δR!ީ�$��wYF\��{6����j��Lu	�8Ft��	#�;}.�&肄@�9�V�bQJ'�TK��-�ӷ#3oq.0þky�� ���{>[Z��&q�Yl��.�$�j��6� ����b�u���cR�)��h�Ma��%�8_�!A<l/���1���4F��Y���W�j�#�]w*
�2R�-�����I���EG�2�&��J��T�G�.���-�F�B�]X�xP.19B|{Ӥ4��T���v�����t./���A8z�
~���<+����nB��Hō��-��c�(���C�N3q���l��d�_�a����>����Pi�dr�2��hX�WUƲS�{y!v�2S��ղ�ٺ]�X�G1���NI0�ǰbg�n������#�}��AUv� {T�n/��ۂB�`�X~b�Z�|-�f۫?Jg����w�zƠ'�������Zc�U�R���!�"t;����2R?i?[���R�˘м�>�R��)șh������=�F���F�~B.�4��y0��ݰ����o(a�U8 q>yh�5�����-3����bNx��ʎ�/rN�]�v�ǟpS�w_~�`���"�N%w0�	���b�/�6���1�1'� @%\pp�$^V�S��S�A��] ���Xx�g~����3��)�+�A��崚��o���$1Ҵ�ʭq��p!vj�y���/�>x�؃��ݸ�SN���R���9~ʫ�f;�\HtU����8����E�.�o;?憮�(�`Ө >IX3��
�*P�R�z-��yL$@�T�Y����d��oXȗ���~�m��i��~-�,�59M֔߼�\
�-1q�s({� !D2�݄ �5�2����ldu�i~n�2Ċ�ۨ��c��,2}��$sއ���j����W�p���B�?������\�V�ۥU�[{Š�Ps��6z�n�<��qU�._.�"ꀙ�`@K! @*$:~���F���5j�
�-��(�:k�'G�n#��9_��/q�~9"3�eן9"�z �{��>v�u6��,ǅnz=MzM`騳5S���4���W����A��cR�c�~DQ����)�@O`�c�ḱ�?�� �7�`,J����t��` ���|ro�y�fI�P�NK�Hd�9��3�K�� �cF���`r9Ij���4u��'^B�1T�"﹖G�$�p���4���2��ݺ/�`.�NO��K�J�6��gZ[D�	T,SmJ+�9��x~��|�|����m�`Jc�O�KdO��Ͼ2�D�J{���媉���?qv.B�ܱ�d)X���`��� ��8�#�����n%~�@l�g��+�)v�𾹨����������Xw>	�BSXɭ�|��o���>n$r�X������@[� ���L5\�QJ���~@t�/T��3���q���j���)�t�R$K(��5���L�vP���Ͽ��ɞ���ReM`�ӟë�c� �Y�LE�w�ESO둦��*)G�j�s�ŵ�D�`����fw5�����i�b�o?��0�����w�R�!�	�^�s�y���H�`Ф�o���^����>ɖ��^���LK��N�1���L�e\(Tu����;�������d:n�r ���b�r0��9t�^��sPHڰ����8��1���M�\(��4�9�2//����3d:�#|9_L�܌:\Uq�n<Cn',�|��l��[t@wǖE�{���(��1�B2�P'>�����97����|�@�_��:��K����;1�U�lPF>^`��1cukn��C�XW9���R�����KG��������#u�;V�]`>�1	ȜJ�Ak���>�$��pӚh�/�V��̔�����r���m	�zr� �Σ!6GB�{4�t���y~~iCn��5u^e�G=�t�1�I�/�h��/��n�-��r��@se���rO���A��&����XW,�b�:�UQO�U�$:��mj̺�_٥x�	���2j���Z7\ߚҘ���N����y��zӖ�i��o��C�+W�����X6��4mZ~`���fq����OE�n�)ey�̰��9 ���U�>ܙ?A��f��u/`{��d-,��s���:�*��k5�1�2q�H$Z���{\گF��f�Ǎgʞ,/{}r�^}tA|*�Dr���W�ݸ�.���.��P��F��'�ӗgo�j|6�Z7���
m��IU��5l,?(|q�	|�����YǛ����Ãa��Px��HT2��rVC�=+��77��RS+4�f�aЩk���d�@�*"�?�3^��Tj�#��JeqF��������j��I�aՏ�XZ?��,��&B� [��0`��S���3���.I{���}�~����^�,�L��C�d7���/�ו�sV��&��-x@�#1�;�C��+��6�n���&�g�W'J4����P=g.�4l��F�OV�
��:�����G(:jNug�F0��+�|�4r��?!�E�(.?s�v6�=J輳<�.���	n��Oӑwd�D�{��[[��zZ7\��@��|<D��k���ӷ�� ��ļ�|�Y#��lތ�C�|	���- !��UpB�T#%x�H֟�0�p��(�m��	���f=ep��%� ��o�kh���7̻/7zR_ğr`���R8����C	���y�䲫�S%F� �|��XjP�ykUN�M�j��W�M+ǊNtB����-�q0�=ԩ�;7��z�"�]���F�ґ�����J�p�R�I�)3��@pC;��Wͥ�Këqоf��W�p�i-5ğT���{��l������I��L����q3�-�!��`<�w�����k��Sm�C �_F)�5��z�����6�7C�W�l�g�a$��/�\O��zxTY��7�nHdL�蓚G/�/s��d�ӕ�h�����I̥����Gɘ�1@���޺|��^q��J�ԓ֬�'i����d�����mCƮȂ���[mD#��RyU�d�K/n�s�ہf�H����Ah
B2Y�=���4bU�C�-l7<�$�B:����_3����!<Y�����o8�� m� kem� NJ���������A|�AN@Y�p���Yf�t8i�0�]�&(��f�WwT���D�޿Xci�ʑ';��T��`��J��I�6AnB�DE�� l�Э�o�v������آ[�Z�����0�A)�2/�$�J����Sk��k�yL�7>BIw���	�0��h�c�`N��!���F�n_5�va2ҹ��H��z|d+�ܑ�L�?�/�]O��9M?���k�>�Y� �P�`%= �2��W�K`�8BK��H�H�|��۠@�kT�o��[-G9��q�2�FB	^���䀯��-�ك�Y@R��4��O�e`->��n�>"\9�|�BI2�>A��ے��	�еa���Ff�9G��I��'���L���i�$�����ɀA��x�Q��ȼ�yH�$);�T2߳e+e<>@���hG�5��#a5�	��7Yӛ"�鰭��؅J�8X��/	����
�wi�	Cö�yc_�s>2�������v7��8�F0^{Ja�F�
�v�6:\չ����*�%1�H�XYL���+��J�t�r[,:I)���8z��Ğ�{զ��������9X��I;x��>�6S�?mmwZ7*�bI��1��	�L2|��>�|(�ݼ�z�*D��MT�ׅ���5]�7ĵ������ �Īґ����d5W���x�����k���g�����o��
�e�-`�;�L��⧼���fWTb���^���������v��S��`����[,�{��xn���,�"Mm�%�ᆅ�4����@�_m�0�x���L�ܙq4O��x�a0t���������P���u �t_��]=fPu��`,��}ڔ��#�G������	�e9@)��1;s�g�gv{_��(��L��u�S	�p����~�OZ]�5_Y{���^J�+HTt����;RQHBJ�h�a!���Lz���8�y��&�(�n��n���̮�+�\<���2�!�|��
-9j��qx�|���]�*?�䋶a�!����CP�z�W�WK��ݶ�6 �E w�)rju��������,���ź
e��Bֈ�����5`��w�Vyah.�R�Y�o��*/�����yJ�]��2���fZYAĵ�o���Lʓ�xb�t0O���'��g��X�u62.2�y_��Z�LEd*>�J �M[U��������ߙc�b+­ \�W
�/qq�>�?S���Mz�=5�XG�>U�g�����y%�j���D�B�x������b��R_X�Ւ�U�17���\I ڮ���rC橥kX��l�6O�$�c	}����F���K�����\\ᆠ^�6�i��Zז�Ϝ��~!��4l9�X��-��B�^`;���>�:���e�0�oW�. ������Ȗd�0����A��3��گ�-S��4��M��}��!�P��m�{�ʁ7���(�̀ȼi�@AyO=��J�W��L�L��Imj�[y��g#���-�)��u���n8�e��-��c�=$�6�0�1���n���IL����GB2JݟG`��a��Y�I��Ժ�����G��?!�7�8�<a�� B$�A�67�:f���.C��e��Є�<���_o?�pߛ4�d�ezBb$Ķ�Q]~��sή�73]5
*g/�;�#_`��zq�۸�ߞ����6;&\ӡ�M{Z�#ΣV�h4@B|��r!������cK��"o�P���`��N~(�#&�n�x؃�O�K}ϐ�/����Sj�RQn��N�v���/x*����k�=��S[�1O�C�Go5��C(T��������LV+���Q�	���xBK鰬�Z^�Z��z�
)���=��L�D\�5ҠnZ���ijsdY�h�@m/f�2ka�6k��~�f�$n��P&�r]٬�����1�\��T��h��_!͉E�^Ab�P�_5��2hâЅW��vM���w#�	=�a�Zm p޷@��a��o9��` �Az�>?����6`{��@�O�h_��ۊ�=���	��S���4Y�f���I'�=3u�wU9G��{KQE�%�$�>M�`C����-U�����XR�cB)�^���p��6�r��z�,!z ݊��F1�����+�S��Ũ���+C0���G{B���z��g�@���8�a.Ō��m�����Xڲ�h���`���������e*b<��%��B-�9�*��[d�:��C�L����3��<7A �uj�/��7��������7f/�T_p:d����D`�щ��/ɗcH_}	uq�����:�G�	�Vj�-v*ȃ�N~��H�Ep���Qё�.=3�KFh-8�Qo�3kc��t��������]	��:��ˣ(2~,KPD\��0�	f�i����� A����x"ߺ@{J� 2Z�c0a�2�`w���^�'"�0�>C�@��FS[���yp�M�;�d�!�AQ�r�]���ֈk�O�+Ub��ɰzS4���>G��3�Mz�B���3��������ܣ�ѫ�� ��*5ׯ8DD`������c�;[��5�2�s���"��E���C���?S-�<�tة�e��T���m����J���>}�Xv�=֞R/��^$��_�̅W�`��غ<�$��SC� �v�߂1j�m̫7f?*��ic���xw7'��U�l�r��m���f��D�f��b�ez"�Zp��O#�[̙��ܑ���ql�Sna��Z̘�ܜD�y8>������h�ΌBmm����LlE��;����͔�B�&Jxs�����F7�mx��@�f9\ڗ8\=i"�Rb���$$?�&h�q���g0'���?�+e��2�4ŃY������B��t���h�TG��P[M�	�]�f�jxg]�r�(6Ɨ¾s�Frǣ���ᗵ�d�;=8$�=U��4����s�Z��L�R�^B�6ߒ����d(j���V��
~3�~�?���-y�%
��0F���]C��� }7ʮ-��:��q���Wzs��WqE�a��qơ�c�̭�.�]g
|�$Y\ą�k:.gR�-���*$�`{���H����X�� Cg����g�
Dn 'N��'��v@���	P��	�@ ��n ����X�r�������&:*��Y��SZ	�هB�=�P�V��@����i�-E��C�d\��z�����2��Sɍ.��|�	r&8_�����n'g�n��"y;/�߳"9��N��� �ksv#8�=%�;��)��	�D۵�������Zd:u��bR���|{E�8������!H�$�e�,~����x��u�j����;��zZ�Ux�"`8j���̶�Y�z���Aw'P'���񓵃?ω@4�W��C��;��6�:����D><8����▣U��]R��(�u&a��/ɨ� .�X�L^(j>�p���&�XB.
� 2�\�@�M�
.|�+�:[ߍ��M�5ec�"K����a�Z������][�����(|W�
Gd9I����wY���0z�Q�J)������l7�̸]\:^�5˾��ޭ���{t���5+��]%[��]�����N�Q��N����N���v#$������ˮj�D�@�?U�h���X�9�,X��]���X~�K�l�������>�S��ȫ��^�*��+@P�L����l�N���h5IM���oOe�;�[1�*y����5Mn���S ̲]Os4v�r�X
�	��щ�G�����J��yB�,����M?|�����<��WFɢi�+$�^'M�0����ӈ+��lۘ� �
��y#�b<�
0G�����~#�N�o6��0D����w�7�6���d䐄���Fܫp�l�S�ǖ�FOXݟ�ߏ,�=Pm�ⷆ�c)�s� ���ջ��UȁSuĳ�t��~2�:DV_N�����+2��&&���@�ҽ���#ꄲ�_L�mJfOks�~��� �c�K��zf`��6����P�F��V'����\U�)L����ʮ�pG^��;�y�r9�B��P �H���'��Ũ�e� ���� U��bm\Ǉ
�Q1��E4��c�yⳒ6��|ę#� �O��?7A1��D�όj�N%���l��C�%5�'��=�l"������r�G:�DbjKc}��WD`����)╖{�����pk�]i�&5�C�$�FiV.��Z�R���H k�����,/E��������&x��k�9^>�#lo?�����E�cm�u�����#�zļ���3�8z��*Gd�m1�O���	l�����p�1��ZթBy�*���
���B��Z��� ��{:*L��w��&?��GN_�Z��jn�*7�х����;���1�3Y^Kz7��4����Ri� JM��N
£@�T��m�X������tz�����%sr�t�'Q��ul�+�3N��[9s��s�_���Nq.s�k�K�
���`�$bT!��I�5�J��Q��oy�X,"�d0�X�Ǜ�@�k�o���*Fn�5Nv5�<d��U&���/kM��>�|7(�A��&���b��M0������r�CW)��Rw�B��l�$���1���rC���� 2N�t��*�= r�����5�Aa�4{��nA����Z���w���rm<��E�Ej�%��$!J@ӏ��X82,5�kR�8�l$�;�kL�7gVu ���f+1D���t���@����8�l���� ��~h&��RT���B��^9+�}T_U9��W*�¾�݀��	��6���k�='��es4+3������dl/�0j�c_�-���)�X�7������BAݢ�&;C� A��	���������n��O�E6xfH v���
�=0(Y���M�Va�|d��x�/nې�����G'��Q]E�}���nTY8�MƗ.�
��o9���	�&Na�_x�ݩ�`����x­r����4��yR4������nݭ�|?��/�#�˽"g��7R��ԗc�DSk�(X�x�#\��oA����s�pM����\�B��4ٺ����yym����K�$a�p��[XdQ�E�C�۪E>	�H̕EQ�\���W�x0{�b��&CW}���Z����sz��;�T{1A��eB	(�wO�L$kY@�)�"�m���+���Mo�+{g3�,a��g�� �_�حԨn�o�S��F�}_^��ɇDc@������Z	�#���>/]�)d,���;����H��H��j��G����j�g��2?Ӗ�r�M��@uvv�uZIZ�Q�]
����e*����X�hFB�)�o���x(�0�+ �L���<Ďs@)N���v����\GҌ���5d��F������8~6F�U�3�#�LMO�+̐� In���
�����柨<jE�UT�K�Q5��zR[�Zdv|h�C����S�Q-
*�i�#�;��F��d�Z\�<�R��C��3\�����#����;N���%f�oQ6��L�q�,C�ėx	��G�օw}�fK$J�T�f���"�����3B��ҌW�C1 h�k�cH�t�P"��O�~Cέ�7
xni��
ꗆ���J���cx�mb4�h��a������8ޅ����ղ���p��<d<�=-��V���쐿��d����%c�rZ�t���M��2G�W��]Yƻ/|;ֱ�	s#�)_�{��	v�5������~�X������&�o��j�h��X�oLgu�*}5n��'H:!䂻�)�;�y��S}��;ѝ8�b2��x���K�>H�Nh�ï?��R�TKr)�W�(N\��\/�8g`��f(���od��b��@^mC�������(���{�l���G[�V�~+l�C��ytF�����%����͇�R�A庥�'���
�mk�,�[�#ʽ�g��YxT�sWh(&�z�U���)�?keW�So��|u	h_)��3O�(�]��Ř��+�<h�s�I�m�����(we�멀U�F���Qa�a�]LдWD�S�%��1&��ƾckMoE`ථ4�F�����s�:���MGw"U} 2�����.�Gh� P��U!b��;7?~�?a�Bm�V �c���C�-T�it
�,���ԫh��9���'L�|'pYe޵�Ҧ�T�z�{��ă��Q� ��"\Q�,�dN�\P��i��/���ܢDj���¦��JQ�{}��	��ZE��qXըY,Q]
,'�5���g!���v�F�|�/Vʤ��CD��e3~� p��&3��y�6�Ԝ�ڃ�xᖹP���7�v��a��N�w5s��`�O��x�d�1(<��9�@g!�7;�\��4F��&$���
G�γ AU��u��7�����^��W���ao�v�l.����#Zܤ�@�r��e.Gap�F3ڰ��G��<��+����)c��Jj+F}�kڜ��:4S���ͺ��?aL�'=z�>0s���tH��2:���uCx����}p�z��C' #F�SL+��m`τh;�qQ���"rd{j�X�_�g�}r�;�ٌ�Y�Ɲӯ���U�3&�  ���Rx���GC���W��� �7�$}�Á�:�k��:�x?�����O�=�nJc�|U�~P�u�-Ԥ7*/�m�%�MAX��Gc,O��kmE�fLݮ洳R�E?��Тu�X������I������v��{���~��B � c�<R��J�B����n�)�%��Qo�5�D�b�)��6��������Q�yq�Af+�9d�S5�^"F�N�w�%{�2�[|&$�
wv^bdb��7w'�A	j1g�qW�'+�n
���>y^֤Ӯ����eŏ�'3;���^�簯`1>%�V5<҆���W昼���h�D����(�{����,u$ؕ�g^`��� ���P أ6��w�̹���y����D�ͬ�~s�.�U<y���pdg�2��/���.��I�\���`T�5�Ґ#D�E�j�@��Qk�������s(/��Q����Z�2�c' >4�wd:t�>9�:;J����=����~��Ձ^�&���T��b�簯��$�l9�lq�O��תF�g�^��Y��H¥~~��:j�#�<��y[�v�j�(kt�꾀EP!^~9Z	��ll�I�J]}	�xI���U�����y�%�dר���4q���$���P��;$D�@����6A���͋O���Fr.b:��幊~*/U;P�K�,��T�u����f�$���o�XQ��n&�nw�^����iȇ�yUI]����=���j?�����`5�-n��Z��������?�ڰ��F�B��&rY�o
�ew8�88qU.��!lbr�hF״���K��@Z��=}u6Q�:o����1x�Y�o�).��E������h�	�K,>�^?g�ڽ�^X��T�K{Vv�wl冘��ז�����W{�cN!Z	�?	���`�������uhgii	R�f�-��F�5n?�t$�(o�\�v_n>>=�cC>��`#��xZ�d����=Ʉq}d��B���)�������4����⿬�m����qJ�+S[�G����ϫD�l�����<4䟄
�}�+:�lӤ�M�EW&��r��bv��P[0)]�L��F�?��2C� -��rf���݁���°}�'=��u%Lӗ?&�z&h��V��̶Xn���:Q��i!-G?<�L��v+���,����yX��$�Pվ�o���ܞi3qeH�#�����4��D��@��x����7Dݧ���Bv*��̾�ۅ�f$�/��ꄰ�X��-�����s��4^ߍ̲��j�
v�vv1譪=��sk�{�CRv���8!y��c��t��>����w�̣��$}�y�ۥ�Ս"�l�Đh�sm���y�Q����� �� U��Q�zM�/�!����~�g�2�5A��f�zQ�����FY`.�jRO���jn��~�n��GB?f�/��h��pC�^G�J�ݡ_�����E
cq�yZ��n6�$�e%ѹ�����:�,��ۓ�H��
�1f���j7���V���2�Ҡ~A�B�y��G��P�@/W��d1�x�p�?|���"_����#=�頪0y���K
�Uv>�Lw��K��f�J�cT��n�֊n��n izu(ƪ1ܑ2�����E�F�����)�S-A-�̸=�H*^�����������=�8[�q�}��:%�Hx3���9���5]���X��U0�qU�o��OA��<Yqi%����@�6�.����l�8�9T�����A�-=u���Χ���p�п�&;�G�*h)@:�d�Y:6l�v�C��<�5��t�A.����FvlC�wj���}��,��1W&�дDa݈�KY/�J��9�s>l0�J��&�z~��������0��Q%�Df�!�U!j���H%q~��a
��;�\\Q����-��墏�IV�+r�҅&���)YU	Nr=���_�0�e���e,�F������p�b��:��; w�\.� q�4N6���4��-Ap;�4��#Yna��r�A�_!�g��p�O�w�=�F��g�S~�CY�% �$��Y>o�\��[���+�@��p5EL��'�E�(��S~ t��CԘ 
����l@L=</�F+�f���w�%떭��i�Abx���
k��骗P���j���� >�0^�z�q�I��N4㢁[���u�����:�,b1�6����B���Q�7�/��k�`�e�#���4F�����M�����W�!�1�`��k~<g��Wy9���u�m\1Ci)4����yp��?�x!b�������\�	�ⱡm�둯�N��4_͢�-EKfX���).����P�r��n��mS���ٯރP�r5���Nv�xs�ɇS�j�J�}����G���A 	iٷ����l$�A@��uv�Ķ��>��D��{��T/�,Ҕ�X���w�,�����`�c�
�����Hf>D*�.��Y��]\x���{����[��==l����u�6����b��b!BgӡO����P�� F��<|�N�r ���g]2��g��g�����=oZ���ϡ��Z����F�� �jF���Ӊ�b�����1<_��,��n��d�,�a��1&��EU��CUn!&f=�D�b�mǀ_�� �� t�>����[�z�	nRs�$J����4u=�_�+z��#��Ȥ����<%��L��<~� &o1-�l+&�&�����v��eI�j�3���|;���Sy��07Љ'�[r��-�����@�Kt�'D_���g���Sf[0N3b�zoy��`�2�f�Pu�*�t�oѻ2BD	ZB�%`x���R�g��M��MG	��=M�u�+T�����9o.3�a��ʔ�V2D��6�W���ڿ�W.���1x,r�Y�@���U�7�eūka����h���c^T��X �m��~�#�^qb���T���iR!vWs��Zb~�k�I��I��~�"Ɓnp��i
��ů�W�%Ű`M3UIHBZ�upx���\4�+�)d$���;��q��a<	����i����߈����7��������l�S�����M٤��K��䩕�N���YJ���W ����N���o�^Q��@Vi?zh��P} ����?�.����]�����k8���Ҍ�	��fϚ���5!mL��.h�\��*��
�����&���*6r��Zu��c5M�(t�x#52�n?��5k59eC��� ?�}�'���U��rf-KF\���u6[ʹ�����ۅ�§��I
U�!�5���=�m&��{'=���Þ��$�Ԁ�k�/<�H_DGd�%R�*l�X��*f�?���a�	��}D�A� �[u� �OIՠ�K r�
O��a��b����jv�AS��7l#��RO�|���T�Шܞ�&;��o z������(O��k�<w���\�����FQ�}T�bv�Gt����f��8<�/��E�t���0��ُ�r�u�l������Dֲ��(�a����O�砾�5�G���v�Ъ��y�>R�Y��:�B'�ߜ$jw��q`FC��?L���b�"V�&I��D��E���1��ۓ���I�7x?.��=�(�ekdcqj�w�ңșc�7ՠ���%�U	�4B��t���eK�u97E���wi��z����#%��U�h�ι���r����}���?%�>@%�t����:�'���F���~Kev���H����h��^�g�;���# 7eH����e�E��)p�Ȯz����^���MсM�S�#1Zg�%4��`t�8���ݹ��Knl>�X	M�I+�}O��~Gi�jV�%�F'�hȹ\[��i'f]A���V�e�Ͳt���AC��S"^@)i��=�s�����
�����R��:
��c���4�}X��Fb��וj#�����$��V(��G�㯼������Z����6"0�|꯵f��;m��P��/,�o7��X�Λ�C��w��G���}9�π�i7r�����,f����J�,�}��(C��?Z� ��=H�m��0\:W1
p���O����R�o?���~e��HH�e��f�.�3������-9�ՅWcL����By/CY����:)�,�*��j��bg<i���v�R�D8���O������M�gd0u����N5h�t�lB{�.�p��介��eE�|��?R|I{n�g2W3�g��៕�
�4`E0SF��5�f����{ ��A���!��b&���kļ�����gv�(�
0���T���sf�'�\S����b��1S5�,��M~�	5o(��!�*Yh�k�b8�b�a{�-�F�pS��0ݙ���*N7���n��$w��9Q?bR_����sc��p�4�)�TE�Z��b)�,����.WPuR�E;02�W��ȌV����x{Jydh��.4����z78�Pg;ui&���OE�*ƭu��i��tO~F�Mz���-�#�79�O5<������V�{>�H�Vю��K�$VK�c��d�$�W������ۛǌ=����	�:������,'(�����v�Z:��%B���jQ�S��wM~z�˘7��Ʊ*<����U��5n܎q�^�z�(�\���i㪐�> �������_R|Y����*���yzIiu�%'�Q�ay.g��.�r�X������*�46d ۋ�3{a�[ͯӤ����.�)-}�-��OT�c��ܓA��\H�;ۊ@�V$0[��,��~	�+��}ߏ��Fy�h5���b��"�4�qĥ���*A//tZEeX��~���Jߏm V�P��i%�gޒ�J��L9\��z���*�1��YY�\��#N�1X���}��ڱt�G[�.����~I@��I����3�����c�~|���X,k��GwZ.�\d|�Bvl����,ͽ0�`2k�y��Ç��-�c���g�0�20�6\��lUј:���i�t���Q4�E6�J�AZtz�'��v�@f�"��-A\{uz$R+ӵ�����3��h
�4�1�I@���~0�M���z�H\��z8�� $is��왁	�2�?S��Ȕ���?��T��	t��?�}�|ӏe�6,4�fb]hG��d���xf�(���<@��9�0�E�I�2��o��evd������J�Z��e�{�&�]Tkܱ:�����:
 ��u0&��K),D�-��Y/���t�W)$x�7&!� �M��:>M҂��ae�:kz<u_��|z#��'둄��]:Zc�϶OCB����?v���b;L1p〢�EW���B�������h7Ξ�)2DW	�N�D*��P�w�<aɝU���6��iEǟ�hL�(��!��蛍@kC��P�)Gܽ�|3M�Ă���&I�<X�g��\�׈<vo��Ob�Q�������&Bf� ]�X���� �E6���B\I��}'����P �m��K�b��
��t>`�6sT�^aσc73Mq�'3�y[�ʊs�~�.�S3�%� ��蚜���T��Y��t�d��7����^sѳ�~!���!�aeg���c��s�G�;�� �\��V��Q��\:0FYl>x�[��Iq����@�A0Z#�o��Ezt~��f�|r�M�^)���f�p�����*K2��&���~�������BC��?��嬁���;x_#�]e>S�B��*z�5Қ�@k�O)�W|/=�>'4	��2��$ۑ��1���@y���4�t�*�%��D4B0�����w`+�W�(�xYc�Z��2$W��1� J2U�=�7__sx5���rX��*�`d�6�!�� �
���7s�ͥ�� �ŏ�p<8��B1O�yQ��4���?0�x����I~�x��'9��e��aGV�;�݌_�Q�ۂSq߰Fɟ���^q�z1�@�,�C���ԪK-�]ٿ!O����#�-�._�)��"���[9�?��E�X�ptq*]rWK4�����$G�P$Ε. c�7���Fuv���<_��@2ǽ׈xt�s��)���|Go� 8nO�۬X��K3Į.)�Y���S,a�Ć~� �5u�P8��}�ԑApO��9��	����`ڥU��W]1f<k����|@�
�:��]<��gR�/w�.}ɦ��仁 E�X�� &�ʹr�㒡.�i/KA�u@M�0��@lJ��bn!ۛ48�=�g۷V��F:�ŝ�cV�&�$	??�'��U��غ�NշRk�H#QbZ}h�6����o�i��A�aK��0��NTl�:���J��ר	�� �I˹��!*&L.��\r�2�)
���=�6�>}�Kk< 8���g��G@�h���Ml� �����sp�I���fij�Ư�`z,�me����I���ut�����/��'À1���G+Z��M9w����㻚�Џ�5��]��U���;#��9�����X�dϟ���/H�')ae�y�m|�y���l�k�eO�7V".�ڔ �R���4T
?Ԫ.i�3�@�/i������OSԝ�����А`��	����z+Ǟ�p�R�f�*�#���$�r�����_eAu�ɜ>�Qxj-������ʚw�Ja(���3��'``���	Ü�e'�t�_s;I��+e9���yp��/�(��<��톈�H�15�� 
6���I+`^��De@,��-�h�z��OO8S�?z�\p���Ĭ�-֋���ԍ��ҁEiW���
���z���2w�ܝh��v��)�pAɅ����b;R�Y�!p���Hv/���j�i�0dJ~������Mż^uBC7"���n���=2�!J'j�':�.�E&$h��CcG)��LYt%�\�xl�. V�`��.�K��:�(���8#�0� '���K[d��r��:���Z�8�:/ޛς��P�g����U檵�"�-�մ�D�8��\nt�o(ؼ�o�U��L�#=����� /�D<���~�BsF��7v��++��+Ç����oڣ�M]/v�It�!�ڞ-�Už@��t�� J������gf�P���E�b�mޜ
�ƞ)�z\��D�Z	�O��"cɲn��VPF�����Ca�0������@	�	��^�b�����p�8Pb{��ts�������劍>��������$�=+��J��s��>ܠ���8�;Ee��v;����)��8^A�v�n1S�$߈5����2�ľ�I���*�����9>%
CY����#E�*�����!�X#��~���L	Y�z�rQ��=��^.ݗ�����A����D�
t��q�1�	Xg� �{��/+^B��Q�ߚ�z�>��7Uɒ�dưЉ�~9+��{���?�ݙ�\�����K<VИ*8r�s�CI�\��4�l�Ru />��ou�vl��cG��%��'J�]jD���*j缟�}�2����(N��;IQ04͑�;R��!� UX��~�6eT�9�������4Rm">��ԲN{���2u��{���Bk�O��?�Ҍ��Ϗ�9"�X����=I�`�,����?��K�)�;	��Q᳠�V'��9�$��R|�r�p�����u����ۼ�m��~l�_>x��VW� C��o�K�ro_94,<1�K`��	�NyQ�z����͸�3	��R/m�] T�ߵ��2l�a�8���g������5��L6%τ9�p������s�5�1��Q��T:'���$D��ƹ����تTDk����R��z��K��V'1/˚wK��BFH"1���h��<W�X{�g��Z��]�J�hhB�����8K]���&��Rxq��n:�����&i��(��I�! �wCi�����b�$��4�=�+�R�H��CQS^�*���m�ۘ�n��Q�9�����W��薥W�� ^Ed�1j�}���6+E9�<��F+����BK�I�}R�0?+5&ǡ���?!�����v!#^4�oLA�E��<��ۊG1}�׌Ԕ�
�u?�ŕl,����7���W'��Pm�7�C��!��6�w�{v�5~�d��,̼�N�M��W�r#�8�����.���v���=��qy��2���M�wh~��
hx/�}�6�?2��^7Dx�O@f�oit�K�:ҝ�=B���(_�+�����k0.�������U_�̹<u��R�2_{�6w�{Ӥ�B������4Q�) 7)J��%Wf���������qq�g�'�Ӛ	I�堠�Q{8t�瘯��4_Z�8���`�?ŝ�#��Q�W�43��nMH���]��Ȫ���6� ��f�y�&�N\�w��j�	/��Xn��#�r�O�����rI&�S�jFrSxs���M�F���{+�������4\b�zt(!w�OC �@{nW{��<��8kϚ'�}+
�C����}���-"C�e���ᝥ\�����Yo��ZW�t���g�s�����{E/���^�P��Ϊ�_�f����Ԁ
nc�5ﹷ5˪\��� ��#��y�(5;Mo�ס~ |��{狸�T�.����Y���x�g^//����au!����Ő��Ɉ�!Q�iM�E]Gz�#B�����ʛGO��E���s�S̛�;;���rM]��
k
�x����b�=�5;l}�I[��4�RT�@���aO�<`a�cD����>��;�I��'����#d�k�!��Yrћɉ1�a��1u��P$�VZ�ʴ�L/�$���DB����n �q�/T���آ������Kb�P�pc�{htO=�.WE^���?g�i��q�����B�0~!Xr~��E]��/��+��`��.�o[4�Ģ1�B���/��4@m�fV���C0"���ԙl�j����Do���������ڬ"��nLJp[�5ws p�m�]'����J���<q~��<�&�vr�F:,��1MKXg�޴��8ԐU���G(o��3ı�B�xuY��ˊ����a�L4��"�0"�O~!�Ȩl��l
�J'WD�4�]���ѩ8:��!v6g�YA�/ٝ��H?L!-e�9p���[���h��u_��Tc^�N�	9���r��t�@��q���uu����E�[;4k��ݼ!�¹
�P_��b��\���*6G��&s?0�0ps�M��n��'4Qn���nB���{� �tn�\ �t~��71��H[֦��dj�HY�V��Z�r%.-v���U̎a�n�HL4�
v�̌�x��#�/��]=�_�CAȊ�<�G�p�W��>�>
�ƴ�K�����0���}�	�$@X�Ĭ�-	&�ܶ2�7��ȝ��9Q�v���� |�.���򳈃��=���D���ꮀ��@���H�ؿ��d��\:��/ ���Nn��)�x��ZD%M�9F	�׌䫟rw���~�ӵ7x�t4��v�4EH��?�a9)�����E%\�{W�C���/X� ��LZ�Ko��o�����0�T$M>0��&%@��OMk"�3�C}�R�CHS>k�h+m�Aw�״��A�j��҇`T�u\��h�����0$�ү�a�!7�]J���K��^���ߴ��va0ٚ~V6g��[���sYD$ и3�qɱ\�on%�{d�1�%������4��HySy�.= ��d�m�о�pbT���&��>*V+�9��$���ڑϛ�ȱ2+�o�Mx�U8e�~ͬs�{��#��ǧ������(��`e��Z���]=
�jՉ�z�/�r��T���Ka	b0�z��wK��-���RýAG��HL�S^]|DV�ƅhD<I�7W���}�@"����W�ϗHzm�8j6�5�m,2���h�>gF*z��>�PvK�=0�����n�a.,�(j*_��,�(q6d+�e�!
:ṻ�3�(0���S�����Z� \?�ip<Q�T}�mC�� ��QV�"�����k�3c�1q$U�_�t>4v��Ⱥ�z,��x�M�<!1�y�_�W��P\������+u��7��%��G�pʺ��F	5��W��9��0��=
sx��xA[�bw5w]�|ã���"_�y�4��L���U�ޅ:1�^��?��}g"F��ş�#j�>MTU�ؒ��"5�$�_��ԞT�a��J�z3,�ۡ`:A2�+|����x��z��А0s��s���rP�����t3"]�Q���<�d�g��?�fP6��Y�4ݯ�XU�H�ve��D�f�^�v�5?d+E�h|՗��=��W���bY�iSGD�ddL>��&����o�������5�>-g ��wm���	t�����IS�n�g�G����
rJ->���1���V�w=;�Rq��F���\�Z��6,r�����c�AE�e+�:�3�{��;�h��W<Sڑ0��k�՟"*Y�9�;p�U�*�ͫhy��W<!p��{��[(�.��RdÊ^u�j��(�]���p]&	Ǡ���Yo&K[�X���۱��k;��*��Y����),��'�@��/�p��ce/w�@s0s��;�M=��D��+�lK�Wy�%k��T�*�'Z}�=��a>Y�S�
��%�:s�?*�V���8�:0V`���=s~����C�9m}���u�!�{I3%;�z� �,�}o��׍˟Td���9/~��SUC�F=�p"��ƻ��`KM(��1�/��E�8�[�M{l�1��/��X_�͓��Ǎ����Z�G��6���iF'�(d��sXf��2|�A�(�{[��CD�����a��u�Q݁.����g�i�p�BRK�P��>���S�~g�5嚧��B�h��W�|.n'�ah4��5��D�C�>$�1��Q#J�ms�p2癣KK@�����}�P���'3G9�D�L����zTY��T���F��>?2B�5M��d�dQ���_�=�։�Ⱥp�\�X{��̎��@���9�1��g����D֯�;)B̠zEDPZi��p3���ו��+���Q������Zb����b�X'\ ��1��u@���7�'��3�^_:�>�$���7�6�^���%�c
��W��$��FK�	?o��&�N�Z��J7+�SI;:m?��/ޟ>�G���xF�L�R
Y��X*މ�G�"�QR`�`] �Hwz���|�x�lg��A��:�4��S����&�u�U�B-x�s����=���J�$�����\48��IΞ�Fe?߈;0��~�@�Z��T;�Ih.=�Z|a�B��d�H������l�q��GR�%�
�<I?�8�/�f���A�zWr9 ��$ �uh�(CL�E�&��	�Gt��M%��,:�8������ہ���-�� D��<+�D:a���%Ջ�I}&}�*�&hzy�3��F�!$�k��� �YJRu��--5W�A7�b��ֲ�S�QB�}-�Ŏ)�Oz��ے��Q�F+��ۣZ<��ʨv������5Щr�71� ���M��ژ8���x��)�Rj�w�kFq�xdz�46æ�I�T�
Wz�2:M�,�Y�p�]��n�w'�d����̲ӄ�b�W������xҽK���
(�JU� q��ģ��%�����[ДW�]��u��Hr���7B��&	��u��|&8��h��;�;�u@�`��/�(j�q]��H�{X6N�`'齴�k��6'k�$볱݄5&K9�8C����B�@-Wq��:/4;䢭A R��c�g�:w�O�U��i��ƪ������S���x�(�:��d|�i��c�t-���B�l���*��b���p+��#�7��l��Pt�=n��)3j����y���ѩ���L;������^�r	Ҫ�]�i`�]�/~����l�1�is3����ƱD�f7 �K�aq��0�Z��@ݨ�8r[ÀsZ:����� ������ؖӊ*Xd���K����t�Ga�إ.��D�����h.Ҫ�#�ym�<�|��@����P#�*Ѓ�BG*w����J�!��fɮ;���i<K:�uN��pu��^]H��M�箖}T��Ʈ��� ����t���`�=��}��c��#�$���
�h �aV�̓���p��۰lO�!��d��]
O�Lђ�+K����3�}��#ɐ�XA�ɤ!6���ϗ>��@��Ø��t�d+��iVa�����@���7}��3\�R���buA>o�V�]r�����$�Ɗ'�e��HUR�v��k�cIP/��@#*���"Ɉ	3��t}���yFA�1��(af����{�b�ʵ.�\!|�a�98ǻ��!i���u̷�<�k�t�<���ǽZ�YWl���w��;�h�Ng��n�8�ŵƚ��"M 
ܯ��J�x�-S})+�˨WY��F�5Å7xV֩�G{ͨx�١��t���(���K�>�bn�~�n��Z2E�ݘ���,`���l5d�#LQ�U�c�⮤�9胗����b	����EON����:no�ܗu�a�*�O��
t�
ҷ�N��zP @��C6E�ُUҰ��mG�J�k��z���|�HS�p��m��Ġ�`�>K����H������T�NР���3���;;�ޕ�����D�˙�R�f��^���E8�(I���qUN,��ސ�5�Lp_�C����5όwl~�^]��S�O���ⅵ��*��7�"TY��հU@a�Sw!޺��=9�������=��5Y��?�D7 $|h}�;��dޏ�v���G��X}>�>#�7X��fHRu�f�+E��#%�$�] (��>���I�����$��$�' Z�4��4VR3 �]�H3��1G�C�2��r7�O�p�k�hZ@������Tyu*"���U�G�G�a.0f$G��C�7�K(U��\5�}m�Ǳ�9X����^������x�$J�p�Q"뇊��)� ����l�X��9$���簥�����V��0��>#"�p @��x��D��r�������:�o!Cm�a�Pmvך n�=G��^6�De����wb�oY�\�c��Z��e5SK���
Ǳ➯���,�ADq�p�]�&�a��a!H��G;.>��`=Y��S� �lu³�;:;�5Q>�ر
����1�$4��9����5�!3�e���?����4X`M>!�[cE9�ivz��4c$z�7/"�`���>�:�pP�M2�R3�\\�U4���.���d�t:X.��=��Q��u��'�r����J��2E�qX��ͷ81�����A%������9���z�j�	T�\LɌZ��6PI9�s�4K����P�0�W��\�a�wC1�D�]G�Ct2�}#o� ��&ƨw�s9�i�.��S4o*�&�= �� )-Y�m[�V�Wf� t��q�Bc��j(<ӑ]g~w�Z�X�BP��(��g4Ћκ��gK�BQQ]���7ťA��T�M\x��>����F�fQ�P#o�X&�ܔ��Y��f��S������m
���^E�ܟ�$�:�tY:\}1����LN ���	��F�r�2?���i6z�Q���$�ݷ��1�
�׎��;U�i���	��H�Lɭ�`侇g��O�X�U���߾Z�4+\�{vo�(�i���b0E9 �#��-$��i�#A��#�nS�h�V`��B{^`r��.��~�*�gSgu*���� ���Y�e�+�(V�Lo�2�=y/ބ�koכs]Z�����S�T*4a��loS}�(�LXvԢ�	�����py�M$��Nt�����������渴�Χd�vVpC)HV#��Z��vIO�g����ic�\�Z���<��ϫֆ�zn�� �P�:��x�S��Q�:�K��ߧ_~Ein�VךW���A���Ϸ��R�8����\.h�3w�c�jw;�_T���Z��׺k�Bt`B�b���9��G�b@���1��B��Jri|��ue��,r���Z#]�mv��Ob�E7E�ypn�5���� h�t`e����`���f�9zL��bQ��̛��ب�zڅ�a�%G�����I��p�}EK �Z�(adĩay�g�Z�f�O �~��bbtn�D@}G��`LѺn�c�c�(�t��l %PCR�"7rJy�,bYc�3!ښCZZ=�m���)�QC6"L^JYF6�V�;��o��hG*X�=�N&��.<��nhJ)'�5W�`��M�����%WL��[�%�XC����	 (��.�Iv���Ӵh@
_�r�~M��.@����I�L˝����ķ�0����[3ϕG��4yv��W�-�S�6�]h�����r�.*��݁a�����[@kf��.���911owj@Ovǡq1��{�
�~��Ё�/`}�������˚�w_�X�{���Y�B8N�_�;-���ů�^j2�G^�`N怚�%�="��`�DW(j$�6�'T�s#z��.����2||�N��f��L����2<"��mvD�lK) u�����1A��Z�Y�Q;^�&Xz���!E{�����(D�r����dnP����vv���fO^P<?Tt�2P�p����,D�O�{�eFX�u'il�Fk�z�ws����	�C?y�+���[��\늯*�O�bp�஥b"���p������~��dXU' Dn��_�Ȁ~)�~���E���2ǹ�6��°��
�vL� m\��b����%�W~
t"����	ӣ`Uɔc#KBSyX��%�e5�566d]�{!�m^�����J�1Ж����Aq��@�G�b̖�n�Y��8i�ELR֭���Af����FW7�t>N�\��5�O���0�˼�}&�+�iȧw���f��Ki�%,��2�[q<�'.��	�.T�Xr֋>[��$�+:V���Oa8�_�܏��&}�Yxv��{1?µS�$�4�|v?�u�|l,�ܬ���a�
��؟�� ��]2��=Ƅ�ct6G���-��wlbHD)� *��(�Eܡmc����m�?a�B��M�t���i-jZ�y�.�6�{R��p���c��������Z3]���v�ZE{h�&;:5j�#f̂w���B�^��9mA���O�8��k�.�7�3l/�X[�UV�߽�=��M�C���xE��y��_
� 5�W�S\�4ұ�r+�X��jf�4=��h�U%��#dj��-�8z�ٟ�-��7��_�kw��Of���e,25�tݎ�-��[�}ʠ�i���
�F���f�?�N�[Y�$	m�%��5;��a�T���Ec��4�(n��s�����Ė�s�!�j�(p���H?d��D3 ��,1�5�	$�$m�P��� �k� �]>V��͘��fJ��W䵹y���6J�{�ID�%�C����VU :���t���2r丧l뫮�g��a�m����-6����+���$�����i~��ψ<l�ȗ ()_����rq�>��m��M��ƍ�>k��L�Z���Y�6�/��(�∪:ZU�s=���=�^�^:ν���_c�a�[T���o��O۾3@��`�
�#�乲)P�O�Y�t�V�Tz�����r�:�bf����_��v�]
�8��$�0��X����L�57%�\j�1,��+������VO=U{��KD9�,�)�k��d������/���=��A�u9�=}���Wl��$T�V*6X��1�f�C����χ�"����ե{P��͕̕q K��L�zR����ˀJ#۴�����o^��0H���^�y����;u���Q3�B0eـ��5�_��ǛN�ex͖x�[x!xF<N����n�X>F��O��e-�^�C�;��XcwĨEJ4�}q�1�\�2�i�I�b��$.f����_@��z�5���P8��L]�dx���a/��!�4�\�.���}2ԛ�v�Y䱕S��.~�h���.�a�ҮCکs��s����l8�Uϡ��8�&�`���� ��C�醂��?`�&]��MV�L8iPG]�Oy0�ь}*�3��M��_�w�b�;��c+8@��Mj�6�o3��D��|X:��}p�^5�VU~2�2A��/詽>�r�`�9��MиY
��<��czo�,��ժ�E9��N���l}�6�ؑJ��uS�{�d����8F�o�>��!� �~X���lr��#.�hf�K���BX{B���E���.hJ���$�Q�����IN}�08;E�d� ��%#��T�I�2�:Կ��������J1�5)��JR�2+�zX��K��/*�J����(����E��J	���p�����N�Kq����S���g����#�l�Q�����=�G�8C��9f��?5K�s
wX��CRʌO_lO�ę�GOM͠F�E�,��ȓ*�d�T�cS��.�z��Y������rl�a-���c!:�p�_+8�����(�<wT�3̷ڈ}�� 1O`k��wL� 5���!)��}%fB���G�hwN�:Q���{��py�Z�;���>f֨7�Ʃ0{��U1V�?��r��@�~���-��C���/+��OQH�;@?ؿ��X있
�����U�|h]iS��P��V���T�ѽ���k�A��.>����_��8l\*g���Q��c�C�|~��J���ft�ds �I��yp#�g����qP�[/�}��o70�ޣ�j���MB��G��.�a���L���5θ��<�;̞6�)��,��a *d��O�\9J�5*��;���A������f�<��6�-������ǫ�`U�o�`H��U�i����ˈ'�����q���c�jn����򂯙��"lо��k��������ˤ6�(+���d�P]!Tg>hi�9ro�^�g���1EY���jMK���LҠ�O��=`�[���g"#D~�_�"d��Y���]ʉ�!��)�/!0��Q�ʲ��å�g��^�Ynf�:I����iH�]�=IH��<��tj�?N�v���'�٫#��%�6JE�~���*��T`^b\H;Gì�O�a���]�ݴf8��e��x�{����[���Bs�DUaz7�"j� �[��'z۔m�mv�)j1K�6�.����p��:��F-A�L�Lu
�`�B/TI`��CN+�s<��t�,�g��+�0=9��YY��b�n��۝�-�`8vA� f��V����d�Jh>�u�o=���f����RE+kh
���?wWc���vE�iM�G椥ߝ��P.-4~��<�ɩ�3����>��3-���N5��Z��:�uE>�Z���jc���]ù�-�m�L�U����N>���'SAe������C��/Xz�Q(�d̤u
Vd�A~1�.%i
���&e���`��o@�؅��BG��(�0��{��@�|R������
M-�䈮�'�J\��x���B%��/�|�@���z�~�dֲ�&��Ӥ����x�Ex�"�BM����b5ޟ2�*��[�ͣ�[�S������E�h�:c�#-5�\l�U8�p�0�c�zA�$a��`2c�U� /�BO�ȀbT��؂�F�&�Y�g��	ZX}.��1-'0A
�C�S]�lN%fI�\ԛ��u���v��IZ*��P�:q�kw�_��Gמ�ѓ|�r�F���W6�g�Š��v�J-a]a�)��δ/�B���&�x��l�J�ai��:�P�Jd��iD�������	��"@5�Q��4���"�i)QCkv��&�^��F�D�!����$�uLh�
H	#���#��!�<ѣ�=����nRI��Zl7���hR./S͓S��S.ڕ&}�V���k���T�p�f?�m�G�X��r�*N]Ee@FF3���8�V��7�ö́���!^ևO���֓]��R֕���
ua��%�#)L���FնQ�x�<U�$��Vw2���
r����y�t\�!t]����\�b5r�L�wj`Lá�n�BN���3ʌGP�M��#��)���_��=�\�/�cҤwp�aT3`-��.��{q�کl�����X�d�"�)ަ4�;0�ސs�s���q����n=���͔7_��,BYEXY6:���Z�B��+l/C_������i+��`,U=�>���H�IgM���(e]�����j�%\
t	<�p�I�{����!�ېf;���+½l{lm�_��*���E�h���OH��Ъ0�xF][�rm��z�
�څ�֣����iD��9ذй���Ͳ�u�&�8xĤ�>x�n�_El��#�tRY�d���K���׎.�H��DK��7~Chm~���m�얝���W�~b��ȣ�E6Ⱥf!���_���{�[�Ō��q*$Ch6t)k����,Zd1	����Р�
��]�:2�I~��bP��1p���S��p0��x��*a���a5b2!��V��U�&1��T��K�<�����|ԦX�\_ �M�����* �NS��0�P�ŧ]��`��ĀqP@%���thIx@[�7p��[[A.���4l�%�K�x�o���Kw��mS�ue�\f|����P�������z��_]ÐD���s�݇�d0�|�Jj�p})0�:��8e3֮ӗ��VIYY{��p�%��y�@e��x�{�V m��GhϥѨ�ƌ$	�O���ORE�_�Ԛ��9)h����`�%u�Q�#���I�J��=z|���UGm��R·��x�(x�[4U<d4|�Kx����TE��I��&�9��-YҬk)9��?��T�1v���I��B!�9�!��y@�w��_AU���~��զn�]Ͼ	�a.�2�I=�ù;�~�p#�F1��&>�my4��L���p$�;���=��u�9�?�<1�,���qji��8b��%�8t��cW��zV*W�E>�-�Z����,�#o�|�A�Y�6���k�Gΰ<�����-��ߓHZ�{�b���JD@ܫ-� �U�<���2�6^W~fv�ʌBϊ��]�q.3C����ƍ*����Z��1݉?�l�ݒ����2 �
b �kt<���z��+�%&�]��S�<p�|�%_���? H���ۛ^UeikF�*=,
����|�\۬�;~�֡�������t;7�W��s�$1��AXWс-t��(�2�wV6*�EoԒ�Y�3�����r.}K�=x:8 ��J�X�ĸ�K�R����N��.��U_�G�A�g���>
���v2Em������c5Wؐ���P�YD�P�b�M_L�:񳍴ā�!@F�
QJ�4�|4B�^�q�� �[���a�z�ӑ�S֎nE[�e	y2S���;u`���z6���˝��L��ŀmI�������W��tN�f:S{κ��?�!������H��=Jd߂�����su�c$��ȱ�2R��4���������+����ԉ1�,0w�1��R�i۴Nf�7����'zŪ4�
Z���o�t�4�	��(]���~쑅����L��l��r%e�'���%�R�$>�%�%�����BcW�R��~���.@�@��Nez��kKz��6V�����!��3��T��z��zZ�k�1��Z����� eo=P5�b\~�ϵ��ڛS�ʢ�i� nd=P
q�2H���Ӷ�L�(�|Xb]Po�	��wߛp�?68S-���ޤx9!XE��0=D��b\A�_�8���_��I��/a�
0����V���yfO���� ��^�g�$�L=�@Q�i�MC�B�ga��PތeV��lj�L�����r�у�8��˯��(0�]��	�����В0p��>87�
Q��Up�P.��#���ab��ͬ������( `km��Jq��E��1"Z�ĦƸ�ݨl�)Ź�O\j;@־�#%����	Ā3 �h���ƕ@eB-�;G1�⺝�s��Lcu��2���>�ID�:�Y�k=Щ���=�_\E�^�x��T�w�*�W&rnZan�`�XG9!R��Mw�Z:;9:���Bl��_h@��t���v���[z�d?��fҐ��V�{�j�p;���V�lK�T���^@����-���Qߚ�95�e��85-��hO2�� �K���1F����(��2*��{��OG��g����A7��o���2�K��9���w�Ou���jf�ϡ��˗⸶D�,����;�k�3�����i&[�n���I�W��!.oc�N���&�R��@*�M�����?B�gs�NPQ1N�"����o:�M���-�緉��]�GL.�*��C�"���ۥ���yI��
<��;��2��rk͔��E�$ߨ���7)�`6�&'a�x�k��D�h�]�|�ۦSV���!z΁W�L�S���@ń�ϖ�F�?e�W{���q�KB�,QT�9�Iv@#��C��]}.,5"��r��P������tUh�����4ś��s:5�J��"�eڙ-��5�F�R�H���.���wxbT�)�'l�]d=��^o�`H��=YC"ߑ��б�,����`���)X՗�U���Iˤ"�UЯ��n��κ_T�3:�Q���&�ԝ�=[���1�9�,gd����<���g�/�.tc�)������ܨ�yi�5�4&s�N@��
�82I���Gv��?�Ag�*T�u��(0�K���Kt_�֬��>O��Y�ƚ�x��B�ՌA
p��xù�+9!�h��~���b`��$�& ;��DK�V��n�<]��!F��$�e���v@�G�^>8�:}�_��N�Խ�j�j���u�"�t��))�&��S��غ$[A˚�X�}G��~p4N����s���|qC���Gт��C!���l:Ò�!��]Y�S��T��;B;mJ���}�[�2��˿�:R��I���$tt����Y�����f(ʤ��&��х/�1j����.�&����������wS�Z�_���nP�:�k���W�N��!>cO�t�i�bSL�����Z�GЊ�wX.5���|���Q�H�|-��lھ���>�v�d6K,��3,�z,��m��u�.��,�	L�y;�G�� #��5�P �&�Z����$w��?��e�Չ�����{bYz^+�4d�v��nyL]�8r�̯�Ps�O7�,64?�������Hʸ ڹ����l�=���Am\�;DS��g
��S�D�07<��<!��mx��m�̡��p�r�qp�|�B����%,��Tv��l�B�ΡAO\n;��!	��2PE��qB�U���=w�L(]��m���	A��� #9���7��WOg���3
��*f�q>|W��dV��9�1Y�����t\h|}tV��aH��{'��+;��b�vr>��k��Ⱦ�h�
���E�8��݉J�j���?O�]�7��y,<*}vj#�֎.���'�T��X��}�A3�����~�|p�$b ���eܺ އE�%��`�� [��+Ft�ٳ�������vM�Y��9�5�i?���ä��VZ�Z=?�Z'�s�$����t~ULۭ�g�5�Ԏ�io�c�!\y�s����Ƚ�qG��)���h<��X������v���lݿFD���l^�)��¸�u���<7A��������I�2�-�L���"�e�Y4�@J��|I��LY�ы��W�:�+k"����VP�Myf�`���̈���$/� m}�Ɋ9+~�À,5�|و5�^l�\[�q ������ �trF�#�LH�*\�nC�9������i����f�u�O+bf�.��M�`Uڹ��gó���v̅����wZ`1��^��Rd��Y�b;6 �q��?�{�%�_���%P��ׁ��ʏ2��^)�U�%V�G}%�A����?}_u�;Y8A��:c��N��+˿�\2�X!�/�<gk��CW��4���j�>-�)�M	�Q��Ӯ��A�Aa2i��O����R�9J�]��
@�\�M~�>Ѱ@-/�㓹\����k��W����`�?�W7�L���;�p�B^���o�N�F���%�K���m��g�{�
|���;m��a�k�������@�_}����S��(�T"��:w�g�~�ƶ��(C� �p����I��(�<�G�<Z���wƨ�Uq�3�j1�L��b'ɉ��M�o#�;��%�ɑ%J�H����n�|] Q���@j��|�4�S�	p�jt�>$O���0����QP��tJ����n�f#�f?}8
�b�P���7�*�d �Y�[tP��T<l�P�GZ9>��fKb7XTj����J�d1P;�6�C� �Q=��m��<!���k�����>nЄ����Q�����x}�_�dw�m8�0 ��8�������p5�AT�)��X[$i9�?���YE��5��[����I
�>TC�F�}^��H:'�ʹ	.����t���@D�4C��x�E�\֟�v����,JD��ۓG,fA4E���F�x�_�ξ���~��X�9�RYȌ֨��P)1E�ٽ��w�g�ױ�.|vn��=6³̉J�aS�hje���/���r����NP��vv���T���Hx�F�`��������S
���|F��	j�6";衢|ݱ��1g�؂���v�2;ȸwVX��j#��ǝ�ƌ��eC���_0��3�g �X�u&�P�%Q���T���Qcp=ܔ��\Zfݝg0-�V�XW�Ô{�A��f���;:l�L����n�����%�[��`�W��֢;D�'B�L$��u�zi��5����y�{}A��M-�h��Dq䊿���6 ޏ���l��t}������7 ��E^�L��UžPK�6M�%�q�ϓ�-�
�S4c�e.�E�G��;��*�J=�p��J�1�Tx\�\eQ^A}������������M���j�j]h�s�͢꺫� 
p�	�ϚqJ'��o�b��_�^y�4��ğ2�%l�)$HB����&�*����n�Xn��I��.�`Kh6E���O
�خ��S���I	{�Q؄�GJE}�O��������IT
f�wC��plE��:��	ɳ�J'���x���Ga��2�#NP����q�_ M��
�r| ���O��Z�S�k���i�����@6�q,���a�L�f#��v�r�T�ہGe� ��]����E��+���h8!��@e��������
g�Q=����%�nwaw�k aS��Jc�'1@�C5Z����Up��u�|vh����SZ_������ȫZ�m��g�9c ~���1�_�j�h�I�¨��AO�t��l��=��,���R��SN�5M��`�!�e�#��s;xC?�:�'bѬ�%��u?�ޖռ2�2>tPGm��N���x�x3f�4��$,�f��)����Bz.Ȃ08Ɔ�+B�X� �;'zu軤�s�>��>e7��G1GD%���~pd���j�T�N�����<io�������^��[k.�T;5Ս�����Wd�)]���4D\�v�(�T۸%����!8��)/I*��f�6���B"�9
c�[��$��G�m+�q$�X(hVD��+&1ّ6H�śҹ��+�9I���N�ͦVR�P	(Sr�|;��)�*v�-2�d�3-�ݜ����'���.u�h�/O��qu�������O�T�ɗE�A�xgR���x~E�E11�x�Z�۠͘��꽆�;�ӺWF����y�7��ͱ��R�T�3U�>�C͐V�3�k���0:�{KE�����,GH�����7��R���@o��J/����|��?gI=u砉Ʈ�S��g_��Ӟ�6�r	W��b�E�k �-I�[�����?LG#
b�R��o0�X��t�#�>݊r�Φkd+���r
ǂm�1-����k
�u�MySu�Q�܀im`��;%͑�/���lm�J�˱�9M�:�]gl�� � b3u.#�Wq���.E��t�p�}���1:A�5!� ��i�z���7��/�F��ۜ	w��yp�ś�G3Ѷb�LJ��7z���)Y�����)�9�w�7�ݒ�, ����EZ*�̘P9���>F` P�uA��~e�#�Z�O ���.B���*$��({w�NLɦ�<�[�ݢ���k���
R��֯�p�T��~b���+L��h�4���E��A��sLSB�!��$�޵�)L�Kn���!	S��e)P�Б�s�G�Bxg)D8������],zTt��g��~O�w��r�d`�����i#,��Z�ݭ{�
HY��{4q����.s�R|���Ѓ3���;����F;� ��$%�d�8�l���/�L�Ű),���������P"�g�%`���w�z=���QOc/��dgZ�7���̕i���!1Yl;�7�blٙ@��-H�@��ΩD���ԣ)Z���-~w�k�Y��� (���e���&�V80؁,�95�œ����������x5r{+t�	!6�\=Q�|���z�9��AD��У�޴�2�����F���qzȖ�#q"�D(_��ȇ��o�8�H��9(�W����o�N����Z~8q^��j�mlAqI��\�#�Ɲ�Yn0�j��/�&�l�vqn���/�*�k����ʠ��ѱ�g���<�}�g�f�ik��\�U��&+J��*ɇW�/Ŗ������HF$m(w%f3^�b�:������Xb��� m3^$���٧S ��.��>��3�������&�KAK�d�(TƖ-��j� �dH"�ъ4��A�1�*-]H�6�k�H�wPi�m� �u�z�y���Z��R������	-Jo;��W�m2�ُ��: ���Q{6� ���U4�?��i3��
D�3�R�����k�G ��qçea�{u��-���CG_b;��@w���QW�]��nJK@%,��`�����t>W�d�r�4>��/E���)]��G`��%7��T�-	��l<<=�'��PJn���^5���c�;m��+4U����Kޢ��8�SFc@��/�{���&)��c�<��s��c8����;���Iqlxdr�GG+�[ƈۧy�7�&�H���T|Y����GN:��49$/Z�}�!vџeS�̱�s�Qj���ڰhu������Qn�"����f�uGA&�!�,]?'Z�43�%xC�)	DĸC���tSm@�4:6ȿ(�%���r��1x��u d�cQ�^���p�ڶ�?,��{_H��-���=�v�n�|D�(�u��Hy<��p��|��Ȍ(/��L�.vA��˰ܨor ��ަJ�3���R�O�G v٥���DOb�B�U�G���6���5���.z��!,�(���I�����hJ*��S#����wO)��h��gi�����Z��F��)���R�[K�!��
iwg�
�]{S#o<�sw��t�EH����NV�wC�Ⳉ�kȮ]oI�	3�V�Ny�cՄ 9�yĩ:�%�ؠ��T����u�Qi,������,�qr{i���MO�
U�L�9m�)����6R5j	ٮ����H�
��X�:���),��T���Q�=Gh�q{� $3�=`���^��q731]��\a�Q��ʏ��av���7F���g(�W��j]2���V����4��
������f)U�K��.ͤ�D��L�K,A>�p(0CV�a�g� RI���*�������|�Z�h�SUD��@w�[�����$�&��K_�������%��D�13�4k"=�v{
�� �[^M�P�F շ���u���C�R�Do��]��9G�r� �;vO�gqo�r(�?Ǘ��InSJv���]���q�3h��#))L7�/�<��$�DFܥgSg�4=��'Z3�>6�uV*.�x�Ԟ�a�)�m�h�}�8�0H'N,Sg1O>���"O�`��k�+�k"�`u��ه\�J�z�	����}Poq��8�w�r?��T8���91U跩���Wv���{=-�8K0�'~��x�_;��X���K�4�����۹]���j�]$/Օ��㵎+���nɕ�K��?�.�
(oi�>*�9.���Z�ނ�,S8��f��s���'�3oE�C0P��2�.N�4]�<58D���.�Tn��o� IM�b���8�~��I�:ξH07Vc�
;����(AC��Н�F�L�n��\|�v�������hB욳zG7�.���
�;I�0�	�- ^�X-e���@J���"+h�슄����)�`��@�G;Qs�cH�u�L߫�BF��9��>�z�82[��G	xJ�����q�V�2��Z��W�FG��i�@&Hˁ�9�L������TcV��C�H�r�b$�~���,$.�n� 	^���|�a��O�.뒅�hMn�y��f�]O��%��r���%!P#'Z`u��7�<o��*�/E¼�MPw}q��{��Iޠ�Ev��u����yG�o�83��1}"�����F�@��X�9��Ԭ義֬�{�j�h�B̖� n�tvu�·	U��VV%��M�6���;��r�$j������F�R''�B��#4�=����M�Z==��{R�#�)yo��-S����6�5�(��F��#�	{�k���]��pP��[��d���8`y�q_Ζ̿�TKڀn7��
�{�/`�\��-+�bhj˰{�
�2 6��'�Hԯ���CZ-ث��cA}#F��j���^�)�o�	T=G����r��?6#�/�&J�s\�
2�ф�v���tU����S�����]mo���ŊQ26=KV��q	T�:F�Z��CЋ����X��N�q��z�[<F���!ͻoٟ)�.e������nc����D��QGV�
�	ڔ������N����2t�>��6u|��_�X�4u���b�^r悁ޙ��]<ˁ�<Z��č�L9M9A�M�u�CYP�?FbmG����/Veޤ��3��*�j�$�JP�d�Aw�`*%H6[+��p��]do��UͶ̘�]=�2q����?� "��P�Q-�1I�1�&��~��	
t�3MLڏ��|4���T1��*�aI�<7b�Ke��}ou!!�hbcFPc�Bg�P�jT��V��%5>���T?�ַl9�[������tR������ɲ��X��7�!c���pϫ`�|�,XA	$��hf���Ҽ��jx�O��?��-����r(�:��`]e7��i���V��d`.?�i�Ѧ�&��@$[���Mk�l�{�A5�]�[�K�}�Mb�ϰo�_�����p�+�B��H��B�կR�:��l=�YL���X�jI�S��1��f{]��T,Z�.2mҎx�2�`��'=�×N[���_TEt������N�n�r#�7�������GW�hP�6f#�f�yÅ��y�P�5eU$��D���8����ٺ����n��ig���]u�����d��/�AAW �8^�,�eW������Kؿ�4�� �K�9�۞��x��q|k���)RH��[��&���	�<�Ɠq��;�	P�k��h��$��q�#B�S�(�f��F���hkY!h f���m"o�O�g�BC���e�����y�B/�V�"OKl�'���}S{�^��td��:Z1V\Y[x��_�7�w�ݕ��Z��,~m���r\v)9�����͜�n��m�#�	yw_���@���/J���9��y�?{�zxb�a��/C�k�@ڜ}��IQ�b�a���i�?���Ԁ;�H��}�b$ц���䡃SsDbAP$����Hۀ?��u�{�91��6�s�pd��-m�s�߳�/:��])�$������q��(���~�6"`p ��3.K�\xP.�V��|��M��f��f����[��Ϋ��"�V[n���m_mNg��@�di?������%�ln*�R
i��>Q38�w�g��t�����1�!,@V�")�}���l�p��F�6�4B��ã����=)goA���Ã���<iS����[��J����ȾcD8D�2<��N�]��MҌ$��9�;��{YuS�7�vA��2d��/M�$�F׀�/�=vޜ�Q�Àm�&̃91̶�������g��0�8�i}*�L"�F2����^;$�f�oX	:D�-e�c�Q�~H���=�I��P���z�V�g%��ĩ��y�+44H� 6�P&�?.��8���y��Tl6�'!(m�	�y{A��)_�P+2L�ʬ"BG���QB.���X���Yg[7��E�=��G�[������������I2����O�n��b��s7�8��3�*:�&Kك����c�[�[�����A�Dzx�~��o�����R���������/p�(z�A�k��և�ef��EOc�D�����Elc���Z��Ґ~ܺ��8L��`�AF�ws����4�5�G�؇�?�M�/8Lk����)v��n6a��;
��<�{ ��C�����M���2�C�p�g��e�Z�x�bq߬"~ fḤSz�b~*�V,��c����˵vz
ᮕ��l���V��m,�(�d�xH�Fpk9�,iQ&*s��H�ŷ�x�. ?FA��//� �O��Z�/����U���r�Wr$Cf��r�a�-����Q��S�ʉ��iT{�c���X)���wvD���[!�0t�,y��
RW���s[ԝX�bK,5�<���X��q��!Q�s�:��&���$��`���ڬ�O�����EҢ�Ѹ4����I���3B7f ��g&⧃�6
b�\]��غ�`���{�y�����/aߦ�	�/LI��Uפ�:g���	?�K(|���Җv�2����!�y>F����Z�p������+],>C �4M�/���vh!�wz�N��*<wx�8Iݯ�R\,z����x�w�b��+�/=����4�в�����7�p��*b�
�](�/)���o�p�͋����Pf��}��57_`һ�p#y�7�32�.|��F���W�9�<i'�f�)���;�Y��~:�F�&�����1�(_��ų�F'��{(	������#�E���:3��r� �
�3�$ݢ�6��O�q���A"ċ��"G��/��-��
;��c���Ei:��d��?���h	�/�s=E2PA��`�\er�
����$��+�]e�Ր�V�&N
l��X.�A("U:�#��p⢙+���46�������-+�(U�	7�`ߊg���s2=G���<��[�V���7B�3뻽�&��F�5�n<,�5$jK-�Jqŭ��!߭��I@�����TdfȚ��٦(��ˬH ;k���;�!kfO3�63	��R&�w��c��Я"AX	�yr�e�oGA��5
}��f[��'�e��&b瀇߳l����%ph�F=��&��	��7�x�r���긔�Wh7ۈ���~�qBTGi����Ѧ#�`��~U�G�a��S���5��O��O���3K�ll�P]��;��k���L�z�� H;�H�!I��I�`�~o3��2yi�� 7+���pq,���6H�5ܙe�(l�y�\�E�S(���'�n���)��l/�+�Xi�I�=��壌���G��6a�s^65g-���'�̥���P�/���> �����,7}(��Q
 �����=�GoZ;�����
�X���A|i����B�U4��1x؈(?[z��Rd]p�zG70�
�,�򭽪eɨ���Z,��`a���O�~9d���җ'���cK�\��n�$��!��1?��@9������rS�\X�/Jgi ��h�Np=����1?"^-х
jY�q�m@(�q�VЩ�/��N���u��������2K�^�ҧd�[��f�ҟ�?��IdϹg5��{�r<E��څ�䐈��R �.KJ��rɄ8_����Ӵ���^���/�5���hR͙������ȚN��}�v#�w��N��m�B�ر�O�Y�@��d\�R1��ڷF�D��_��2e�ڝm3D�⚆)^0-�;�r�R!w���s;٘nbe������w���⊩�N����o���dU��E���{�e:��1�"bL
�m��E��Ҩ!Jנ�Y�0O&����8H�d S���~�fO�	����z!i��:��(�\�ɛ��_��'���#p����kF�	ִ�\�lӏ"��!��規�n���r�1�vy��m���B�7��0���|��/{��~�z�c.��:U+�Ky��ۙ/(a	�=�}�����M�$����w�Qy5�֭}
V�$�}v���_T(
I�]�7����As
��s�K&A."��eb���;��:cf��!�`���0��剭�+��=bn�eW���t�����;O�ֹ�!zP��N��Y�F̆�d�$#���~�A%
��t�h�M��4s�^��7QtZ�c9��O����7�\{�.��3��-�4A-�
e�x�%���|vz��8"[����!�T1R�=���bG�VQ?� ����2�xxY�|�s�@�J?������r���U'��|ZA�{_�g�6TDֹ�MA��c|
��L}H�)�-�k[f����Y�^��OO��X����k\�H�M�X{�,�N0�]�a�2��Q���\�7Q�!I2�rb2��L�	���`��|d^��й>(t����AMԐ�Ӵ�Aw�a�T�c�i�ܞE"G�YiL�_�ə;LX��@N��q�R�^�elx���8>��3i���ݩ �|���O�v9.;�Κć��d�!/���a�/	|��$h(�<������Fغ:ƣ�&RA���D���~dU�����.����,�2�3{����� �����:vR�m&����ҍ�N(�(�S���*A�
���0&��E�3�|ܯ~o_��c��D?�"馬;�[��M'���9,�I��$�R�F۩��Oj��-��{=^��U	{��,��ǵN�������V��`Goo���A��^˂��S��.-�E��]�Rg��O�m�3҅N�P�������P�����x|87M�y�~��1�3���)Fg~I6��b��'��|k	�ϊ��� �t���b�9���F�U����7M��N_���}_sؔy`1�ճp*���6��/�[�p�P}� o��8����Lɴq���d�-5��x������|�F��}�2�E�Z%��;�ǡ�)��/,><��FU����`�=e� ��L��g`o��%;�����)h�JRS�8B���bp~�Ғ�0ǜ|H$,St��?���J��N?sıw��Ծ�u}�;��!���^X?�8v�P�T�A}�,4a�$�ݤ�����@��燺zS�\ٷ<h\bd��I��%���X⤉d�ƊL�:0���n�]�i��5��~�T3��x�����G��*)QE�xJ���+nF��"_G{�ឩ+)t5�W��o+�m2�����e������@r�t�}���v8:b���0Z��Y9�5Q3�co�-��w�ƽ��Oӻ�hd�j��g˽��⛽���z��<$^|(�&��Y2�K� 8�G�}Lć	��~e �Dsy:�~����D�xdD�'���x�o�*�?߈����e� ��a}����є��Vyvg�]�9����{D���I��V�M���lW��y���>\��e���\�$��sj�������D2`���V��@0��D��o���g�`�Bh֕N��:=�u�!�q���3����nbh�� �ܹmDs���Z|���))|������������f��m���$�l9�����~g0�~k��]�����3��oҰ�T��M�Gݬ�$� �L����h�u���A��þe��,�h�JP�W�.�����~����x�Ra�?�o~+�p�i�C�Y𔈐��ȉ�'�aT��B���l����՝�u��Ԗ$��Șּ�`n�������ߜ��X05hЁ��e-Q���X�@�;��,�haTɇ&�G�޿kON�'��/<�x������r��B��a(O�,Z�����(�jS��dKcg��iK1{<��!n�X'5HUOX;f��vԽ����� �>/Ն6�-/���)��H9Q@�́4����4��y���ܼfz�����9��C��&����/K�&L`��Y�"4,�WO��Q �6�R�ð�!�)Y-�����
��",����C�+��F�H�!!����3c�w�ܾ�wD�/Ꝥ�2��.}�r����|�O���>/Ґ�36U�h�1�}p��8���D��H[���˖Re�H�^�?Rcl�y�⩯e�hyui�f6�g����t�D��OODLpp�du���IA�d�D��*7#�x~�����Y���ߗ���ȝX'O@���6���S�d�`�Y�S<��$iH[�v-U�{.�09q�b\
/qz�q��̉���o^(R�۾�_*��m@�]݁�^ˁ��"��胛�M!�j-V{/��C�O���ɲ/�[�s ���\�;��W�Vnx�ѾV�NG�cn�djj8��ŧH�#�Wh�WB����yU��P�[*"�䫹}�$'x"}�kѨ�]y��A���7���Ï����Eo�a�i���  x�@�Bi�^�K�z���:F��D��j��"��l��A�yMm��yO���@�|i^�܉�e�6U���pর�T8��M���nD�N�-0ak�z�bJ>�{�T�Y�^'�Z�G����\2�|G+�3�űj9��D"|�*�����^�7k7��Z����Q���=�'�}?��<7�h$/�2�}�M^ �We��6O��Ãow��r-�t;�+�X�y5��͉H���*=�w��#4�í�b�F��tb��������Cݲ�����c���g<�za�=b r��ɯ[�����xXI���Nb��e�g'[r��ҵ�����c�f��[�la�Փ�Г���$q�s�����'e��[(u>��Rě6	�N��fq�p,윳�^m/�P�������P�G�����������>K�~S�ɂ#b��_T��!�$7n��ȳL����_������4>��<�S��g�R���Fa^
@FM�?�oˆ1�Nm+���<b��BP�kk�T���e=����$,��o=+�o�0UB��(}S������\ն���kc}�M�G'+7�#=����PE��2V�|{�/�uw$":��dy���{�^�]�+,S��	a}�[�)/lߙ���A��%A1�AP�����T�2��$p��WʥG�9���#j���Y�sڳ�v�,pQE(Yf��Z��#�	�\z�dP��D�x����ƪ&D�6;Q�>��or����W��"���w/p�w�qh;\���#m^�ʤ� J�N(c� ��$����I�(��yJ�W>XX�����t_�x%�᷸?���$���}?�
�j?J[�&���w3����ڹo�����ؔ��f�_
������U�<��F�`}-	�e'�ǌ�.7/����,6�a6tE|���=���E����O�F@�pͱ�z�؀�ǝ����:�<�Qɣ�"l]�0���`���p�So�k�v���\p�}E��&�����X*�\�z���6t&�nU�[��ݚYD�|��}����2@�,����A�#<�`f`��Q)�!�pn��]�[�벝�:���4X��5
]�ݻ��8�́)�0J_٧���T̋&շ.��)k��Ɛ���M��Aq_n��q����%:�����.�^TF�7�<\W�rhr�M*YF>^�6���o��ȹ�<�5E�[g���o�^�X�.CЅ���-C�}��`�ٕI�Ԡ�mO��R-�g���[[�tmD2�4�v����W"��#�������_r>�ZȒA{u�.Cl�n��Ήv|���2���m�52FI���7B{���'(Rt�5����R�
 ��>l���|�I��9�c*L�ys�b��RLwi���*�pA36:�k|3͍[���y5�Þ�_Q��x����xP�`�KG���q�zd4�d�E�Z�E�)u�[�<��Z}ùЏ�4b��b�R,Y��Bd[��uO�S�G��#�hq�A���E�W@l�#%k�i_#�`���%ݴM���y|�t��(r���o�<Kڙ��u/G����>�5,7�7E��8<����ȟ)q�v.Y�
+@i�[�Ȫ�;`�U�����OP�|�θ��|-��FEA�����x�X+���R��`�e�Poz����������h(�rDOqĪ�\(�}`SNRup��?���\RYE$��7��"�~S����vXDo}�_��G�m*�l[��1��Y$�B�oz��k�����p=���S�h@	9X�
G�|Ò�Fǀq��ϻ
R_�3�V���٬��������kV�Oo�����o�8t��|>X���S1,�)K_>[1fӸ+GۧԶ3=�0co�&����G����Ǐ��SSaӕ�6��ܒ]|��U5
�_#�� �S�����b�>7�՗�Z�Ռ�6t�����cP
T�3�^��Nl���=��,=�QI�=��J�[q{�!�E�����h|�'�xh9K$݃/b9��8�O<�)5S�չ�Y��,���&"��˷���8��g��DO���'��'|�p�la"F����Z����D���V��z���X��ܨʠ�
�a��#���{u��s�f$dȞ�\�s��ۓz�%��`��D\�(������v- b�@�@O
�5sh�w��'�����_@"�I��9�����3��۬�j�z����w��r��-��)��c�����2�]��B?��|�Iqd���!��
��YZ���#�fc��E��,�x]�i�c�c���R����+(���r�3+Dj�_��e�c���U;�{r5�T,��O��'Kdq<�e�	�Q�"�_+6@
��$#�
���8�*�g���6�Ҿ�w��;~�=b��U��O͔�VO�4v;�0�o�_"�T��w�h<}�3z�݃OY� ��j4l�>y}��������������fܳߢ�a��`)̭�جVU��%��̲�UX6�m2M'�yL W!�Ψ���32��5Q9S��E�d����!��y���^����_r
q��-j쎑'Dru<���/SQ��x ����'ƪ���Q��-������E��1�o�q�rZ�ˮ��G�YgZ����s�B �!�ܲ1���������Ǳ�<Ʊ��_n�<��ʐ��x�~�@�7)>�t-W��VNC_u��[˶���� ���Ө���΢Ve��acp�W4��e�scڍ� ��
\�t|��$�}�0/���%q2z{�m��WǊ�4���;��֬䴃��)�����ˋ#�G%.���뜚���I�����-��׌uv���g�鬃50%TK������3�ҁ�v�c��&�1�o|[ ��``����ʈZ��
��P��i���tB����U.��k�4֐ߔ|���o��7����9)u��Y�~�~u����7�Ѩ���n{�u�=�U��_)�A��7���pFc��Ry�K��.F?��N
��&�Ǘ60c�a�%p	5��'�Va�L�����:7���:~�l�s�{�;��oaou����|!3l ˬ}�`24��@����c�g�-�|jR�LW!�	T'z�Hcyٛ������V�r@8_�Qg1А�{ک
���Q(�X���U�D�&�ճ��L�5B��N�=�C��nxmU(9=��h#�r�F4PWX��u���!�������	�fb8wLQ�u���rx,��խ_
I>�!�m;D;�J��{g�OZδ��{+7�I�6Yg_��YU����� Z�9bm�,�%Ǎs�+�I�ޢ��-�|Vn�����}�Q>��d��L��Ɉ�m
��T��0��:J�kS	�`���z�>O�܀��.u�MF+�(�t(֎���Я��~��tlݼO͙��F-k~��Ѽbro�v0 �u�EJ�.=�U	R~+��U@ ��08)Rp����D��l'm�%���W�����߫�&����*�DPV��F5?$^����Z+����N!�kJ���I@Z��X�Kq5�l�����e��F����T�%��\5�/Y&w))��ˏ����(�������˿Qɧơ,R����@}̥[oj<\R��-:F��G��(4N��\)�����cq��w:G2�|x�[_O1�
�|S4{1Z-s��:V�&�4B��@Y�y�I��3=ځ$��Cަ�(�����"
�9$���GNv!�d�T��%��jN���.#j<0���i� ���q�]�򸠠�:a�L@	���3���QLó4�q�����T�Q���e���(_��E�����ɩUp��w��n��.��|� �d#��=^ɼ�E�j��mE�ƣ���DK�-�II���-O�_�`���(&wȶD��J�\{."���^M	�շ� �]�R�''�8ykN�����h�U��x�Cv�r������<��b�锚���Q���w���0t �
�!_�b[�8�*|l�%�}�F���o!�=�{=�wX&��H����U�j��bT�EGN���1Y�wI�g������E��q0M;c�e�X�?otBAs��ty���y��^� ��]Cj�q��321��wO���~��Z��7V��lո4k��@C����r�42h�.�(� P	6X�Z镅Jv��J3jzY^ƗI[}�C!����޳ԟ����}+(k�L���(�B3V:~9�ۺ�[��e.��q����,/������u�[*13�5=p�?sM�Y��-�rz�$��{��`qe�bW�9f��=����}�c����i��H ?��y�^�!�"���S�Mס���g`i�� �[՚$�&�Ѳ'!4p@�I��~=�[��nУBH�^N���-{�7� �� ���W�GR�-����g��JT��!aGMAEd�R���	�¶�x.�:�5c��s��1MA^�f����KŨ���.�4�Y�'+7|���A�)�7βE�������ˮ�R��HǦR���"��J�Ϳ;H9���I=M�t��dZ��0u!��u���riCT�fz�F2�}Byٶ���cŰ/�T�9AoC>ZN�Tg2����*��|� ���>eO>��v�I������zC4�7�8���S���i%Rr�9$޼�ed���x���Po�)|�%ֿ�l�H���H������+��"86g�E؝'0w$���+c2����Q&G��;�f^:�-T*�:O�kC$��Q:��+��J��QE���
��ӽcp-��3'5�ޏ���j�[p6'��2�i�T�F=	��	4��K��[/��}��T���~֬�?m�H����y;rH*A
T���)�M(�$£�&
t��7}W}ҊE�ZK6Ȧ_��~�.�1���=�D����ζ-y8K[����V�ɂţV$�ÿ��r�� �Ȓ��0��՜((U%#ć'�1���O�,RJ�#=�S���U�q����ɼ�]-\;L���S�D2AZ����KV-]�+�{�v�S(:|c��Ӱ֘4R��v��$�&���&eF�x��	��d�F5�dem3�jtY���Ԯ�F,�R(B�˖��b���-H�=�]���'�t�� k>b�Y'#����1j��	��]U1Æ�2���
��bX6N�M� �Ƕ�2�}����d��c@�5S�� 3P�����y'n#��ߺ��;[� �2����9KG���=#.8��evj�Psyvt�U��㼄�<3
sً��0�\)8�U�d>�'fk'�	��i�F�NXA��
7�3�`����`f3���� K��q��	��p��z��V�q�ӏ����#�K8]u&����t3'��Ͻ ˟u6.dz"���L8��-�_�%\�����g5�j˥��Y���`�����*���^e@��p�]Ia�<��6�p�ܫ�Y]J��,6��V0y�������N���lK#�Sb��L�����]���`%qu9��^llvK:�w3�b���s�z�"\�%�VA�f�g���3*K�91�ݸ��l��"�0�Yr�a)�$�N�[��i,�Ν��IϏ���ٌ���NJ|�A(���(!fђ�?-	������p��c~���,�%����$�Q��-��R�\Vq�qפ�y.� ��U̚eV*�[�%�D/Y?�C��c[A�E��_�k7�w�Z�X��܄�\z3s��F�Ae�I�	_E���u���tӀA�'���Q4x��6�1�%І`}��T�Wİ�M�7�\!���k��2��m��U��3+KcI�������Y�钤Cr�Ti՛L����5��jU�r�Yk�LoЧ�:w�ŖP �0n揢�Q�]��Y�� ƹ�*��W�������Z�TK	�2���D�S��0��>n8�M�Y�Th��!����:�"D����_�OUZq�뷲;�ȃ�s @Ti[ƕ[���2��¼v��҅J��w��'s�(�P��|�Y�����݄m�-���ͻ��L|hFR����k��$c�T�ŧ��h�%HS��I����H ��_]��_k�YE^믮F��4��8�"|>��%.x!�Gt^6IJAH���E��0g��D�M-nܙ����LҌh��ޜ�!�a�Q��	!x��d�N˨Z�:{ʔ�\k,I������],:�gdqV��M���Di���iؖryq@F3�#t�#B�Z�g����V�$��E�=� ��pz��EK�݊D�-���1�M=p���w��,ch��>5�����*������! ��+(��2��^*҉������x��v��g�
`-����l߽��;ʙr��N�jf)?�&u���ɖ�5�U����22}�:n�8z�Zv�pM�I�u˫d�Y�t1ՠ�k�G���C�Q��
ڢ��{9�$��*�Ьh�Z"��7��� aK��?d"/B5d�a�v�8Q�>����Z,Z��$��T"F��%l���$iKNN��iL �T�&�<h�)f�*�s"O��Ԗ4\*�ƒ��fm�|.E�������Q)�zP��]�{l��̞V��Y��V��Y<��e��_��,Y\ekv�M\��}/�ϐ�u��%i>ȥiRT�Qd��M�@]���O�
�c�[�B���n���Rk��Z;�-*�i��	�Ȝܞ¥���~�FiV�laNz��:$�	)���+F?���5�������{�L�a-�(]�槊�OR�<�	��DiƓ:���ҹԻ������
�i/��N�=�����z���N�UE!��/$�U	��� u���>X(��B�
:ħ���=��q+��	��7�D����,-JB8�ǝ��X��3��b����6��{��(��^����8,c3nay�Qُ]�T?�w-W�`@/�3EP���5`�Q��	  o��p]�m�ӂ͛q͉�����|��īn��~٬>P�>�a��f�׷U�{�*��c�'j0itೈ��M���y�l�Ќu9Z�O&U)Q�L]~�_���f�@4�v�X;�"��Ɨ�]r�L�|8��\>�G[�"{7�r�ṔP��Zٰ��־q�\�
ݩ�nz]M��~$��ikWg�<�	�7͔N�
�Y��l0�3���T�̫�<��_U�r�Hyl��<6��v����`*�<7w����X�-��ueX���#�3"���[γ�缑	~9�R����Yڐ�_��Y��v�'O� w���'mm�����7���A��99�n��<�B��	]=qw�V��I,�#W�T���>��1����m;�F~U.ϼ�CCΒqMu��y[�9�MT���=^��Q��Ͳ�����ʊ+�f(�z�r���ls��o���T��ӗ��$��Ѳ1U�ѽ#�6W)�R�UY�����*�������o����KS�c~�M�ɶ�(4#��	�
���˶?���M8b��Ǯ���}rU����<�F�&�57nؚ��n�"]> 3�$�`���hQ�QSwm�ǡ5��:�%h�8"uO���>S��ʹ8�T�VU�?Ī�gQ�����h(� �#{?��P����	=pJ���1�ܐ����#Y�1���[�%�K(f�u���t4V���r���|r���H�Oc��Bh�5��X�_��<]�[��/��j�$D�L�	��N�^�r�1��&�R}z�i`�
�0�gwE>�T�� I��ձ+��.B�g�^eg��������943�="ˡA�^×��|
Xt�s)���HΒ��YoA��������g~c�&��p�49/�b�=�Yڼ@P-I�\�x:�Vo"\�*)q���M.�������#o�c��ϑ*���7���j�_mJ%�H���}��\�Y$����_7�_ 69Ҩ{Ynҥ;E"#x�~��Q6����q��-���x	g�ל-aOY��O`�(:���4�l��`p�/����wl�2Y���2SQM����*�_��ot�� ���6���$%�āK#}<�k�R��-�Ԯ�,:0���K�r�Mi���W8k���4�$`v9��.	Mv\�wsꞧ�x��N<�p�v���Y��!��;�j^�2kWw?�Z
ӛ
����/Ed�����-�+�ް���K%:�.��$�և�7ob�ܱ�	�cj�Vp�y�B�K]6��_"GA��p3��	7=r�^E�L���+Ǟ��l���-�@��[��)��GR5T��	K���%�Pgvy��(�&��r�L�y�1.�sZ�F�-��̗��q|������|}J��o���#���ߦ�2{��<�yq��$�����5{f9~l9��=}̭��kw��*B��4�
�v�ظW����qΪ})x#EY0���w��V���.BZ(�K>�rR[3e�'j�>n����]t8��q�Km��6��8���~,���U�C��R��ߑ���]
޷����u������D٦l+�Ǣ/GV~�:�-�{o!Qmu�U���Y ��o���4΀�d*�'u�Lu�_��4��i8q�Rc���;0ϥ����B�h,�C�Z�k�{�z��Ly
���t�f�U�ٖP+���Ԡ6��d�r!���"��'�cf�\K)�����Y)�-ZY��"��X�H�����5��]Nsa�*�$i� ���ǇyF��N���d���.��c<�z�P��9����Q<�3�WIQ������ne{�����Me���PI}E���h&��5�:N0YN� p�&����*�z��k���5�'4e["t$|��3�VF5�,�a�����^��VP�����=SyY��w��`U�,{�RU2�<P�S���\iڧ������1'���y�x��r��KS!���__���^j�/pD���6�UR
���UaO�*F�|��.�K��rlm�g��ئ�q�NpI��sZK*u�&��Hrb�eWoqŃTZ�|��F+�B�ZL/�ܡL�N�����QP���&Q��C�BBM��N��m �y�K�پ�Flmx��4��k���_JF�2w��UP���w	g����Q	�����w;�&(��Mee�aJf���9�c�Q�a ���>�δ�@wгn^r�+׼P���kg}a-�E'ˈ�O�����:H�9�D�v�>�� �~x&X���OLmgL ɵ��,��O�{�P�M�<ʣt����k��-O��w嬬X� lE%�b��CT��+_�-`�Q\3�6�r����{��� �![p�/�������R&gn5����*�h��_�w_mG��"�ȯL	���p�?Z�]W�p!��mW�%%z~M��R�џ=��i�${#�p�˥��ץ�ԣ[4qլ�q2e�]����:���M��Q.�l�"�@�b7���Ӫ������^�t`��0�X�>�����Sϭ�/E��B!��K�y`)2П ����C�>ƅކ�9'e�4��u}���-��@f�v�8�g�0��Zb��p�'�蔮�w�I~������Y��ӱJav}u�.������P^\r��Xnoz�afRʬ��y���8z��9+��g����o ��5�Pҫ>mGӉ�Y����A�+pՖ��}�����ա�sr�Yv+X�E���OIՅ�y���Z�:W��S0k߲���(Wy�������kx�d�K����~�O�l���U��C�:'	���A�!�H���E���C&�lLҺ,Y1��.sa�aZ��Ó�]!�4*.�q�~�gQ��=����؈�5g6� �`���aڙ𶿝�E��j��V�l��L�ÖیY�y�|����h�\�g����	�)a�\�� ��6G���jo�#°��ۢ�Α�6Ö�`��%2����q$UVNJ��-�7IԸTt"a����+�͢D4Lq�M��<�a,F�Iv��B���f/{)>�Á�4�^�R"XEiwoC妁L1�_jmdM�V���	0N�gV�A�2��l!����w^B���D���+�BC�ʽLԐ�"��7�6����´Ʊ��x�D\T̃���K~��'�E��l����U��]��	�^D6�,��0�.|��{�>Qp��nx�$:z���o$��س��N�=T�d��X<zr�O1횈�dn{��6�l����u.W���o� S������E��J}�lU������Tn�Hl��+��R۳~���o`l5RLz�����4T֗ļ�NS�	}Q�JW���\[��ժ1��Q@.�����b�Yb�+��F�8�ϹI�+XОo�����iw%o{ ��G	a�o��t��cw*Q����<��EMU�m�JA�����r��J+�"��8eb�g�;q��4�?���Md2~ى]���y��|��#^�ئhN#$���'ƕ~ �����Z��P��h2j�*?d�פL�b��?��4�]JW�l4Y�Q�lWZ�uI�!��9fQ�Ȭ��@uJ�I�Kތ��r#�t�$z��}qHk2� ǽ�N|6A���Mt�*7�z�Mԇ�b���p��1'�ݙh��|{JqJL��r��)ݾ/��Z~��=�p�M,��|�?)n����ݼ�g�CN���!�g���ݹj�K� k�n*oJ���&�J��c6�();�]h�����M*���+�R��/QX��4a��՘�Rc�,��	�2y�b3GO���W��Je_�( d���Ϝ�M�+��H;�ź���E�l�9�,��*����=G@"�k��F ���:��((W���tZ�r#��tHX�\/���[������hM���\c���>$3����;~y@�{���p�g��j���*i���݉p�0,��:Լa��䴭���y�u&����z��7�SU���ӗ�9�.0Y%d�n8[��d:�Iw�*�Q�2H��Q7��Veo���*J����r�;�nL��K�!2�r��p\�XG�ܺ?��Z|0kۙ�Z���P�o�����M�v���+1VZ~���.Ek�eB���}��Vw���Vb��Jh�s�n��Yt�=S���	�d��k��g�����3#A8��lvt:[`�Q�i3)`����D��9�"�����b"��J�Q|*mY+�W��}��f� �s�9>����z�;���]X��(WȜĆU�X�����(7��R�����(��6:�nx���?2��*��d�H|"�(gG߂�� e5>�~ :�s�d�	���X�x(�rh<��|���ۭk���ȏ>W0OFo+��5��0N<�{h�
�P�P`U�����A��n�΅��qx� �W����>�`y7�cW\U#��=S~A�m෹0~��P�p9��]&�ړ�H�Z0�/��R��\RW���V��⣉A�3�"q�{��Q�'CZu�����>Z��rL+85�]��PeE��[�B���m
Ƀ;`+R4W��؛�d��1u�1���7��/ b��,�Z�"]��쪧������
��>�������S�(�0��U�%ɶE���e�XX��
��x.�W�5g�"j���]�2���;\*/��_������	a�h������J1��Q�*�Gg�4�AN健K樅�kM��=�@l�G���������}&&t�y�Ͻ���;�_T��[Z �;A�o!��5L�F�TO��Ӄ(��w�o�@�k���ٿe'�?���f��|h>��F��%�?瑰ښ-�۝�ףuj��=[��{�Hn2�K��yDo��/F�6P7��W?��֣�B��=%��j��c*�&{�&�K衩s$0�[�v8�g��ދq;�L1��6�e�7HY���)9���v\]�0 ��y��w��'�����x� 6��2�u~���/`C�~�!�X��߿Z�,e��}�sY-7Rߨuv�_��`0h�)?v�}�M^V�[��Du��v��O�J�&ށ�.8��d�����F9�^�	!�;n{�AT9�~^���?�+5����{
�n�@sm@��(M_��w�<���B�\bf+j�.:��������t�F^��u���DX��و�x T1��^n�Ѥ��(����t�,jC#��g(���^�R��9ϵ�`L�����9���4,䐵�� ��lA��4\��U���L�[�i�Kګ��>���"{X_�_���e�ӏ�+~�A<���H-yJ�
��Y3����@�2y��;�v�f�n��K��q��ў�C�����w�����}Sm԰S���Y�F�Og*[�O1����+ʙ]���ȅՔĘ���������q1P����%*��)Lm�=v�u�,ɬ@E�0��� ur���3�&�hwVJ]OAm�k ��z�I�� ��5JP�''���8��q*�5���/������4&�̑8�y̑��Hp�a�M��F�u�	m���e�'I,i�h��0i��8�}�>����d��bEB���tQCg�P�y��\�5ّ�"s����Ꮻ�.�s`�a�$�P�o}bI�|f�3Ŵ�u\t9XY�g5)����d}F�n'L\^���G�yp�� ���#eW�w�>��
G&��Χ���s�s�?Ȃ@�Se]*c%h�=+��\x�ц��X���
'����i��Q���X�3�B�����c�B��<�m��ق$
kI<��6M���\��������;W�Z	�_6��u�u8	����tĞ�OF�ěV� e-ژ����ޱ��<����B{)O����k{̆��͖���9!;�a'�qY:.E�D/~=*�� �;���0n[��\~ ]��Z�B���ɣd�F]$�)۟������}º��G%ֹ8��!�Ә?���ۀ���(�5�No�1U����%���.��tz��+IL���矌Pդ?+�!��$�KbM�.Ң��䡽��5&�K#�'�>����岁��keQ���л%�zȦS���ߓ~C����7��j ���@�W�G;YԊ9~�r��%�2���A=N�g&�Yc5$�P�8���{|Oݥ�)-�B䮍!`ʊW��ە�RA��[��q-~!W�i���М@��${`��k�����Xm��L������UaV��%���ﲓ�G�{��
4���)Ew7�{t|�����dX����o�JE��VZ �U$>ۦ�=�7��!�#�X'�4��/�t���-����0�c�'�U�7���H|ZG��B$� ڐF�E�<��ʎ��~���`a�;JHҚ;z��6��Id��Ut�/�	4t޴�UA#���ۑ6�>b���m�a�	�&r3�*N�%�f"ȷDml4��-�;	��l���w7����?�O�!�V�D\e�c�}�:z�d2j%�����9v�G��fԠ<\�?W7��>�'�#ςyug�ʨ��Ԇ�Oo���nGIaY-��-�2.}ϙ���'n���kY��4(�4�R�&����u��A��
�3�D|���Hxϊ{M�� �����g�]���[U7͋�q5��Э�Zc��^A����+1uW�U,��?���@E�B}E�=υ���~'y�~��s�J�ve��-Zrؖң����c�P�JT�K�>"gG���{9M}�-�{�6��̝[*�� �%�th�.���Z?ۭM6�O�K�v_S�- e��l�4��=4�h�	��Qs޿�4*gF��a+?���Ȋ�{�#1�C����!E�t��b�V��E�5��>��cW^��5}n(Ѱ��8S���-���vj���Y�pDs����B��W�S�WPX��"����W#�&1сJ�<�WgƜzL'E���62�#E:�Zz�k;���[�v=#_���p�5¾Z��磠�����Q`(����50vD$v,W�*3L�E���H)v@��>�P�i�����W���堸���7���EO�2��o�t�ĕ}Ǧ1�D͠�8)�g�����-*o�8��f=l\ �r��{������E�Iyu��-��~��55��w��j�ҳ']Br]�z�����jZHٴ���%�&Q>�P�_}�7^�6���J����F۝���ޡZ4N[����@��ޔ/�I!�)�����X����ukaZ-p�r_���ǄC?���]�[�0�{]�~Ze�uP�OCΏB�Q��o�����E�v_� �8o�M{�*����(�O�#�˪�D���#"H���-v8��!t��(�w�5��c��N�K��w��V�%��Y�9l�~2!����U��Q<�FE�K�P�kRwf|�
,�A@��	�PajY���-��?O����:�7��C�G�S�A�����r�|��ҡZ�.Y�m�v�Y��j|J�[�)k���N��t��r��|�h}[8t��%��F���'j�*�J	j����`�O�2_�Bd>l���ԝ�?Ps�Q5����^W}�� HC+^,����-U�c��.�Ґ�ȓ�����V��kj�r/j/ �����`�}ĺ�q����<N-�l#e�ץ�1������.h�q���b��:�<��W�7m=P��#������I��ߝ}�F�5��c�%g�&\�N�'���r�п�eף��L{)�C-�gu!�x���-�J�܀'y���Ha�b��1(>�F8Ѱ�&�XvJo��j��]ı?�F��hӘ�\E��*�I"�k�����[�S�N��Ω	E����eT�*���'\b�P�X�	�ͮ�}��^,�6��h�=��b��U-�Ei�g���>�̪�MT�<�]��q+0�oQ~��������"��h�$64��}_~�� �=�Oj�s�q���^*��{�4C-HJi���N�t��T�ͽd ڿ���5�U�Y�U����J�fT��z�d����4�'��j0CT�t8pc�>x����=���5x�(0��S�%�Y�5��&��Z2L!��C��=���Ґ�B���[/`�s�K+WQ�o(G̿ڈ`I�.*@2�q=��O��7�mL��!f�5�qk`�Q;����Þ~6؈hY�C�N�jOiIg2��� Sd�km厷+�3�&������ � ��]�#Ӟ90�[M__�;�'�*�I⫃�4=@���;�xW����um�9u��-S ?R]nH������@�R4���b۩�#nZ��+�5�O �Ң�������=�Ju�L_����3�7���mM2cT�"�
}�Q�I�ÏXn���B�`2�o9�xPH�lc;η�}�0�^Eꄍ��mk`�#�Mhh'�i�*B41�l^+���TCKm�1�I3�@���Q\��[Os���_b��2?���|�a�dLt���=Lώ�	���Z\I@�[���B�#������ȭ<�Z7��^�/u��)�:�U�kN@�X��Hr��� D0�_�n`]&-�c�	��`��ɝ�3�P��Ok�ypk�M�1ҁ5��OxdZRE�yo����	@�c����=R؂��}\��@�w�uV�?��Y����X���&��YAI�JT�H��5u*HP�k}'z���h3k��pb˫6�ܟB	�FI �%T{���0���¹>����[.��_qݕn�w_���5*�h��O���)qkx�پ��00���w�Yny�>*~��IS��A�jxXsU�޹�gUR_0�o�������ez���'T���
�]=`�ے_zLUo�
%g�u�~	��S��h��?���i8w+;�"���I��t�^�=a���0��+��di�oJ����^0�⋄��k���C^Cכ2��j}�B"���
+A�Z�',�T��6[�ٙA��aB���9��yQM������%<����iɺ�
��. ��-�͖��e?E	X�y�Oܱp�̆��ė6f>1�'b-쪈��F���_�sw�@���Y!�a��9��#6<���vLs�=�A�qF9�)�̭�+q5U�Př� -pc�8�'Eb�1��`��j�Ɣ>Y��H�ul-���QU2�a���ƽg�"�Z%��ɉ�Ib o���z���*��`5���1�Y��6FO$����X��>1-��EFv���.{��b+�� e:m?���o��q�R�cP�s�����م���;P�: I�#WB�&�1�t}'!����M�6����5� �N3��P�x�$�
�ͤ�P89�ch�5M3�͡����0!s'[��M�����6g۱!�%��+����i���pj�]���a/�~�$������̣�h��KR��V�i��/{�����Ѹ���L[�~ЯGtP���}�̺�9ǖG�<����i��27�
����	$������:�rTs2����R|�2/�<�Z����?��a,�G�������A��Rx����b(�i�j
f�����E�TWXZy�S�1u��;u���ͦ�%�i�I�IZV��L?�r�ؚ��dq��r���{H�jӒ�� S#CJuz�Dx��ZoIo���؃!t�+�.$oN���Q���0�rs��Cm�H�$˰����}�F�� IPJ�	�e��C��(GZ�\Eԩ�`5���ڎ��S&s0����ج|tF(� �ή[~bID�11�>�۫��·�&�WȔYs{":��`q�����6��-���^���xrHwP�[���|$9`:��z ���a�ߗ�.7�\��{��1v��%"�c y!A�-F^�L���'�jc����t�뙒����S.+rK�[�v��]`����mOҩ+� 0�9�Q/�B�3 ���s��$�x��IQ��K��гJa�ͯM����M���l\���ѝ�!�u��n��3_��Q��t/P���x�F�A��'_�|#Ufܟ~z�-��Ufa��1dC	[_�)&���Q|Q�<2L����,v�\(���YM����L�}�DGq��ڼ���mT��j$H>{�q4�6e���*��)�N��:9^��rYm��wS��z���'42p���t`�O(�2-�d���F5,�l��U&E#��M�N�Ǧ("��4O�M!��ÌeڭS���ZB�,�M�����[���b��kљ)�{���7Dߙ�plP�[��R�˫�J�Xŕ��7��2(A��[)U�(�A*��d�ta�$g�=✠X�ޫ�]��U��;;�D����g���-�P��^ޢ�7$Y���O>���S��BoVN�U��U*w�����ҽ�+�ZBx�-��3Kؓ�!����C@<I@�����D�!�i����_#�KLW�x�a�1��@K�t��e���.��4{�C"�WxT	Q?fF����j1��$�S�E3��ߢS��)�+yb��F������	y$�[+8��օ'[���0� �V�?�O�����$I�����gS�Ѕ
~�1w���]�������̽��`�Q��R��x���qs�� $�(|-{J�@/�vq��L2g]i��W��6/O"� Lڻ4��kh>�[�Ի���":�h���K_[�D������][��s%�����2�ΐ1�zM��1��s�<�P�ۄ��6�t6 JHz�<.�^fN��7�U���|�e����Tm���8Me ���7��g*���_˯���M�� ��5�
f�~%6go�2~�]�_���.<��[��9���>�۽D"��w���/WJ�>���s(�l(����{̙�c�y}�C����VP��c���y�2�z?t���5�켴�]8�,���������#�'��'��Efz:�/��D��Ȋ��R�M>�#��[tpB@HMr��\��G�����ġl�`���� �defùg�����q���J>6f�1)t�����e��	F|����|�J�v_�-�0$��Q+f�3���M�%�xPp���TF�:h�x���2�]-k�Q�<�t�b�$�^��e��f��>�nJ�Z4ϯ�L����U����师�0P���' ��m��Y��;1W��˼���()��!���Qe�.C�o@M����oz�Efʰ��H�;݌���Z��h��J�w#	a�N�<p�d\�����`*�T�V:�ɷ\�Aۉxc���k	��<hD�e����9�`�ӨGm��km��0������f:ݪ�\��u�鄶��6��C��5��o*�g�E������.��Y>��P�|y����0�V��혩-w�n%�S��f}��#���(��]|rK�=l;�EǍ��� �;�gk���ߑ���<"\-ۑjw�j���/X�7����$�yP`���:��2��>�͓��IsOT�J��g��HxRc����O��}���9I��QzE�J�U���Jw���-G8��o��{��G��x��sE�bz���2��k?�Q1lK���$ *��/���˙\�*2�B�2k-�^���ǭu!T��;�כ�)ԑ�ʬ��*�)4�퀮I���$����U��<�!��O]�A�m�F�*�.�2�Έ~i��[x��0X'��GxUAD�]�S��4�&�U�. Me!�Œ��a;�S=�zik�8R�dc�V�!I;�|��f��No���m:��hY�-�ề֪KR�-9�+a0"��-�_*�6��$��ҙ�4|om}���:KKۚ�"ȭlb}���ST��:oG�:w?���Π���(`��U�k�H
E�7c�=����9-���T#�<�!�&�J\R4���uj^�C��^�}mQ�%2�h6:1~z6�� �͝S��Z�0�)n�����4�r}��#}��Ə����ٺ�ǧ7�pt�Az�8��!��i�+��fm,g��{�Sl���R��9�m\;��܍cjfoGQ��,!���fQi�=�Ӕ�VdΫ���|cp�]��չQ"�>�tIA�cG	��3+�#���w�3ǒ�(^@;i�#�o$]5[P+fn�d��^DZ���Ƀ�"�g�i�95r+8L�p�W��F����M����Yj,!Y���`_)X����+�t���}#��� �sX�%#��J��;�E�U���LO9/%�d_:2�w���?��w?gfu`DH������B�?�v�̅��o��܋=|��R�s.�n�u�S�D�5�C�7�+C���o�=DҸ�^y1�UiT��Y�(���l��&�̪>��X�ș����;�c�^�Z����a��c	J.9G�Eb	O��4���S����~⠣��8�C�x�3n�MM��c�E� ���>�S�D�o��<H,J��,�^:�T�{������D��&�k�w����zɫ=�p�����k��i���^�9jxݜN��2��{��+m9�
���$�o�:XM�E���ƭ�$���l#vx���չ��:�CC�,�%��M�hGS��	�x���k���Ӑ]�A���<����ݬ��»C⃘���݊[T�����l��SO���\�9/�*�*>~j��4��$��"u�+r���~�<�կQsBu��(��A=���2���n���h~H��'�а$����(N��7�O���Gl��"���vga�3�\U��(��A?H ��6hE���+��Y]15jٶ�<��m�zm�h��I��D�H�i�+�S���/�f[��6_�v���Y��y��'��Nk+�#<�զi�dG�v�#HMԒ�+�G��'��b�Br����W�ҽP@�\D��e8�z����Rs���]��$�"'�����~��I�(����5��P��7��;!b�hA{��0�t�7 �S�-p���c���Q����>}P�?`���^���)#U�.��SG7GGOh"�����\]KN� �= �N���\O�/nG$���[1�'��[�W�_�*�.BO�x�8��Ё`��kH<�m�Yb�!��@�)ך`�����|[�N��B�+��騪M�u�ү.�U��hD>�`��5&�����CU1�F�0v�� c�?�k޽L��r��[��&��C̚����CZ<'�iX)vJZg��b�e
���}���W.q5<�Tv�}w�b<h�NV�)m���U���1����Q��}��n.~ke;�m�#��ԩzɘ0�7P�_�Uʞ=z��ũ��kщYQ�n�E�~�V�u���n�F��TX��[x�uNd�ʭqY�W�ߙ�G�Vi�g�nS,8o����"��3a��`|�A�3���.�ٙ�#��-7������Ŀ"H��{���,J.�]�'�A]p8�<��z���Ws�Η�-��5~�ى2�f+�ྡྷ̈��wV�4��R3JP��֤�M��%�b{�Q�:3XK�����9Hh�zv��0̓��� X��I���	����~O^���a��eU!R�يss�jBC��R/ t"�
.�@����C#�l�L��='Fҽ\t�'�[�߿����`ޝ�˜�E�d���yzfi6��G2�����Y[�W1	J�5�
=�_�a�_�b"�V��y��B�-}w�	��WwJ�;�9�~	�b��Q�X���ܸ�3aKJ[�N�Oa,���&��~L�W���͆�fh	*ˍI�<L�9�Z�Wڨ'��_�����|5Y�6g4�)��`�g,�nr�?�* 6��fLDÚ@0��IP��e�r\���EVZ����n�{w�^	��[cD�TU�o-�7�E��Z��9��,q�[��I�g�z��D ��tm 'YK�D-P�n�6#}�q��2Y�PYE��R�n䰧
��|9�p��G�S<qu����.fTٚ��{Χ[���E^%#��옞�޲b*^�1�}�5٥�e��TY�(�^
^��c��1�ű<NF,�M�e�S@r(���m����$��gg�G \1�����[�@��]�ꛨ��g78���o�W��~�lL~�o�}��p[�6N7��d���[$�9Õ�*cDC� ��&Ƙ��D�Ջ}���ɝ�!��9�G���R�&u@��}�i�nh$Z���2Ur[�4;T|�,�=�E�(%����S��d������ڥ?��v
��~aA�.rA{�U�K��_�xl��k=ϥ���'��ӳ���t����4ͱ��l�0@�Y!�1���%�w���1"N�����w����46��E&H�@���=rxq �:�랙?
5�h/���$���Pc�P��^eB�1c��?����T_Y*.�Fh�$?'�����/��d����6�MJ"+�}�
{����ʚk���Ef-s�Aы\���z�TJ���Fe�f�#rI�Lp^s��$�Z��]uP��.�*ߦ���^�F�V�x���=�KF��������x>-9�[��EX�16�����ݨ22z 9�χ�~���r�̀��^��ɡ���͢�,��!�z!��>���`
U�>,�m� �7z�F��<\���	�Jtl�|���%��h�߃���~J�cS)��#���k�	K�P�+���K$��Fw��6�8)䣯`�!J ��{�y�gM�rgC�x��^9�q.�yC[��\�pm��e=Z�݈0ⷒד�ݨ�m�����v��ܑ�T����Z�u�gF�$��YI�a�]��)!��d�S�K�Q�m�l{���T�u�,5T��8���IwZɡs�#����������Q���ʇ7nٺ�蚌�c7�d��7�������+**;����N��*@�S8�8|P=X�RV�uVջզ>O�������qs���Ȼ�Ao�f�St'D���KKoG�(k#�������?U��^�J�� ��+;��~gڐ�`l�&W�u�el_��hm����3��*���䃶<_�r��0�6�k�4�sRϥ�e�����h��5�J�c�v�"۩z}��Z}�~��+�|�\���?���^�s+~0�d�8�r�����цM]����Wm袅~��t0��ޅr��G���� H�y�P0��R�p�W�Q�b5M�.�0�)��,�B?���`�I��?��$'��=]������8X�:9a]��:�&�/�+��F菩E-�*��'�U"h�ϐ���W?����� 2#S��8[<[��=���}5�@K����`��p(^���Mք�����Gqw�.y�̶��t`yت�=����6*p�'�Q���+�>F�m�c��j���~M���Y�c���R��p��h�I�U���e�yn/�KF�U���d�cC�$�	�9���iѷ�)�����jD>w�4��<�7^qa5L�gf#�
`�ʾI(F���ՍyL��HQ%��~[�I�~'Z�h4�غ�]{��,�ؤ%����(�#Z�'{۠�+Zm�k��sw�Ğ�4��j�2�f���*3�~_Ӱ��<�/[�5��{.G���u�?����Rh�D�<�.�K�e��4�1*��=�4į+뽇�e#ף��#��'���H�X����v�9��[����d��jn��B��=��-b`�P�`w݅P���ӜgM^��X���9F�S;V@��+Ν��˩��/g�XM�X���B>M�r�͍{�^�?��V�#W5���\k���f��!��z���S1Ec�d(?bD��L�Z����gͷI���q��ĭ#�7�#��p��ĩpI�@Y`#KB���g����^���x����_�'Р\���F� kR�*nA�p3����d.K��R��h��(=�G&�ߎT�
�v���ֺ�(x�Z�Ƙ��ų(�9�⃒�\��X$�P�H�����(|��k��y��oh��)��tC����8�\�A���o"B�h7!�TP�m�����C*�'99;�Nc���-�k+���Q؄J���)�£r�ִ�NRa�~=x v�S�=8��4��vn�3e�f�dO�q���W�,�r,���B�w)�X�p_	Ѿ;���J�B*�'�a���F-��1Hj��K���A�P8�������!� r
����*x%V�_����%6��
�6���]A^��}Ⱦehd�t���˹���1���8��ۍ�î]J��BQ��
��eCSU��9�+�$�yl���b���4�0X�
w^�X�ER��'�!�,D�$�y6d�+�z�)*��=%�R9��M�-����S�=�7��)����d�_}-�1��Q�7{7S�Fl�'`.�6M�}���� �Y�Ӭg�c��j��Pxs�P�*�[bcU}Pb#��8A"�şD�a����D��b���y�PG����
�Q��|l�Yp�\��k(ԑ[m�e ��x�)��JnU�m&�#E��ַ�b�\!X�a����`��6�=lP呥C/ts��(�|���)Pݕ�S�,��&���K�h@�oS@6��1tf��Z�>�mp��bU�;�|O-*n�.{} �(���7�(@D7N�"��z��g�q���I���5��u�w�±*��k�l9�S�2�qb�m���;g�i�4ҋ����lt��8�(�������Y5���oSR:0��[�џh�m��*����ULx��g�ǣ HSGX9&i �#���P��!Q����:�ćq餰�C��bٲbE�i���sJ-nU�wP�:��f���AuM�w��-#�<Z��0�3�����4���`��J��$7���u/&��s�۷�|)��1��WGK��b���o���Pp- ����)lXc�)th�s8�@��&ٕ��0?�Vv;�n ��;~~ìzD}��n[��ӡ@;�Q_)b�8�R��hV��XՉ1�����@��{�������E1�nJ@c���e�8�I	�ƫ����bg"���oa�&���g�wC�n��y� ��>:C^r]F�N��$N��a�B�|"@oЌ�VPS+����uKt�|qD(7 y���%���(�F-�1�3R9�������R7ch�!�u戮�y�L�|�?��\&�L}v�~�I��|Hba����(2�ʉtάIP���$>��av���m�����b��0�px���١�Ob��fNn���'�y��AQ�0�W���?�x�Ǔ���� ^}�m��8���0�8�3��63�&r_�C�E��[K"G�͐�:�-�Bn�`�V��`L�XdAs�E�C�@�h�qZWjBĽ���f�oh�����椆2XG0`[������ Ӈ��)�9���Y�$�z���t+��1+�)�EI�1�QoWNI�������.I<������!�%:m���I9KU�sm��H����"R��ٖ�Z��EG���6wT^
����T�n����X����^IX�����Nt��$��h̽ͻ�U*�v������ka��IR�b�����Wco3C��g\,���L[d:��5������!c�n�N*E��It��,_|��gR�3��Ki!�'�ai������� ��<��?��d3~�YU��R3�n�yFF���f�X���A�OR�Awo��&gw{��:S�/uuFD��O���b��kd=0�k1=2�	,׎KiA����R'Y�r?Lk?������Ž_�Ax�uG'���XWI ���:��?H��pb��}�Ej���V��;�QЙ��>f����1��C���0����C=C_��A�Ͻ���Βĝ\���ܭ�A�~pi+����A�d���j�@_?8o :������c:�=vhg*c��iA��Xtv�Ֆ�gH<��4i��s����u�uh�Tώ=_i�qg��-L��!��i�(�\#j9-��9����`���������9=;�:�a"����	����%����\O�sf#�/=6J{/�D)'��n���$s�B||�ap�u�iRGF�M��'8&�&�sfug�:����L��#*�U��*k��J�M����A�/��_��(lś�ď<��e�h�H#��鵋?a������zs��j�0XOD��1� ��16X�>σ���9e���tQ>���{ћ�����p�l�����*�4��M�������K,ۛ�B�%.x�`ߋ/U|�>���p&����"谒��'�M ��*��K.�jP�wUAt�Mp.ڣ�_��=k�*I-���"-g�mM���hf�8w�K���������f�1�<�r�,J8!L
���X=��뀓�/�D̼�6G]�/�W� #�R<���#0�������`����)� =�������3i7��&�q'LI�	��=_���{��*#�y,���\�Pd��5���.�ڊ��`v�!� 8I؋���C��� `)k7�V�"�x .����\w�aOB`A����*C��=_�V>�C����-G��G+QQ�nYD�~���dR���>{�vS-��-�n�s9��T\�~�3V+V��^愈��9��$,A�U�0�I*�I����p.�p�΀N?I����$	4��SH�������]�sԌ����*�f�{3x�#ѪZ��E~λl�	6����Y��IG�����Ĭ��6_��q������|��D��r�Y��$��������o���(����c�9uz ��B�S=A�(� ���\����\R$,�z����j�<c�ޣ���8A}�&}ͺ���n+#��Ȣ(�F�jt)�z&�b`T{E�!<�-.lB��G]�r��_���}8�8�%�d+: �u�oj�!K%�*�y���1�����-d�\ߢBm�秼�9��h�m��b��E"i��;?7y^RvW���a5��br�~��쯚^)φ�Zv�n�Su�Lvaǧ��bN�]�Y����v=��%���V��A���7��#�l̽Ĉ�(7��NŞ>�qx�z�#�C�ڧ�T_Jm��UI2���U����yc?ԑZ���4�zFrZ�U��V���i��&��,�ߤ��|�I�W�=���˸����M/���dю�7Q�[������@#x�ie��o�:Tw������3^
\u;'��P�����eD>.P^����*��St�0���vOפ�b����-�%��+�������x��6=�+��Y��v�����!��XQJ�D�~���ZF`�����5O�7�L��?N��У������&�ڸ�;�K�lh�r�!_��P���.6��v-���(������l6�>�Y{���{|��;UTJj��CE[����^\;ף�/+O�/��.-���@ M����b4�,���Z)ҡ���Ei�&�/����%�\�(��;�f�{���E_��~�ȰB����O#z ��߆�v���3��|^A{q����C�`ڿM5���(��^T)��"�X��i"˳��Uv-Y����!9���ӻ���CY5�=���]���j�(��C�0�G<�zNJ� ��7S�V��g���>b�s�~��� �?׋Gs��r�AbRRPU�!��Ls��B��5���g�� Ǧ	/��h�!Y��J眗Y������)g+l�F��#��+j���W�a0x�Wb��Q��'<�1��XW�5�1���f%�(��(�}��Ǐ��`�j����bx_���̤�'���e�Α�j�E�]"��m�sҠ(D�����2gL~�NZ��p�<Ԡ��"Sv����>1��N�B8]g�����k���U�V�ܣWx3�	�)��
(;��o��f��i��[B��9�-!,�^Z��Ү��!LE�LM���.l�f��?�%*����u�7� ���P9����"�>�'l��c�����cN9�v��Y�͆�q9�w}�r��i�<B��BN����akk�d����Z��:�l�ИS�
�K����oo9�y/�^�,c�!����R�}Drn�^�G����E}t;�����,���dg߉¦��	���?ch�J��26@�_2��[p��f�3D�vLU�z)~��~'�'�V��;�_���@��g7�LHW�ytUB����R���O���U��mU-���K2Mh�E���_.���}��E�6E�ho�Ul)��HD��*��sݗ�ǖ�t)P�D�f�*��&�
y#7!Q�f�뇖-�2���凿����|GiCD�PM�"G��[���Y�on�i��	�/�&�.�
w�6��Nm0�5��ns�0bea��e��6d�(�	��y�n�g`��3k�U��y�)��_�(��#��p���{���sh��6>�����'��<�?��;��o�;8�oT�P?ET���Z�k�]�y�\��e�f��:��]�E+�C�w1z(��	��K��7���Z�[b1�и�@~�<3�Y�\-*���D�ct��Cv�S�>&�%2�`8U���3<�'zP^zh�zy�H|�P�*g�V��4f�ڽg�`����^�
�=�Ȑ���C���򍻰�t��c͛&줧܀<�Vvʋ�U�6e�"FV>���c���fl����0� ��2���s5q���A2?(���w,�le�B���q3N&�Ŋ��p࠯]D;*"P�
�/��%G������ؙɃ�����f�K���SQ���· 6)I�r���?z�C9�ڥPP��h�o�	����a��F%>έi���A����u�`��D�¬���F�=�I@�_��mx�؆�b��f���:��G����#�55��!H����-z?�hƴ�A�wU'|�QM�+���B��e��=� zEɌ��H4-Q�k�Pd���ƱI$��;��4��Cs��!.�#�����P����5Gs��3Y��0ȞΌ�;:��6��h�r?�MI�It�q�ڸ�C[�e���z=ޭ��W\�ư���� �>���!�bjH`�å���ZeS�xl������9��'��Xĸs��5d"�ĭgG-�w��r�C챜5��2~S�m���BUo�����q����F[�`CQ6u��"�,Q�CU~uU��.S���/:Z�c~]_򾫥C�$<��\�����H�)���R��L���0�4}v]���s���l>��L�@����Wܔ�tʙ]�ʱמ��
���������pv6u�zM�1J���Z�5��!��( �,�3��	?%�]�~��pZ� j��Ծk���<�s*��Vu�>-����r��je�F�\*�w"���x�B�����(�{��z�8�����U�fmSP<h�q�)�B�%��B�8�P¯ ��Ўu�&ąG:��Ss{�C�J3����S%c�ko�8���=��\yG�YK�?تC6���x���aRc0�**��9�7�'��b�]�W�������Xq�������BHgh�Q4����3
�v�����h�2��ҳH�: �b#Um|_��j��"9:2p��<�e��� X�Ǧ(f�x��X�!v��#������P4�'b���z����;VP��F�j�y�Y��<�)����AL.���H��z��Um��@A���,ge��d̉ѐXh���06�j���l��V_��)�{�2���u�Vl؂���8��� �|�����@1h�ᬁ���ƠnhbY��䢪Q��0�P���K]��-��Du���'2��3b[�g�`�T�a�O-��)�c[��� #�8Re��À�SJ�f�a�eo���@�Rk��~���?߻���T�.>a&S�O�<{W	J��ظp����L����F�iE�镲�xJ�q�Y>%�ͅ|5G��m�L��8ܴN�Ȯ�ꔗ$w�!
+\Hxݦ{o�my���s}��Ĵ��󂆾r�=7�����i�i�WZ�kr�)���7׌(��}�K�e�dl�V��>�,��0�t-����k��Ȍ��U����{����*Z��E���({���������-n�fݶ��L[��2ܿpX�����1K��t��c�Pp�b7ґ��D3X�C����
ȩMd�8/W�ʴlYpJ5ɣX��P^Ｘ���F�G�w�����cQ��y?����*�M��2P �$���5U��\���b���Ԅ��(��9<��T
���t��z(R�)\p
Ba��:�p���͊�Y5��&2��X�'kn�=�T� %6%!̡��p��@��]�9�Пԗ�7`����H�?a9r���u��.{f}D�0�>3��ٕj��[�[���Q��ƈ��j�/��S�*Ȭճ��#?�Wf��\��M�rK�©�HT��d�vl��qb"��� 8��kY�V�3���wr�'��֣���=|�����
��#��2cy-��r�S�3
���a$��T���y�*�h"m�d6Qm�|R�"Y2tm!o�e���(vM��o}�X�"��p��"�3�[�`YPtf<W"�.�����ф|r�u)�ϗ��C�]�Aq��Ҩy�囥xF��NS�8d�>i	�E�8���=�	n�,]*K�م��F��F�b��3�!��	�$5=�E��2M�
���RG��PA7�2^�z��$���E�R��%�ñ��Bu}�]	�C�29�<�T:��d���@_��[�v�Y����d)�u[[�����7s���O0X�v_���Ů�w�aS�|���R���bTrsY*��p�+�LQ�m��X�	a��x,�˰/���ꛮEϺ�n
�Csj�JV�9�6׉(���*�ݧK��с>��4޴Y��v�1��z�m��XfU�������A�h�-����a���K���q�D^�J�g�W]>P�C��LV��%���Qlֳ\��ZKK��'7����+�L囖�T�*2����g晰v)������L�,х{G�}84�o~�D;�&.��t�X����Զ������I���q��j�.�n��W��c����Y�c^���l�b�.�q�eɖ���3�_�꥿F
B�BB����ɮ*��6I�;P.&GqCO2��nM�+�Ep%�s����p��� ѯm5��=��_��J��'AS)L)=�|>\rhX����d��u�^��
b���w�i(�lG)���p'�K>�
1�I�zD�í���ƅN^�i��tH�!l���\a�D�|CO��)�l����Y�`>��~�����W�.�?��:þ!�W��3�C\�Y��Y��p��6���;��0��)�? R��'z���jg�Cl�Y�\޺3 ��J2�ls[�m%N%k���I�Q$'i�N&} ��7süs�p�b�bS��L�ޡ��Y�6��:.d[�۠(�@�k���W�L[*Ti��z����c���Fҳ?~}����Hb�k�-�E���Af�R?��z!�a�{Ǜ��K׹�aj(M�;%���Z�$�-��Y�G�&޼�@�%7,�S0�>���/��������%� z��	�4����)��{��a���ϧ�iZ�!�w��>�z�dM��eS߱ww���yBNc��:]���Sx�PyO�^?>Yr�?�t�[�S���YϘ"��KkC�g����(,���9r�v%��jj)��,�_�`�ִ�ˆ��ϙ�5XR�CtP��Ŕ��5�@]q2(� V�\q,r�ӆ�!���h�Y�"S������NXﴇ-�����Y��Q���&�n�w��nC	���m�6M7MoT���7¥��o*~�=��/��\�r@�.̿YV�1����fo����-��߅���`~���������ci���T@ľ���l3�I����f�=��(�W% ����<b�-�2w<�a��D��9��W�/�c=(������x�8P����k�`A6G~w!X���+��VQ$v_����h�ſBl4O�#�Ʀ
�{Ws�R�F�*[E�Y'\˵�Mx��N?�S��J(yҸ��_d�/*�u��V��C)Dm͸�n�@6Vu�R�$�b<aכV���Q
��_u�:dŵ{gL���g��O���V�!XMFu�b��k��kֶ���("�%�B�t���q!;hǁ2Q�C� ��* ����u�H�ߜ���6x��E���"̠3
R2��'[��'�/��\��]��˲���O'\��)$<�FĴJ+��.Bt@M�6��ﱌ��y�z��)3{�;X8�������}T��s[��I�V����{掹�d��Q���;�o�}W�_�{5|�a)�G����I�i �:�b?���ۖ^��E}�*��|��gW�: ���������nA����}����#ۯ���p5s�i�2v%�'�T�61��k@�J"�ŏD�
+x�6vF�Ʀ�̋�����Nn�xP5p�e�����mǨ�X��Qs	�֥�B������.ȴ�s�5�����ij����Cf�%���..@Ib� ��_�4��6����x�s��Q�n���[/P����/������/�6�f��妱Ө���f���ՒE�����\��SsD��ok�E�����7��Z҄}�3ի&��%�,���ɫX�:7�2���ʆ��_W�|��b�u��}���=��BP$gcn��M�y��Ȼ~�4�byǃo�XE��C�2s��Y�������
�#�</| �M��: �YJ�f`y:)�a��z
}
�yb�&+Y0g�y�&}��v���'�"���EO���5R�����c
������S4,=Z�k�aE=bx���I����h�S�1���K�T)Ӯ���G�ڥɢ.]Y�ǟ�.��\�<�)s�hmU�$d��E�����HR�QA��~�#wv�>5(�L(���Ř��&"\
2DTh��N�%�s�S��0��?�G%�ԥ̥ޝp���/��6�By��5k�(AV�ǥ���h�T�`ޖ�[y
3]g���/ւ���,M7���x��nn�P���e��b�pl�O�Q�́v��.�>�:��V�0�-�|y�)a��`R�/|`�S��m��K%���!87�>�|�ZĴ�� �:fd�mLa#-y�c·[^}uq�пUǪ,�Pb��Ӣ���Q�=���U}W�7 8�Z�\�B��k��M����c�(��L���%-jlF�\�M����O���oiە�ūr�qG(��ów�X�G���%���	u��/Kܝ��jWl���h�\0�/Z�Xf��毪�'U� �� d捏��^f,��ԇQ�m�r-�]�m����.��#��	����9F��[�K��p��PQ'���SL�E���3������Iͦ��?�M�V�5LlFF���� �\Wh�1�	�&r{2�����|���Y�r�v�/�K��>�/]���E���ɿa�h�?��se	��P���d7��Ey�U#e_6*qP���4��y\r9�p���RkIX�^���D|Aڨ �Cz�ts�L�N9Vnbvm��U��:SoB����NGN{����"��D?RmI� 2� @���=PP�w����L.�c��D��C�@��S�5��(��Y	���I7'��̅��+�X�����ˌ$�h�6��8%��Q? �^�Z�z$�%�М��Zn]�P���s+F���^��F"5��7;���>T��񌇐G�`�Ċ��-s���4>;�sB���r.m}t�=%����Em��J��'��!��475����
"�S/�������8��
�Oa�Ǡ��8�m���*��H�4��x��5d8眔���K�Ca��,���J��\꣢���7�=B�X��[�灩��WN��t�B���w�.�"5��M��vXNM����ܡ�4�.���|�&V��0�3�R�4�v����Jw�ٛ���O[˟r#h)ʵ�dp��_�oFp32�FEQ���L��T�m��@��0�hh?-��ǎ� ǌ`+�8�=*�䟣:B�1	t��o����l�����I�X
���}u~�w��N��B o���YI?+�d��1���=�"��������p�UNq�<���}q�4C~���~�L{�>v�p䄊�3�EJ;�]�p�eo���9�^  X�ᦘ1F�����L�]s� ��b����8rQܢ�~iY�g�8�%�̱�Ǩ��)�὎�h׶w=�4a�i"�nLw�8�s�]py˛ˠ��e���t�:ƚԬ*M�J�����˕�3��r��t�Z2��g�N�9$qӺo�q�ʣ�hgK��q��5BJN��H<�ƺ��%5����a?S�u%=@��8�â�O�w}6�Ϲ2�ݹ�8�v\�Bm{ކ[�����UAcohK��0[%���OFe�(t�,!U�����DM�:�����h����:#�Hۘ��t
�$�KL�U4�'�Qr2���;�Ҙ��ܲW�<TW�o�U���J�8�j/eRm���ʚ�*��CN4�x&]&�f�n��*���Z�v����!ut;L��Zo!Pgcr�P�bZ=#iЫ�E}�I���t͚f��E���&����;��E.������1��|�1E^��樽[���K�LSa�^?��N<��()�E#��z6؀и?��z��g���5���;^1AZ��T�'(��	5�]�n_w�EǷv�O�t��^��M����#ʹ�7@���m��H�Nߍ=К�^�ő� ������ä���X�����n8U�k���^d������6X�e;Ց�dM�e�����֊9\��ނ��+��͗���$��pB����MKs��	~���UB�b��25��ԵℏX�l=���k5|�&)�Z�?�����p��~Z�� n>O�7��?�*��z�t�����(��Z�p�WѼ��L��@ь�����q�q�����+��ב1G��g;f���'����O��+Γi����p���]Zp����GHBdqب��O��-��H��?��B �ϻŶ�u��eؤ�"��FL�� ��$�^�)�[�F���<���;�����J�x�*2o�Ȼ�t�|bX�ح��
Ng���Cf�m���^�3�UOƂ�{,{_�H�^.�%Z�9}�.kj�#�<B<����p��	��9;tg��Uv$��2�F걡��`�G6h���gQ�w��%z��8�0�G�G�ʰ&Z�\#��i�S�24-ENRki>�_G ?r"FίN��SX��k+q�[2IW��ԗƫ[�Nvg��B��1�3���PO"�)�ĉ��-*k��m�󴞒t����A�<��rb�����'&�u{�~M��2���	c,KE}�o�� ������>ι�Tr�?�i��9�)�嶏�D>������z���מ���t��=�����kS�z���tZ��7�"�w�WMtR���,ϧ)����v6��͓ [�(���d5ZW�S��i����Bk`{��d5�����4������(.!5A��Hbp�مr��������=;���F���4],�Ӊ���.����('�ٌú�=���U�Ek�O<�k�68N��{�zcTD�PY��2�'C46:hW�<�0l�rM��+#qC��Ntm@�A������ƙ��"�e����MC�cŞ���rY3�hHZ����P���z¾o<p@v��gY��!
D�d�"�g�!v7FHp��BJK��2R��~���v���ԍ�1��Q��[E}O��P��ͶP�˦�e�>�A�j�Hu��(��Fr:�,l���W��X�-��-��==�a���e�1"��N6/�K��"'c�eek���AE5'�ځn�!#M�$^D��x[��L�����0��bi�jM��ᢦ���l{.`(@���X!"�Lr��s�=A��͊�!������"����b��&�S�m�����֪���7��B��tq��Y�:�dGWq� �^�#nF�w��+ߴP�+-�>hSl�cAG����ʝ��&%ʍH��B<��bV�΀,�XvG39��4R��C�l��.��bӂ�~\n`��J!Db{�0mj,`F趣u,%�&�E�0�fAG�T��ߓ�х�> ǸD���<-�p�"p�d�����:�=��`���k�6N�����}���6�hW��ݜ�i����۰��$v+e�|>�#��U��f���s��8x���@2�����d�
��V� ��')|�ηqV}Fa�Ab ��s��@���Q��pZ%�mV=&�m,a��AC��ą�m�����d��ߔ:�S��Q.f%��z8g�3�j� <i����W�V��p��$߻4u�w��P0Cxu㽣9Tb�Ħ2�_/)XFsa�\/����%���y��u!��@;m:l�^��0J|�
��� 7:�¼�B�!��߯������$� #�}>�j�4�3��~�ы#�x'd| ��� ��YX��
{�l�5��*���i�N:H��wM�1�:^!�j��Wo/�*u��X�

�$%G%IW��tvr�	C�+T�Na~��v��N�>��'�uPbױ�%�g{V�i�jru(<�P�D��d�`q'�?��]���t9�i�!=4tk��]L.����R�!�����n'Z���&ƿJs�4�H)�K[��)y�Q6�zkW'��U8!�k�����	��m��m�,��� yFN!�0��4*3���'��� �^�Ŧ�*��8cLg��*�h34502�0�f�D���@j}�����&��ن�}I�O���[�d;�N���:���� [q��t��1��;��g�XF	c:�|˛qoJ�p@��Y�Ck�[��(m[�,����o�N��5H�މ����J5��o{��[��]Z�d�y���n	~"w��:	�7 �gL��y"�����]�?�Pt�G�������[�ϳ���ԂZk�[�#OLwU��[�#'(�]Ov��@~c�����
��{�C�a�/�2�v>M⦺��^�-��E{4Dū��Oym�0>{���<(+y��+u��G�xG�H_�F9���=U�A}����=u�
R�?�!�t]��@B����O�뤜`�`�3�|_�4��Y�~C��F79�+�#����g����o�[��z�s��9Nۀ�K�&0ydȈ��7�Q.�YS5�i�;�WX�
��H���I(�����L!#��K�U�*x/�W�&���n��`RBP�2c���ԕ�x��E�\�AoG��,�E�z;�8�B��=��B�b2�WY
�EB�-�;kb|N�=��>�M켆D��>>4&�[�uL��;�R� 5/���(yᡳ��U�s����ڇ�g9��y�I���G]����63�����{P�!F�����E6ѯ���MZ%���W���ڽͻ'd��U)��H��b2Vׯ�����.��-�7�:�"���|&��������]��ʭm�п�M��\r�a[&�G��y�B*8P�Ð�]�$=G����>8�M����O�{D#�8�'"5�P�)d�R�c�����f�$��7�i����b'���0�2�ttb&���N���}��ʹ�l�ϫYܢ�`�m�ں]k���|�W��,]�7j�xw���X�Y���/{��E���^d )283d�|>���#sQ��Zά|Q���I�b���xae���~�@�������#����,E��د���h`_����0I��k���Z5Ĥ�����˻*���cy�a�n�X��D.ӆȐ	H�6���'�p��uA�D �	 cRlsl-"W�Ô�,u�O�(�;šޟU.	�/�WC�Aݰ�1���Ցav����� -����8�~���A2d3��S]hD�a��{��s�s��ῢ]g{Rm������~i~��z���0>�E���琿G�`
;}�~^.#�!1U51��x
��i���V7�N�Pz���8ض��0������s_�)��:|�K;HC�W�v1�Q�2?�qmv�͛ˋ���Ð����s��F�����'钇������g�J�C�T���n��(`�؍�Y���Zy���ǭ)��z�����I���>P�vt��r@Æ�|?Z��-7��9t{(��\��L9(Z�������׼[�[I�Pn|o2YB�db��r|M����j��t�͕��������1(�U�I�i�u����9B��w���S��9�?���i��V�������i�]��i�H��ms|D��z�#�u��;��{E���ȩ���)�˓LLT�
"IúKc�9���1�z�L�]_����������u-��*��?U�Ň
��q%���!Ob~Aځ�Xf'�����@s�k}�X��w�U�'�(��h����^��z�H+p��}�낗����wngr���p�M���I�ho3Ba��%=,���������&*��ն'�|BHȢdzpó(���#nv�Uk�m�����	���%r]B=a5g���B�|-���p�Mn����������yZ�LL�r���׭u�C�CZɖ���P�C� 1[@����[-�e2��B����_����2H���� #G:2sͤaX���2A�*w������dq�\���,����)Z�~�D[�jm܊��_�,/̩��<l`�1��Ox�E_iсT(N��5|�5cx�v�c�ОTB�9�� bxR%d�����V�R$2��o��oo�3M#��dl�gǑ�KP�����DkY(�������R����ʔ�Y4X|�4�nYV�e�H�ù�����-���r��Lk�K
S�⧼�ʌy��}��t�}L���L!�gF�+V���2�H?IG�,ཫa���쒚��"	]1}�>�O���E����ǀ�^e����uh�Ƶ��ʣ7��7���1����%+[7�lJ��Ui��%��F��\���Z���e���xA�89B�!!�\J�fk���|��#N���~^Γw�T������4N ��TBܣ'4�%�D���x<�P��+����\*� ���`K)y�=�U�m�����`7g�g�o,���7
㢞�l��n��RP�G�[�$�EwqTa��M������M�Xb�"��bq����,9���+�hQ��I` 2�XtiK~A�(l4}n�1���+"R�Z�#v���/;T�*�&�O��HI��#�y?���*��QY��TmN�d]�{Z%�����xl���> �i���vl��M+!�|Wjd�|���	�s�����"�#�en␇�
�����
�}J���, �S����:��)B}ƴm3������6!H�&����ex9�G���8�U������,�6@��;4%L�x��Vxk�V���QX���4f[L�{O��N��9	�q�����YlF4�uR��B_QT<alg���8���f:�Qu��h2`�5ŭ�L� ����*�,� =<t,~�t-�
����{M��9>Rh�dv��`��l�((8q
�x�M�7��p1a�rZ�kK]uR�������L��޷L`�yO�uy�9 p6��g�b�߃����c_�k� �Y��-�rǻW���ÏKץ�Sm?�B���cE������LJ�r;��F����0ܺ��@�Iz�<�l������yxQ:L:�vb���F� �v����G�w�UX�T3�	��Wi�S��A��ċ�a�X��7����[�O��r_����PJ@� �Ǚ5媪�!�"�����r�kN�~�	C{�����v3����������G��Б'8Q�0��ȍ]֔&�Kb�!�H����>i�[�	]ᬲN�[<,�J�\����:Z����i8��_I�������)Y�2iV{FS|Z��^�o��j���Ɇ?��X���3���Y�:A�y>����.�}���`6�q$C���v#Ԋ��8H4I��L�21�/�*褓ّ��1�	��_g�\4�f��s�v0���lZ16OoMy"�:�3i�>r�<6�;�K=&�-�t����_�+�TF��20�,;6�VΆ���^�+�W(&Φc,ܐZ���#7&꿸�jG�Ԩ�G#�z����~������a���s:oK���� {m�w�7���3Ԁ�O�N�l��~�$nN�q�L�0;Rw���}~�1G�����oF�`U��)d�����w@T܄>���ЌdA"'��~#�2+Q�d�P�S(��e��5��^�*��:%'a0ϼ����#]��aˋ-l��z����q뭩�k��N���0�i|�W���G ���Ɂ��F�\��"�/��N�B	_Ǔ�Fw@yqk4)�@�V�u&�[*��^�@�i����_���D�}�|�+ g�F�?�'��V�4h~ 5W5��nu2�>���Ń�:1_�l��F5]�*wKʝ�	{�BR�C�X��zml�=�fڣ�����g�x�T��&�[-]�i<�]�W�q�1ΰ�����-���������&�$�V�L��\�����!¥b6~?��C���6��q�2z?`A2�}'ɍ�]D'/`i��c%�E�����K��7OU�-��e���(��54H�v�s�ہ�*c�#��J�[�{. 3<5�"UȔ(�^�R���*�R�8,�96c�.��d]�6f��MT3a�Q���Dh�)L�K�$n�g�n珣��w{��'7?�h�2/^�-�.|�5�=�C@�_�)��俿�nV���^�U:̭�gy���V�D1F�}�1�b�M��ڬo�Z��+N�7T�%�d8�h����[����Jp�2ݪq^4�DG*
$�<�n���IY�?��Aj�e�H�`:�"R�K6E�ϙ�X��o:o=�[���J��}�:Θ�ރ�58,,F-sԽ�Nc��5��LW�}q��Y0������/��"f֠��Z\ܯ�S��1��e��|����{�C�VZ9_���q�����*�GM!%��Ϙ�t�]�19M���A��
Ͷ�)����6T�k���#��W[f$ˤh�����ys��u�U �aw���Vp�ԛ���tKy�l��ˍ��$���0�@�5\ӘG5p��U��:���=0�A&م�� D�YyB �_��&cf>�Z�R�ys�e�qUh��e��ݫ�q�
��'�����>�H�j	�풍PM^�i&�4�����D!i���#�'�Y4])�d�=bjbĿ��D�_�';��1l����Z"lty
� z)��}�ۡU�BU��}�3%�gGWC�ă �X���y���A����ak�����f��9(I8u�|�D��O٠Pz�U�n��bN%Kg�eƹM��(r*M�����F<	���]�)��D�!��[��#�*����$B�t���7P�KH]���Z�=p|��b&��$kfC������W��RE��<E�Q����`��a����,��$ޝ����$�<�sD�pٍ_By4B�!�k	���;���Դe^�D}:cZ�d���ސQ�M٧��?��6�{"� �j|�)�j=i��#����@�J��A;@�u�b�T��)��C�7�Ng�[��K��T ��<7���	iGV����Q_��7�W�6W�]3V��@�t���=�\�M��7ij�zΊ�4Hd�? �4<#q}�L�N���_�ػ��SBX�E���0���O@	9Q��]x�$ot�:ް��#^"VP=���Z��':�C˝�#�� ���@וV��Æ#(4g��N�L���:�����%���p'o{y�Cz��x!�E�s��.�c
"�d���Z|b8D��u�����n��Ys��х����kg�Zf��P���;��Gc^Mw���|�^�����@���nSſ����b�J+��|�MN �����ڨ�q�.����G�gr���6��㒇�i���O��Noɳ[+9���xDn>̃�:�tz��������@��/� ����{�7<'۫c~L"��^;@WʰN�A�ʉY�۝��C��5�5u`�%$l�Β� F-�_y9���u�]�����~x���s6��N
�M�C�a�~��{��?�d�|cR&+�碑z����$b���?���L�8\�p�ү�"��?�\sW��,��g<�X_1���l��-v�&S��mB��g9Z��&*�T<I/I=��.~,��#��J�|��@��!�NᏃ�	$m�P��[�vF��ӚYC��� 0���7z��0��8(����rHCj�Ew7[2T��~:�a��jI8M�q�D	��r�РE30�#}'[޸]��g	r��"j��r�JH��{?r!�<�]�r��E0{#���]j��5'�+���	۪�����6:z(���
��
h�*^h��N��ȅr���n�N\m�ד� Հ}�d?%4x3�n|��TtΙ$Li��p�舽W�]��{h3���r�@�ۡ3�l"���9����mؘ.�օ��*V�^������3�A�?k�'<�u�Bs���'�C'���e3�����)8��\��H+Y_t�ί~�EG���=�3�jxa��L	zك��e�����꼲��e�ܔSa؆�%��R	چ�[�F}p>��02�}u,��錺-Xݹ�٫
��=s��W*PW?���Ɂ�Ia^'�¨��i�)�O�J5�!��9��o��� }D2BE������ذ����k�����CJ��˷Z4�*�u2�@�ǐ�M�p��xa��QK�+bfHw��Q�DQ�M͋뼭D��.������n��C/.�y^���@�\�7��>1�K5 ����kH�)J�px*�����!O�]��b��ZpT��4W��k�!M��ۀBjI���F1�##�����`�{"�v*�	��SM"��f�qF+�	(�4`_�I9�og��jm��4W �ZʱϿ4���M���-n�:���]�V.�f�0�TrF�p��]z�+�r��:ړ��K�
&�'9�\2�h�� ����߁�D�P�K=tu9:r7�.�oЂr� �y�r��Pq��(տ�a.*�B��� }Qs��a���pR۾<� ��j�[���*��@�%�=@��h	����u���,�jr�7@�i(�B�V^GZg�w+<��\eF��U���z���~k�dzs���q��Uڛ=_8��ԡ���bX��Y_�]rOTsT�,J	�u9{[wy2:"�=���(}:Q�ν��3c�`��&��l8�c�����M�11.���83L?�h�7��k��xr 7pa�kC���q'��4h���^u?ml�g{پ��nP5 x�(u�(��mZ�I�>t���&_������Y29,�"%���6`7�>��Y͹�� �M	�P2� Zڪ��ڥ|��������`�k�
�ҕ��{lCy���Hܚ%3�N5N����D�#9^�#�f���o�5���J�L�}M���@��10D���_����:=5ضl�%�N��$�rd�hk���MLpOZ�|����?6 f4t�!���QQv2����eP٥�
�܎P
���1Nʯ���O��b�=n�~~�p�=.�a�@��|8T���a���2�a��Rm�%#���B��;_�\d������*�-����	9��~F�ԛ?k��uAEl��@4�yn@�`���P�b��� U�iVfлS�[~.r&<'�E��w���\��Rh"NP�M�0��SxϺu�y�S����'k�&aA��:�dG{&5tq��Z7�S��o��tڮ9����v�:����t'��N�,^���j���R�/6�b6��+��p�C�!і�����CP�� �;#���r��"f=8�I��n�����$n9�[�+1���\���2Ae�8pWȦ�B����7�O���?w��9�N���t��������vP���W��*J���MkM@�s$M��6f ��
�n��J��fr#�a	��������{]:��.����^�	 ��Q������u��n'�l�"4n�.�9	Y�l^�o;� �w	ǜk�E�1�X|�c44`�vL�GP:����4PF���7��Ž��Ɩ�C\��h��E���Ou[��קL�L�g�?tk�����Р\f��5Jc�?\���B4����V`fWH���]o9�ŀ�F�ɻ�W,p$����b)&��Ԭ/����NE���#75�J�NZ�ܼ�}�m��U�� �d�W�=T���hq��E>$b����'�'3-+ҳ�Ə�7�.N�+e�I<�����n��X�5u�������F�.c�K��oח�8�����؇�B���}ȗ�X#8��n��Cu�
�4�ۘ�/[+k�]x���l�#�6�ӑ]%����(�砪l�|�(�v�@�9I��LfjR�`>��y��L	/�q�x)m{B���kv���!�y_#�.��@��֚4ٌge,�Pܹ�%S�M�������?���&R�.`rj��m�o�8M�Lk.�q��QC!��'�$?q_a�������'�\]Bwgp��C����vh�^�&�u�-pY�<r�R�z<�R7���^ ٷw��APoo ۙ�Er�մ�vHh*��'4Nbīp�w_�)�O
�9X�H�*z���X��J�Hf��,������0bL�0����7�!7���m7N��m����%+?����Z��lX���_���U%zK�h��6���2�\V=<?1$�XV��;+M��?�4�Jũ��������q�@iu ��h�ƅP�M#�1�L�<����9��C�G!H��5mT��	�����(!��.r������v�F���!ܼi�w朋m o�Lgw��ჀF����p3� N=dI籠��2��W���������/S�K���A�à~�/
~���|4$?����R]/=b]��,X���j0�F�mCQ�.��@����6�"��JC��t�H���g���48����S�����s~�l�+ժ��8ӸM@�lԞTŽX�g`��XV��x�`y���cz��C�<����@:�T���D!��!��]/�=���C����пN�R�����&j}���0�y*�$׫�[�L�$�m(! �7�:D����,�n�2�� 	Y��[y�3��䩷��zz�*?�M�����T�gq�<x�8q�F{,
.�#4�AvgtV�U�g�o)��0%����߉R2�I�:a̔�;q��Lﭣ�x�����){Af��c�nZݘ3��5}�#/3&<6N)NSQ��������8��r���b�=��p݈�s����%��3�+|L��?i'� o^0S��ڵsN:f���3�S��1�z�����L�O5|��׬�X.=�vH�`8��k(���<i`Q���� �0!�4�:pvy �ھ;��v���.G�|$�)�Q��&�A�<����!�gZw3�#��fju�'1�����(���R�I ,m�nUb�B�p���Ƿ]�����X���T�1���PU�Kv6`���H,��m"���ĳ0!Db��d�G�a�\��� ~�������H*Z~�g�܄�|p�+g�Ї��v(O��[Z����H�$Q�h�bo�C��=$p����C���V^���+�v��.���ãk�ؽ*�%V��ctP2:s��B΀X�D�{5X�U.8�V��`Q:lT���� FҙIJ��aL����>G^B�H�O4�X0<~G�ؠ1��Vm^[Ͻ�@�,�s�]mG�v𻵓��c;��#e&~G.#99�P���d�����'B��Ux��00C�<f	"]e�GHL��l,�c�$!}t�1tS�B�=ifع���-4I���:��Ga_)<���Ӻ4����K/2
�Ly��1�ti�`��QP37=�0ӿwI��j��
�F2=������R�r���$(���W��L�ތ(����| +�2���	�����~u#,<�	�!<��z�+�����BH���sX�.�:��鮗��>ԴOՉ��j2b<I��!u��N$�Þ�')iKpN����eȉ:���{��EΚ;e$��oD�PF�zk�ᨒ��0a���Ix51ձ~�r�5h���VE"��kt�1���(z�-|5������_<��A�P���H-#�R	����Û�+�O [����Sh�!����<h̫�{�ˏl=��ƭ-9~i`Plw�}d��*fuŋ]<��[��:�3�C���Rw�;����QI�U�L�H�Got�%չ��=��?^�J�9x������/�p�n\X�8�qWvF:�o�A1]�Vp�����a_�n���7�hAa�F�e�2ZR�a溓��������0(,D�eĕ�{*�[p��wΕc�����&�@%�<&N�*GS����s���.�-�R���B[��L��gys
���� r%�7��V�.�ex%��ߡ��#�%TS����6���4[hT�e�eѢIM�"��Myc��*��lJ���-��{�
%���u*�=_؊*N�Kɲ�Um������7")-��ڒ=�y�#�W����U������zο�ez�t`��d��X��O����������P�o�B&�� ސA��,����f��uy��bM���k����h4�`#���k�L��$
?���i �U�b�`U[��ou�?�2�$��B�U���ېhpf~$�!�%KY��OE��s�}�N��*�&0a�*���z����@lٰ��GdHv�@,Di���<���aM�%��i����F_>H �h�|EH��0�~2/n������:j��+��WGM���3�LT��_OO:@��}6���:q���>]_|\���?_S$�a�)8j(�|�Ӈ�/�*n���J3L�d�Bmi�OL�G�R�@�ƕ��7ಔ��$�'�1������#K6�%|�F0��t}�RE o�N?�4 ��ԙP�%K�B-\�
��y���9�d������T�<�ji������E�s�v;�����ki�Sn�7D<�
#bwE=�VD��y����)�X3H��Z�&�e�-�H:��)E�c���W����h�YՉ8�d�4��/��s0߄P�:�D�U����40��ϗ<Z��Lcq����p�����&��q��d�b�/�`�)�6S(������ą����*�F'-�Ԓ�ȓ�+}�贍c�?�	�r�%h�>�'؈'�
�*�B>5m���u��l1%��~��C�ce�h�KNDm�<o#�H#|��E��K7�T,|�zv}��}�v�����l�R��o��Lt��	����w�k�9���>�R۸�p�ڲ(Ơ�1+o�U��l�P��3�؍��r��\�.�1p7��"��{8hԏ�b�ݝ5%�i��:��T�PL�0LQ)�7�A���.n�;SA���S�pC䫯��[��{8��	��<:@"��O��e��#��=#����)�l�u�	�����GնdBaKhgɘԥ�nÚ,��?m��VӁ�������r�}����j��J�^�A@��ޖ�Ж!�j[���q��AZ��μ�%�-/j�����&�����D[�@�����G�g3a�.�+��c�1�s��v���������0cG����E�@�Ʃ��Vb���0"5b��$ (����QfT��W�W "ߔ��ő��ʎL�	�UQ ��JR��%=�!A(4����Nu�T5dN�!����B�F���V\w�m�� �\S�ŁW�~T���&3��1&�#��6K��U�H\�F�C�P�*�}𶰩��Awα� �����c�%U-]��w� �Ut��w+T|�V;e�{�� ~���2y$���N؀R��.�z�\��Z��|`�E�w;�A�z7)�M�<I;6�n�䢨�ڷV��0f����Rj�\a1�H|9w!Ѓ�����(���;$��dd�9���"9k-��O͢�irI7Z�M�K����SUc�!s�Q�`G\a`�u��v��ʀH�ǤЭU"���Qp)�m���mP���k`H|��0�T:�t��!�7����*e��5F*�FZM�=I^ :+����[�0ľ/�'(�'�6ѿM+���1�0�턍��eMH[4V3�B���-��K����3{G�b���~o��&���89#���N+H�g��gL��K�]p��4@|�S_b�m�Nb\���n4&3�(�Ov�b����Za��� �t}i^-�0������/������nF�S��?�,.�v���"E��d#&��]XN����S��b|��G��P,�Q�	���7%�J��'�]3+�p���Q��NjG+���
�lVh���2�XQޭ�V/�
]�~�D��m:�6m�}*]�6c���-p�qs▊oW�Bx]��fr��e�޷���	Е��6�;��%���ȇ��?:��І�'�?���I?!ɂ�1�f�2��^.��s
�[5I�Wʍ΋m�G��L9W���	fx���$O�uU�E���t���E:���n����t��Eˮ�R�5�A_x�l��bs��*^z��F�8�};��[$�5,�4��I�)�y��a@��j�apmP^ ��$�����z ��ar�-Xi�Jh�!`�!���2�,%��ŹU\�N��s�Bj9���f�ԝ�`�q!�k -Rl�k@���n�����8�x��;�z���]��~�Ҍ\����e�fR�V�Y�����>x�+�ކ�ŷ �2P��!��D�c]e�I���ͣq��MWl������g�|���FvI�ő�/��?�ҫL]F�5�`L��ڴ�ڦ�������ˀUѢ��;�^��b���p�����b��:�F�{�
��f~�hO<29n��:��*~���B��f�[�B<���w׵�ƀ_@�{��<Q��:����	�.���7���`͌h`v�G9�����`���ҡ�v#hﭙ�c�$��Z�ųO@t�]=L���zuԩ�֪;���v�{�m��LҦNk�"���l��1�m�h�U��
#���h��ej����ȿ��=K���6��	i�4��6c��6I@�=�s:���*��b�_�ĄE�#���
s+`cez.?,`�V���\����v�gf�XFڳb�+f��ZR>m��-����E�F��z��dBj8h�>��N�^�D^�̍qb���ka,��#��z���K���{�"
��/b	&~�G�W�i���N�}��*I���H|�'!�ݠ�p�!2]�����kj7������I{&`g$��
y�������<;��&6}�+��5f2�}�D"Ə1���$&U���6�hsvjz,^���u
�K�$S���t���B�a��(�qurC�����$� !dzD���Uh~H�2����R���u5���)�*$��@�q�^)����V�X�G�$6�qI[�xR�O^�e�
�JU��¥�m"7<2t8Ƌʺ'�*JS�a��(�C�X��$(W5�����mH	�;I/`k���ņM0����4�^�
�
�:/c�P�,c��k�r��J7([�vG��~f�(�B���ly,�:�E��G�/"��C�,�M,Ğ�/�ck af��t��{����l,n������n	��\����L@��d%}�Kns�>�V���P0�#�5��^����_�
�{���tR�`��Ҋ5nWG���w���]$`����h#J���>�,��o�3c1����� �d�2B�2����m�j����re��B;�����5�j}'��_��_o�pq��ֺ~�n���!���6r���g��7]����<�K�:�	7TJwu���I��W�Ây��pĠ�(���jT�돉 ���b׏�J~.��3f���^ڽ8#��@Y�ԉα|�Z�׿`�Z�T�4@~�A�~3r�|+th�_��C��`���gzx �b^�ژ*��Ζ���ı���j�(��1('g_�W��\kxR�^t���DVu۰�0����|@+�%T�:����k3(k^+�1���;� �����2��J@Ä��Â
�o��"�6E��ߔT'��������X0}��2��"�VF� �'�+X�F�7���p�<�	kh	��gib�;���xZ�ʹ!��5B���T��sz
t
��%�֊���JF h�4A]�cˮ�M|\L�s&0�n��ozqv��v���#�\�y�Q�,]��7�[�M����L�"(��l�+tek&F`y�MA�OH]��.��������b�I� �9|!��e�#6'��]���#f�-D�_H�e7�ch�n�U��`lPQ��x8��7��	C�
s��&V�9�}y��� �xu�-#�_����r�y<_���������4��Il�(�@�^uW0[�|N�|����D�yT��zr5eK�XIx�q��{s*��k�,ҡ_��&�jR�v��B���*���ƥ�����RJ����3|���P�;K �H{�weeR���ݮ���Nʖ� )�	1�戀^&D�m��})�%�\�?n���yX!:<� �)"��w��om�g k�NQc|��ܕ�]M���֠���(|rx�</:�j����_-�&�;����,�o�{�˖�� _����|�S�~q��G�����{9�����lb[�F>R	�<πS��1f����%cG?Bف>U�P1k�/>�r�����=��7+c�
tg��O=	�_��r^��` v�a�{��ʌY��5��>�C":�	rڹ$��t&�ُfuj���Nx�d��R.�<k�3%w)iA�i&�){�����H=4/����ĭs*s�6=�wz�Ϻ? `�U���8\�[��޹x_��B8�h0�JT��Qi�8h݂8����ɺr�+���ѐ�K��]ʗW:$�Dk�Az�Ɨ�
�RS�Ţ�T���m��X��G�Y�J9��̎���	�n�؀�O�<b}��(��	mʭ�K�%�z'phVhm�q
�������wn��g�3/d��Y��Q�j����>�+ �&�wkL�J���8�:��HD�N*�H�r�_�%1��,w�t٠Y�W�}�K#F�Ü���NL7����҉��!s_Aʖ�7v�CeM���R��F�K����d�1���3��w���ك��E/��i���S:Tৈ���L����k�S�^9���qq���`é��|���t�Oȸ�}�G|{���l��U������M �M�Q�E{H�3dT̛^�7�CJ*	�1n�Yic�{A��D����&���4�/h�P���	�cu1�n*[/�'.n��xo,�7< ���i�w�Ƙ�!���1`"}s1�I��f{����S)����Z
T~D��50�_�V���uR��Tf2_��7���5�2.�����!y�Ӭ�)�b+P�656UGc��=d����?S�Օ��ڦ<��;��-�K�)�<�������mNw�@�P��kB�ȝe�C���&/^� �l���G*"5�$8��v��O�t�R͒����ۀ`��~;^�q��ޓ�����ڈ=eV�򌞯/�>�$�'�@f�2���,f�9.)�/jV ����~�pl}�d�5�KWh����Θ�B�}�&N�[<ٻ���I�k۷x�����UI�X�?���b��f$����w޲s��(F8��\	�nv~J�4t�xr�K�6y��ʅ/v2SI�W�n)�k��a>i�_�Ez��<�B?ˇS�{W�W��'t<٘f>a &�aƞ�����:ѮP��-,�h�����5EW����b�l6ta��A�j�� D�P�ڬ���v64���L9KQ��5q�!�x��*Y�7C��iB����x��цMj���^Y�P� ����?y���0ls�Jjj�v۝ǰVA3�g/��O:B��EpK)��������wNA-��A͐g�e����Is}��I��E�co� �S��7���L>DC*ezQ���9T��ֿ�k4sʯ�H�/�X�!��Zԍx�jk|�'5&C�̙��u�e��qb��C2�U��`���xzsn����p��ި����~1$�n
]i܏�w"��o�ö:_Kޝ1K�����iN(kgL �����Z�A1��;#C�W�(�,ҋ��d��8�5
62��2��� ��N~�o-���BΧ�2}@}���CI}�$�[N�mK�ҹ�;�2+C	�������ȭ���>�U50�:v����Fh�T �}� R��18���~���H�p��G�7M�Ov�M�4�H����⊯�yEÏ/cՈ,�œ�͝���/�5���j	�$j�L�8y�A������|�Xi�[��J v��d�h9��޷��Y��^ld;�w�g��嗓;�pmx�[����Դ
rɤ��<0Uj=A�y�,1���g,�.����:�א���b^��p��/HK��b��ŐW��K9���G���Vx���i�3g6�����s�?��mBd�F��}@�r!�3�
 ޔ�&��I�}�<i蜌{�9:���K�CnW��p@��!�����̃�>��2���|�"k
��W��,�9��~	�hT���?����K"J&-�&��Zn$�H�ٰN����~'Eɽ����l���u�;�+un͇�?Nz���F�ʆz/�%Z�E���34�ʎ��W�.$�Z��PI~�����3���%`Wv�$Tq:B��G��X�{
ʩs�"�@#�h������t����_0ڡ`��a�2��h�"y�Dc���J���gf&���h��CV��T���͗�����+ρ3w*XaY�H�C�ԕ5e
�����W
�������?�ҹ�1�Ӿ��`�=�`S-���3["$���B=8��4#g�5"�mvW�?I�EN�gg�n���ϭ��fKL�۴��N��7?�lݽ�9K%`����x�%&\�z�:%����$�X�X/��M����v	��g��8�F���������bY��U� �1��N������&�p�^�G���4AX�Y�}�`|?�O�e�(q��-�Tm�5�O��O$fʁ!�M��FԴ�x4e �q���NBOYe�����x��.�6���:�7!�w��噁8()��;R�=�nt,���G��;���]0���l���� ���~�!f�D�X��Q&��h�vJ��'r����骥u�g`X([ss!�����J�]�y�=���������&J��$�{�̛����:�#�0���CZ
�d�{dֺ�7�>ͧzr���?�E{4��5!!�����{��r\��e�a���T
�^~BC�{�j���H��F��ÝrR���u�����?6�yĊ/찛��C9�ot#<���^91�ȓ�9�q���+�Fn�B�y%�������A���2]-�:�z�`�xn�DX%@�Уv��:T��r۰�Ih��H�Y�{A�J���KS���K��p����sa�G�$��D�+i	�)�w28�%�;��y���*�Jm jZ�TP=E�����`��,Пͼ�}��DZC<�^�^�oO��Z���e��Y��lA`��X<x#��ҥ�b�0�(je`&>���N?���4hT�N�NA�|1��<�/��l��i�Ꚅ䍇���{4V�m����a#5H�R��l�8P�=T>�	�'r�6B�^�)���4~q�!��_r5=��1�r�,�	��7�'�s�&�rݐ�?�O�rꁞ/�'J��q��(���	�0�Le}�.�i�Pm����w��q!-j�����(ےS�M��S�M���*|֫:3��X���c4�JL�:�'��Ϗ�\���/%x x� X�7�b$K��Ð�������q�0�'�u�3h�E:]t˗����y�c�{.��6E�؎�������a<���U�مvK�� YZ|��G~$��i�X^�r�+���0�u�S3��B���T7���A�3E�Q�Ĥ��$�\B��,��_�V�g?:M�g=,(�]���-�ca��,o�A���ST5�� 臸@�qb�B`3���T�w��ݡיA�:�fk��[���D�j&S7�*_��=�8�v-���H :�p$�a	�����b)[���r/���
F�%��А�����lG���x+#��hlY��	�	T/p$�M\-���F �<��
�(�VI�1=SF���i��:����W�U毄�C%M�k7u�HI��l�%�BuO��h��2*
q|�����W��t)���9+�1p�(�J�-�
�;����k��d����aن�>�����[W�2�(�K9�Sa��7X�^�W�E��	| L�N��Π�ȒY�cCtd���G#f�������3D(ҿ&=G��*��p�z�	�ޗ���6�,����:�CW�%D�
ݔ�TB�Y f m���A���z'������d��M	7Q4_��t���:8�vm��Ø.XHlz4/DM�[����}mR噷��}��y��@�{'�U�f/	n��6�N	�y�))�)fR[��U.d~P��X��<*s�F�M�06܈H[� ٣�²9V�U��fa6�����fܜ���&|� �;��Q� ��%�b������E1Yx̣�|�k;p[�]`��T��W�ζB%�(��-C�i�o8�ɚ
t930��
p�v81jU5��LG�VjS��1RF�	�䇤�.�͢�Gg����v%7�`�MJt{�%�"�Q~�5E�Z�|����ʿ4��� �$�)3�&�\���d��s�؞=i�~�Žk��Ò=���꽡��
1i3�tקn�A��A�+C���>hm1���zn=�o�F8lU�����O�Bn���15
�ID[	���ɧO:�=9�
�����ց�U����0딫���q[hڱҩ�:�C�=Ԫ���;���,��T}����1�ua�-��>1X��k%�.�?�8a����.Ƿ)���q���_�:,թg�H=������!��E�,�#ZT�
�+�Â�H=٣�D���󸝔�a>DۓS��RK�+u?v��R���k�[O�F�yx�SN@%%T�0�����Ͳ>,�sDDr�c\}���W���݉7vF�]�����P"��c���e]�.�$�:x��=FBd*��Ci�י�m5#Ƿ�#��i���~���ѥ`�mgl��j-h���Q��:��(O:X�����ȩ�9nJ�"�(-3�:���a�N�Sp��,K���r�[�!>d^������]�������	���.D���i�g�>c�D�ӽ�b�����'�!~��D�Y�7u���](��=̹	�l��)l��Hq�3F�s���$�-a6AJJ��}@�8fW��@�bH����_�_ �0�w�.�l޿���,��븘tғgbt�F6�F�r�K�({C�������
 ��̚�v�
$����dT��c�a���-�։�p��}.B[��^���YQ�/� �q?^e�IR�D������/e��%U7L牢<�&޾���|,/��,1oWa�Bi�u+z��
�G��q�y�T�$�"Y4��i��3	i@)�v:�Vr�����	>OPD���V0v�`319M>��e�M`¹$�(���n�R�i�ӣ��3�gT����9nn�4p�����
z�4B�JR���PG��w��e�}�uWe��pۢU���I|��KP��j�ɏ���䫙��t��W2�ٖ�I��T��\��7�k�?p��?���c�1&�8lG�,�C�<�_F\_n����#�y���]�0�?��u��1;Uc����ImEI1���wI{tu��^l�wS�a�BWv�����g��ʸU7�u�]��l�|r�Ҥ�*qxw�3=��P�Y>�c_���G�N07�K����E��D7~�v�P1*�F����Vi��cԚy,��@�^���y���/]���O����9��y�Uv���ᙄ*�43TP��a��w- ����� e���+�x�F��c"8���Κ�R�d`��a��6�;긱��7��B��|��^��&~K��d�;B[o�l3��!�ʹ����c�H�{���_�7�j�.����k�2���*UQs��^�*�狅2��(�����l)nҳBZ�,���Oһ���	��).;&��j�UAM��YLwJbX��+�b��=FQ�ҙ6�*Pت�T;�FbE)��u8��Ƥ`b�#E$ (�ϵR��0J�2`���(���J��{}�`��Є��p��$t�ܑOw�٤v�~�n���F*����?���@S�z�Ʃ���Q!�`Q-�� "W��r�ea�_hvP���c/� �I�.�jYs"��#ٻ�l��|�y˾V(�5m������Z�.砲a��9V�2OB���Y�����Ðt!k�z�^|,��qdN�W��{����-��uO|~*���[g�2ƒ9򁥶\0gOJT���ۺ�No�P_Q����wb�*�E@p����N�
���R���������>~0�Yכc��
lo\��b��r4 �R9�98���Hʢ�Y����_�����271�M��A.��?q�ѱ�����dv�D��`O�v�L?x�Q\3x�v(:�]V��U�ϖ��5�A�0��Ἠ�`�YH�+&��7:oQa��:0q��][�V�*��arE�J,?r�zkmCYwھbk�t���O�ȵ8�G,�	��_)����_�\�w�E>��E��F�!f\�K�s�n_f�[���O�0Vc[{.I5��\I��İ�����d�۟����;���)%%K�O���q��܉�ܮ]����&?,M=f��28h	������i��Q� �z��t/��-D^+��Ћ��k�ɂ002#3�.b�w�����_�����ՄV�K�#�R���}O���^����YR
a��^�-���|wr_�"��|4-mCk�4���J?����'�#�x�2B,J�NU�9���p��H����;�f��I��7���9^�������Qd������վ_I�=��]y��9����K����6�{E�|�H�9�X���2}W��v�j����i��v�K�&3["�N���ۗWNaǶF@�B=+.��d]��J}ê��t�|e0:,Κ���m�
�Jy�c%�&O�T\M׭A�`MZ龭;��X�WPq4����l�aKM� i�!�8b��` ���g�����ɾ*<�/�'�\�T�p�_4]��Pybw��b�Q��u�y�u&�r��#ǀ�����Bђ�����A�����1ZyC2W��w��H[p�,�njK�L���ꁕ~�y�=[�t��^��3��]+=��E�R��χ~�B~�~�$�6��c���R�o��N�������[q���:�K�T��R�Zj==>�Pٻ����8PiE�w���|��%)8��aX
�ZF�9�V�/7 y��?�Q]�����c1]�Y�@�n
#&��!U� +i��[���b��\5G��$�-Q�熭W�S�,'�y�v����*�s���2���BH���l~����[/[��'W;��� %Y�;QmWR�1¹�����܆L��a�f��D�{�Ёʦd;`٬<<8oH5��S�8ƭIIKp���U���;�ja|/���# �nU��|��a{���.���8:���2E��|�Z���$5�O�,�%5�`�4�Z�������sms_��"���5�њ	p�'���W5Xx��^;0��*�+���6�<8�v��i��vSqZ�lz��|]ǗM�
+�-h9q&�3���T�j)*NoP�3h�D�*h%��{,���G��=�H��1}��+�'��E;�^j����5�E���r���U��էP �`�"���3t����%��՟��!���m�s�Gf�V��6,� O
�d#:��D��.(�B��`
�*����F^#�+Inf�\ݗ͖<�S�aL, 6��0�Ǭcޙ_6�Na�3M�=��St�rM��{(x:@�]��8���S(;�� ���Î�z��N�V�N&�	����؟ҪU�tl��b�Rs^��q�?ؙ�KD�H�K-'	����z�"�~�Lñx�|iB>��l �g��r�|i��C���7��Ä�.���>0�-�N!��HT��N$��_S�������+�$%M���u� W5T&ˮQ-��嘛;��;���r"��C��/m�����xki�ཊ��?4���vyL�[N�ވ����`���/9J0ɇ�U Mi��,3=���!�͍��É?�$&@�m�q�^Z㴓j��^N �Vs�8ړd������C.,�������J8�~���Ù�P !΋+�p�|��oC�sd-�x���{?��,�Y��y��sr�������,F��5W�wd|7�,~-�k)M�x�������GԴ��Lx�C7S���M"���.*��P��$������&u:����O���7��0zM��G�Mg2l�h/��3��.�n�c'�]�"G�B�]�8�X�W>!�09��.�v����.����8]��N����H��5Co۞�W����b��L�ƤT�^é�k�ū���¥fk��&�_���D'�Y�d����P6��Q���F,ǏfU����࿹�L}qNx.��6��rp����`��2���8s9��0���j#�)���9ʆQT�ձ[���������
�}OT-I���2|������m�fߐ������,�n�@�BZ�u�0�����W�<i�I�&�ʇ�;�I���]��+�N�8��'�{��A0���O�"ߞ��X^��F�������tA��e���D�t��!�`<[��{���-�[S���>O�m�I���e�����_M��g�2�yF����4�f�3Z:����
�A^�`h>����P��-�0lI�B.���A�
|�����ܳ`��y����F�]I{0A�+zȶ,�f���F!O�ڑ�X�	�x�p��6\R��������2M�G/�%������1�E=!-�1(?�89`�N٢U�h�Qky���6W�Kێ���0QP6xyT�}y;'_8a�� ����e��.��U8��8����f�Q&/�|���Ƕ�#�d���@A�涩+�9�@v@0~'>n�J)"��9�p$��49��+��߀��FGQ�Ʊ����J���;Ӝk<Y#�h�%3h����,�hl7���k��>��Vi9��)JC�t���M�pѧk#$riO�5Z��g��l]5�RJZ�{̇�:��uh]��]�Z}?��O(%ۼ2\�h�[��A�:X��o
�Ҵ�
�p��ɟ��v<�>�G��>���8G��k ��E5%(m��e&�F������8�ɚe33T,lm� ��ؙ��Mʼ��u�_��7�z�lbwfJ �����7f�[f)�X0�B���N���CK�@�g( �KUn�nL_q�b~J�{MZy�x�������aK�>};[����ՀQ��Yx�"��{�̪��Gצg���먅b��>g��Ug=h��mt��i�ә�ު]�,����L�1<V�Ղ��(]hq�Ը>��A�.�|�:�Fh�T&��/��N/��@�,?6����ki�`�1��vH��FMh-JT1m��`"0�@ct��}���t��2	�@!��m6�=D�6�g�2������2�*�[&�/é�E������z�ȳ�_��&|J�
Lࢂ�K�<�(�'`F:��F)��^�@۵׮p=�S�6� ҳ4�BOcABe�5jpT���0t����S�X��֡�&�k�,�Vd�1r�1�z)Z�Ę�a��
g�����t��J��޶�͡nQ�v��O�vx}����X�O�7����%Z{���ňKW�m��^��Sw���+�k���%�?� ����8�v�5�bN���@4$弰�C�\`2ʶ�����HPa]O�z?.M��V+���.���k�j>#�s�����u�V�<��)
�a�M�\�2+hNgVI��He��wCՌ��|�;%��+mGx|��-2_��k�mI'�uï�>�J�ԅ�ְ$�"�z}�Ȃٖ���'˰ qim��z�Ԯ�ԝ0��i�ל C��s�Xº�:�+� �-C^��t������D0F����H|��qu�.�1�ƛ6��CNHiT�dC���ri7i)�Y�lv@k|Ի�� 5'��Sv��HO���Tؼ�O�6�@�܀ώ���v�U^Ѻ�@x�}l�(Dۡ?�O+���|�r�D�Z�R�D��hK3���|�o��6��
�D��x�<x��`���%;W�K�R�cPCU���B7���)�|{Z��Xv�%��e��帗�<�m��t�c�O|o;���������j[�a�?�Ư��P���[^��h�q�3o�|W����t����(|�#ٷ�cP�����@�n��#�Do��>+	�50x�_F+�C��؄��؁CG�t�)�1ֳ��:��	|�ƄF�\�����լ~���b����܉�lM'gf�0a�,ML	���e�F�;�yw�r>�̞2��
Ѥ���w�G�Ч�M�:ѣ��D�}St ���_���r�ȅ:�5��{�Tר7��aj	��0E��x%˓�_����T�d����P�	ٍ�=��\2Q�J
���]B�;�t��#�92b�ا`��3Ɵ�{�V�H�/9�H��7���aI�qQ���*0#��淸ʜc�F<9^�����&�D��4p�q~���F� �}P۠�ڧ �5e�}%�4��B)2���`�)�]TI��t-��>�bM�ZFpj��u�?|�?���T�6-��	7����u���F��o���9p���%vV6}aL�*�T`��k4�p�b�(9R/�5�i^7� �
��МL�/�B�q;� �q��$�Hp��0���<n�
v��J�i�T#�/΂cs�^YKj���
K��9��v����`�
?v����/54W�e�7T�N�Mh��16�u�f��er I��b�l�+����ڮN��L�q�'���]�#6j?�e�gj�?&x�glCD~����k�akꡀ�^\s�Z�]=�*zw�9LG@#Q�AQ�M�����i�i�fa���ת�#�	i�)�s/�=��{	��I�+y��X��7��C`�����,���^����z�������ۉld��^Yߎ�~��+r'��n�͓�����V�����s��Z�S�E�O��~(�J�츕5�(���>�Ih��ݡ����Z)��lY�e4$�ـ����o�
Y����E�yX��8�Ϝ[@�px|���0�Y�S��h�wB��\�� ���uΡ����瑱������l�����|R�gm��1�<}o���v��lh���%N򦯭I�,�Cz��5���@�#����>4UC%̫���9��Н�t����DmҒ�aŹ�^}�ģ��0�eD�D�[��Lg�Ld��������-׼�CآYy*1��^������� W:�ɩ{}��P�v^L�}�����j�������A�� c4���x_��gԴFO4�k��`�ا�1�M�Ǘ5��@���ڣr���e�䲍i;880��u���tب��qS��;O2C��!��:�Z��1@�M�X���CW��\��S��%u��𕝵�ϑ�|���)z�5Y�;�S~�Z�ES%`��%��~!����&�C�~	�(G���IT�c��{c"l��#sX��(Q;�A��2"��8�}�/M���|5���vi�t>$^J*U�"�}.�\����i5_��,}<V!�q��%!�=C�xK�`R�MY�����+����d���t K�DCh��	L׺�����b�G%�z6��R���v�d�KP�Ut-7�߶�p���z�#2�<8J5-�B�I����\/�`_���f�1C񖶰���w�3?�����R� 4m�x���E?vz�?+��f��ۋ�t5��g���J��1ZN쐹�<l�i4���$(�5�~6�/@i|�~����:U "d���~\dx{|��g$~5!��^!�%�%	M<���t��I�f�P���`L�/W��r7�j���W@!3oIJI�m;�|B��@4v��F�L���见k�`��I�n*/��@6���J�X4NX����{�F��,a�a�<0;d}�������+�f:�^&�C�"��ܻ��i�R y��~ܛ�,�|�jy�[�D�K�gՉ�q;� �{��t^�n�c��?�$敭��a�����I�	�s]L���LKX+!���G��U�=�`��έ�ı�"^�w������r��ԱTD���0{���ڒ�k�S�CĤ�ԽC���66��`��ly�r]t>�Y�H,� ���\����q�C1��Ʒ>@�V�1?&E@;��zt�І�tU�I�G��p�2%�g!�X�@�H�>:g�q�����L��q8v��2q�*��+���������b��	9���f��@�Q��M��X�q�����񂌘���U��=�jnl�������k���u���Z�1,����}���`�I�6O,�%.����#&�ԋ�#�б��P����-��m�4��۸�10���T�{[
������ s:�ã^�3��@8y�H�w�
K����+Nc�DM�k�As5�=}��?܎��5e��'�l�Q�#�e�s]����3�E�'��TL�����B����Ŗ��_��>�{�u9�d�swY����j��?�� ����7�V��D��AE!�@��ģ*>���>����!�� Q�M�v���*������(�z�Vȁ���s�<���z<�+U���,p2���HtT��Ӎ���Œ��Z鋭��[>�v\���z��}���b ���l|Ru��]�!�g��i��L��o,���G�"�)�}�T"h�P��:Fᡖ�{����J~��gO��b��iv��i�t�k�EG:0�8	o����[���&�b$����2qP�p�����a!��
ĀF��*�f)X�q�J�y5)Z��E9���wr�rE:��6����}v�Wѭ�9M�2�zO��d��9�xϳv>�hĺcV�ͤ=���&%j�\4C7���GgVAW�f��؂kN� *zM�v��r*��ڶݐΐ��,��꧁�� �s�¤�-)W�QFm0.Bh'۩y��S'��s�cT2 �ş�J<��)B�W�����bB���9߄��c���S䥰����JRS/d��^�n!Ϯe/6�
����u��b������x��]S��Z��i�+�L^ύ�������і�=nR���o�{����Q�)�h�_l��9)���b��V1��'�p��l$�����Ts�����7捙�̅_�4���&��A���58j�׬3�{POC��[����Hu���X�������JB�h��cJ+��9;�}n3��ա��$s;s���Z��%��$*��x�}̦��E�����j�֫SUDpra�UiA_9dJ��x8�^����g�f��){S^�L1�Y�<�OShŞ�8��E���73��n�z�����ӄ��= }q`����z�cwW����*���y����.t�.�a�������	Ra(ۯH���@�-�_�Ǵ���/ʋh�Ocr�O]�|�߆{�����#~��w&9�B���HC�?I�k��թ��w��璳��LP�ہ˳�,U[�R���Lz����x�FO�Ϳ�e�h��a���M�^�f*gz����؟���
�̊r�Ѹ��`�쮬K�H�u�(]�и��Í�cFqB�D"���e㢡ZL=�J��䗷��C����К�J����}4	����z��SdIQ�}��S�c�x��ܧ+aR�P�\@�W�����Gw�s�Z��,�]����6C�b�E۵6O���w�eW��|��+����`	��'*���4�E-�ב�����HD#�m�zp��-衕�����ۓv�<*Ca�b�kM�L�������]&Ĕ�_��I!�]	��`1iQj�:}���zݲHxYAx���r=�!8�fK׽V��ɑ�hNsI��~�QP��ZC|&�4�D�H����J:ؒ�F�<�[0oUJ�ـ5�U��{$*��3�aғ�u��
��;xկ3Ϗ�I=5�~�����(��I7($��,�cv�K�5�!�oW���[1��%��B�{j��=Z��-D�oJ��~���o;ok#�+5'��=�<��l���ь�����;Ҽ��}i�?U�)T�c�b�J��|��)Ҹ�i�|�����ѯ�W�B�D+��=oPtCʹ�h�ա��*��SAA*Y?���n����^����Y͸�/�2,Y�p���I0F$�����O'Ez��� =f~<����q�'�]��a��y��_U�:K���
v^{���N��m(�mͺU:%_$l�T��a��׵����,<I����ev�޺����a&�]�~ث�Ɣސ�O���� m�r�h���_5��筞������:g���3҉ I��0$ä��"y��G'�Fi����*�Q�=�oe=ok&0K`9����<���r����ɽY�3MeR�%�z��p&M��c����xm7�bL��d�+�(�u�qùLHM)p�qE���_�C�85���~ʓj˵������R�\\��T�Y��7���V8�k)�s��	f&أ]�&��@���B���Dn�7|��/u�t�{�)��=�t3�lՔ�JB����%l��H<�q\O�v
�C������:}���4 %o����2#�^­L����z��`�?�6���S�����|�|R�$J��/�[��H�c�� �gL�)uL%���t70Wk- �SS=P�h1��c����^��:7Ҷ6����s��񎥑���6-��1�K�,?�.�_|
���z]<�eE��-Kõ�ĳb�%lai�-����=]��ֻl�.��&J��cY� ��Y�Lٻ$�?_�M�1MN��IR�J%~�o���C��,G���n���<���?Bٻ<���6���p�,�r�a�z!�;���4�"a+I�/)�r�&a�/s�q����,��Z�l�-c�:�W41��bg�c�1#��n��+�ӝ�#*�o��=��C���h]�����j
����1:ĩn���p�#����$��45�X��k	���bA�5���Ǩ���}ׄ�4_.-(���d;˗!~v*J���-�2��<j��]%{��i�h�u,�6@�a,�E<���M�k&�`�w"�J|ޡC��W�� ��B��9Ƅ_a,�
%Q�D�YFO+t�ꪝA�Hx��-�6���)n!X��h�͏�mXE��%�������ro(9�CE��q�s�m.�D�1����zހ�Z!��ѱu�c��߬�f��M릭�(c�X&�~�j�<r-_Z��*}����AGT=���; ������SOʍi���#
r"ҹ��GQK������6��"�QQ��89�-�3�%�|���X�VLOFE��Q�|��#jZ�ٳ�F�ՙ�F���ź�a<\��Cb�t�D���;T5|�~�L2�Ѳn�����6&�PQ�����'@X'뀻("Bßx~���k �ܯ� p"EEB�A�Uw�u���6wrs��/O�R��G��Ґ�HS����-!�=E3/���J���w��Z9��s������ �m�X#��a�3]A�	}����_2�8(������i.x*�9���;��.��O]��sf����|�|R����. 5����}�!�7�,Z�4��	�$��f&�Ѳ��Ha������:��E��D�;�Ry>�v��ܢ!�0��2FB��crϾ�ҼZ��}���)מ:�� �tטA ��|Bd"W!_�/��~�W��:��_b㑒a�s��`�S�<�� ��X��QU:����(Z�\��^?ىck��DľO�8�JY5�?Q�Av�Y�L����j�"MQQ�I@��Q�Hd��}�5�Ϝ�==��t%� ��I���]��ⶹ��}j�u��%�z]�Ou�v����tr�J�(7�0�
�eI�D�kgBݻ&X�
�5+gz�H��:�/ 8T�y_��iČ9�Ѱ5)��,�R �yQc�+2By�lN@���[N_�U,;*�Ȓ���T�tS�w��|D�t��gX���o/j��3�>φeO���ږNUM�v�&<�`������M�ǐ�5q�� ��L@��w0�]1�`d IN���$���?�_��\-���n��{��a\h?ܞz6*_"F@����sH��ۢ�/��JF��������xCj�8�P�[,����I�8���A
 ���Nä8^�*�5Ow�^��3��L���y/gM.16�!z!����F�_����c�G�n�x�=ZC5�����M�S�h�'�yB�w@A��Ɯ6Qqf)�FTD'��J�0D�\Vf��~,juj�D��t�J�����yR��`'��,�����̏��%ꚲ�V���rk!^�,7[&��<�8\��-u�Y��U��x�~fC!�x?l1B��gB�7�F-S�Q�����w���A7h�ƃ�*3G�zjB��
�?��3֡�a2H��	j��6���r${�h2�Ǎ��M�E$ IO��Y쥳!�h!�V��H��<*��-AzC��|��s�M�����|Wm�R��WL����g�n�)m6�����PDf�,k�\���rnC���*פ(�)u(�遣�Zt��^��f�藩9��j�%4*�p���m���92\�����'�u<F�L.��BL���;�֏�=�V���:R�?$\o�[f,�#�"��l]��D�S�S��BJ���Q��g��N�G!An����>�gr��D��F���?)��W�����v���+�"�6d��~��{�'3d�����e�p��V�W��c<Gp��c�)�B���NߌE��4$ �ϖNQ�W~��t�шO1yX4�0�S��q���V
4���>s�>���c%w0�)>��G㈻�U����s��U�m���>���ZR�W����Bq>��讐��"�%��|�����C����sT�$Ŷi�'+��zO?�&�z)N�5���&*z2`SUuIf����Tj!룥�s���8�M�W���^<hz�l�D{�,m]I�?G�_��aVN�:�~�4�W�p��9��^a�G:#�("�U[���.?�6�l�JX�0���B���μ0�1$t���g��7A=m�ܳd`o��OuvRM���/��ω̋�ʢ�y��Ζ{x�JL;�;�\�pB�jL�����,����.fkJ��C|}(3�N�l椇�	��6��Y��=���$Y�Yd�t?���lD^���iS�p͊�w��52>z�_���8�$.�I�E��J`�.��F�\�w
{Q�5ފ܌��w�֑��wj�2���p�4/�=Z�{���aV�x5`���jY�$��U�S
z/MR����x�x%8&��$mu,#� ���r�6�o[�^����'�~���G�l�h~�œSFv:�7<�A���&��#|�.��G�wg��\��H�S'>��v)G��ҳ�E�K���k��j1����%-��6��xW��~�%�(�h��Ôtg(��D�^:���]�BEb���= ���WJ�� ����>$�^#���=�;�t�
^:�+�y��Ά뷽��*�\��LM��P�������8��^R��<gj;*5 �� �~z�:վė�{��tty_1j��~�� ����3ĭo�֐c��p�(��R��+�<��n�|5*j��0/�/qO$t�rWי���b��ý�v�^��`���o!�瀭;L��N�_}�3�]�L������\v��~�71M�U�+uD��)QҾ�#�c�<�홿�^�q�CI?��s�P������2x���B~���q����]s�1:}:�C��ı�uy<j���@�o��X&tIO�с6����W%�O/�]��F$w������:�Q�s]��bח�0Ke�������7k�7� �1ٳ�!�� �����4���D���MM����ΙC��Լ����cO胔�_r��\��1���T>S�?{S��&��Og	�u�����.�6��kD�y���I'�z�ϛ��D�z�QHG�LV�T���j��|��Μ�@�b#|���K^7e� �0nXi��i�g,����1�\�f���7�i���pΚb��u];��x^8��v����fF_�r 'DpCG��6��h��,r\6ϵҖ �k6&��ʝ: ��Tݎ�6}��gp�P�e��5F���OB���8y#��t� ��ҠV�1$��>�Flh�^p�U8�b=n��<^��Ss3�`�C�T���{nL﬘���i��1
&K��2j#��ĕ�v�]p����L�\��+V�_9��I��#h�5"�K��:��t�6L~��������8 n� �ҾY�c.�h��`��
e�	��G�ӣ�-C����J��rp*ʏգ*�Cb���]Zv}�ζ���ﷂ�����Ps9�	�pf�J�X�i���<N}��RK��g_S�9�	_S�
�"�п���R��ta�}��Jy��;��|�K��Ư��-"�	?ô������>6��p�Y��A����$���v�N�A6�c��[�#W�V� QV�1;q����bp�zG�єU�|��A�!�٩�f)�c*�i�v������ᦦ�'��
l�[�s���ۆ�������B�tkXn��̝.V��x7���U������Y���h6�����H<<�D��h���-�$c��j��{���wm�#A��1�׾qЇ��<�������.ޘl:�p,�Q��P,�T^X�����}�zxS#���jV������Y�*�j���g��8�����g9,�`��(���-t5���[0��*�c{C6!A�쐼K4���>�a��:�)��Iܞ�*Ss*_��ˏb.�S��|y���Q$W!��0耚�[����)�B�zЧ��4&��)�E�������	��Q��8��:��\O�N�_�Ь���� b�E�V2[lYR�?��ϝ���,j�XZ�1o���/j�&�5��v�a�:z���8���k��mv˖���M��{k�DM��bb�z-Tcx��[��['�q!��?���2 X=��	�%��f��1�,�fa	Kd��h_)��g�E��]3�6@s����h�/s�=�E]1ٻ�:�g�v�f�-��8��0��h?Z�D�-���Ϛ71�Jh# ZHU��뒦���`��1>��T��1o*ܜ����FX��gpP�r�v(O*ŕ�O�:4�$���0g�'����U-�&�Cè��xtT(c��uD���[F�ğ���9�k�q+OK��k��
Z4и|��l���^�P�>v��R��*���~���gi�fy:��J)	�z�Ui����Wu{��`^@)���Q�ޞ�>���:��c�ڐ�N�R&���{d�z�p�[��"�C��{j�|��^zS 4��D�1���sP�E\�iF&��:Ow^���ڏ|Gp��2ҿ�yǋꍈ(ÔDj��4YdԡI��]Z�yjۡ���D��5�|K<G��	�8�rjQ+�L����Y��J.}�?-���}�\$�����Q	�YB��l8iH4�(�%~1C��0O/#��cv�$e��|�@'��U��s\�m������K���܂� �����!?���0�Yj�|)}��` ���F-Q1dT7�a��y5�젣'zGx��1ʹ�,s2a�
7�bL������Stnl��Ć�����(�������[5t��b�P���\,���\��2��B�{SM#��SQl�������%nl	�C}�<�^`U�� Aϒ�h�p/���Ծ�=�a�X<�R��&���;Hˑ(��D��A��G����+F�w'�>���|a��n�Jy>��xT�'�s�)
%M��T�0�X�����G�����-�,i�3�:Q�Stk.�_����ھ���Gb�k5pW�8�p���\sg,o�嬋��G�������y���Y</��w�~8����� ���&I*�
4�D ��O�Q��_wl���������68��=���K�I�^��#��U�Һn���twm�Ȑ��GY�E�����;$+����xw���Wb�>3�"R}"�}Cu0�G���^��u9�Vz(P�6�>i��`F�R�+�9��|l�&?|@�X�Ů{v��x"���k.�~	e�g�8\��	:�>��;	X�4[�:0�0�r��>陭g��ԇ��E�ݨc 5�G#��H8�u�];l
�{,`0b���u%��'��yt��̾vHe�/Tӽ�CP��E�BA IK�+{�<����ґ����(�|��w�l��F۰	�uM�����ַK��&�z�uN�Z�(:1��zJ�P��<��[�`��v����c|g��z�(��)r�� Buu���)�B�ȟV��jj�:��o{���{8��;ˊ���a^���M͙�"�1���J#M��w.�{�9��+�Ә�B�]Ƞ:�<�� ��%�M��tQz(oX�����N� �\�ՙ�ɞQ��	�[��B�Y����$���J����cE�3��+��<HԿ��r�]��^��X�{�E}��9���z9��y`��hxx�����u�=��|�����c_���GZ�&�e��kj�m]#�ny<?���fJ<A��mk�,�K7�����=zۻ�������l��p[:: ҹ�!#�c�2���xWFu�k��N���"�AY�Z@KW`���Sº?��g�of�Ēch���X͞���0�f)����[��i�p�<�4��6�9�(�Jh-5�s����>HF�ܜТ�ج�]�Ti�|G��zڅ+�F%Ol^62k��Gj��J�w��o���=a�?���
D��rS��R}T )'A�!3[�M�=�K�����q�]�/ބ ]kQ�O��V�T��,���������8�iƑ��[��^0�>�ZF��ʵ�O�ra�{??���� ql��J���:[��\����U��A��O#(�#�����5��U��m�Qj�Ř�$B�F�V����Es2ya�4p�F����x���Ĩ;9�˽q͇�z�i���H���7��Xi�2f_b���������ĹDf�����>�-''&x?=�)�u�Xzpx�Й|v������Apr�`�\4r�w��1akX���
�%$J�Û���RF��Ȫ0�?0�04���no"'k��Y����N5;M�%u��V����٦��[�U�����v�;�f!���
6"ʔ�O�	��}=O�����ў9?$�x]�ߟgs���B�'G� �bf��q��hj����mg�|��X����墰��y��y𝅉�
Ư�4�e3YB���~�7adH`�⌌h�۝ִ�Y
�2�V�%^��C٬q*�&�V: yf�+�sE�Ƭ��&+��y�J-ft]ԭ����O*�Foi��lŝ�8\������&ha�v�c�)�'�5i�%�l \�{�	4���4�'J�*�%���������Ϟj��ghdȇ���R9^�9�Gٙv֞��Ⱦ1�},�-��Zа���s�#�:����򒹁�p;�Ǐm<�J�^7�u�z�&���:N�\��B��pB��s�OpQ3��3Hͨ�Ў�SǬ=k��_B����p���`���އʋ���o�`�$��K�o�'���އ)�yKG��x�kD�aj"[�V7�L��X�*��e��T��3�"���noH��`,5��C�{���p(�u�:��(�|�7���)����h��I�����Q���_����p�Ր8�wQB��*�|Jڱ����+��k��w�������1RJ��(��>�z�G�	�q��{�c��ڊ�,�"v�0CA#"q��^&1}���T�V���׽�R[�Z$��&�`�Ū�%e�d���i�k��-X��� �(�/��������
���KL�A)K���9,=�}�6RV,D~w�6t�q+�xBQ�~��6>Ӱ��/������e�Ԓ�:<������p����牃�3��)ͱP)��oe��s��qWZ��r��4٘�@�.� -.�E$-K���	�=��J��B����$�
����X����h��� ��`F���q�^�Y�z�m���q����S�-����G\T���	�!�O��V0�`�^�}fXK�蜴uک��0����k;\�r<�ue2���V�4O��&���I4����ޡ4�X�G:>����p���J(P�h_�Ǵ3���r]u$PuR$>�,�Eq_񉸤EH*��|�'��6MYm�Ք���a-G��9�75�y̨+��c�l0��X�n���G�߾�Y��4,�(�oL��n�S(���O���!RQ�[�}��>�vx�ш�7�^�g�.�z��	=yA���S�g�����~9b���@{�+HR/:�ҰQh�����;��#��[�S���Y�؜z��r�ʇ��Q�v;=r���ǆ;�A��7M@�0�.[z��2�l4�s-��Ĭ٤�t��-( \� �d�ͺ�S�򻾈�g��S~�������$3�Qkși[tE�����d�]*�J�&�N>��N�;�4"!4&���N"�} MC1ޘG�Ǿn��V[�vSJ4KwT��e=/����y��W �Y n��ݕ �N��v�'܈`�,��~�XB`X�>b��a�����U�rc�>H"\�!׾�y:������gZk��}�ʀ5;}� tI��%�]uK�賏���4E0vw9ۮ���gW��/@�EN��[��=�aa���w0"�bp���#�7z�"�"�׭s���
�uA��"�Ta���C=���ؗ�^�#����+�'3i�	�<V��$/��K����e��u�'�<!,fGۨ%11&��l���,�o��|n@ޣ�]I+�d�Qs��o�A}S�%$����\���-+��k��߰�(
5�z��u�i�>�@�@�ψ��4Vg�,��s!��jm�n�d++	K�֛5���f�g.v���ڬ-2;�D��@��Y��)/�G�aw���rMpFh��qț�:��ph3"Z������/���1�@9�$)�Vm�E��+9^%ï����G�L��!@!�R"���Ά��t_���z��!�.������� ���_�f��jT�s)wV�R��C��Y����j����ʂ�k;���W��0�e��DKS|3�d���B���l	�Wa��h���l�l���Eo�ָC+�$M��r�nJ��ū?���! ��{�T��Ye���(�-m��3[���J��2�ҩ�㲌��釄U6P@h��1IGS.'�b����]zp�&b��n��ܮ{?Jo��-�T��ta��7|�P���q+���<|V��+r��r��?��Βi/	����J�s���N	ܓ��=c�q�����!���y�i� �$�2qY�����VP�I��=LC|���B�rC3n�EtG�y��rUA����,��_� �n_��5:�M��4��J�-���c�Fe
@Mq������S^Ðqܶ�av<��J�B:�!����;[^B��]|%���>�	��6����K��}D����mg�� 9�HC��0�o�ٖx:�"K9��$�g��s�9J�	$O�G�`�M"�����F��r���?��Rt�O��䭋V��r���Zs1e��cKHf>��ua@i��ܹ1{�!�.0s@��<���K�*R��˝H[=�7��*�����Z�L�;o����&�MM��{�,G}t_�Ǣ�/�zeB�����nf]?�vჃ��e̺�=�W(�Y�0�3ϵrh�r��F?e7^̙k����-�S>�U��C���d��Z����zqY���� Q�UAhNQ���PF����r����.�b�j����@��Tti_�N���`��A)>� s����ܤ}ܧ�A�h�ў��[VA�P��Vu!��.����"�`���k_�\�����b��,��U���dV���7�iwJYH]KG��SZ!���(>a��ҹB������R��m'�n�4b��L�d5�'r��ى�گ��ځ�4�cf�r�%j��jW̒[ގX6#<�=^J��s�{\4�{cA��N�H�����̗����',�
U�M)���˽�N"��#��$D��B	�a �Q�q��xaUȍ\�=�ԡ�0Z;Y� �n�tu�X&����`V����U�{/6�er�ZL��̏�z��1�Sf�5�:Ϡ����0&:C�f�9mVe�Ⱥ�Z������g���uy�s�[)�0QO�h�VnW�rK|�'  xM�s�K�`%��y��ɰ`���Xm�jP�8��tY�߾|̉�#��}:t��q\��@n/pQ�N\��Q��б���d@�QiF���@�n���RF�E4�Ơ"/�8�V�w���Cu�\��<2T�h�v���T�0��C�樾�c41q�S{ ���6�׏LӔ4����aFGP$��|`b0�xY�P{��rbN�s�))�I{�V�i��H� #�Q#�[s�#X�{�f�ρ������L�f�`�垽�最��3�j��V����a3�N��T�[mV��6F��g�,�5He:�ب�G��Sx��'��Uk`��3�,ϕ�:x�i<9��O��1*�Y��bv����w��;
C����a)�/�����_����t�6������RY��#'	�=��T���B��Hs�׽��8R���gYv�]ٯ�
����Gu��P��擃X��W�7���%�z}� ᴵ�fK�,��WK����F�zl.�گpg�%���� ��֡OGu:��q^��N�u�����A�9�|�gx��*:0�R����m�Rt'��j$���Y��_��6}}�ą���Z�n��a�Q�J�*׊3y��4k��a*눣ozL+�0t��(�j�y�J�q��j����#>�H�6= ����R�i^�`�R(kVz�U�Cb�b�[sU�a����ǲ�3��
�X�yBR�EI"H�e�/9�jf!�� TL����B�QG¶�1����W�
"?i��6Ĩ��6d��-��OB�dxB���[�2�O՘��]�z��a�6���X�)���&�����/TV����'{`{Z76ޘ�U�_���C�^�y}=}�^��#UMj*�������*�}̪��jUr�駼�P艶j7�>h�j{��w���㻫߿�N V�H�v\l(Zv.�5���o�����J�,p�0Nx�4ɭ���CƸ��`f*����#�0z���L�������M��/�M8B-�>8aG�z�O��&Z��ݪ�lT����G3>��(o�sJ�^��i��S��
��Y�]J2W���LoP���L�#����m�J��"��k#��k�Za�{0���"��X��p�r�Ĝ�3v�Yx�T������s�B��x���r^,@��s�������I�&��fv�q/>�o��>�蓡�f0�g�u�j�"�P�ҕ��@��ӫ5�5ܾ�G�#����}	y�^r��׭��[7��͜C�-uv/S�^l���B$��t���$��!����93}6�� �E�Գ�a�kv}�Z�L�b���Y��O��/bOG�y���a�����7P+9��Gi6���#N��r1X�߿���	).�#�2�T;/���$ �j;7������t00��]"!�V�����O�~FY3�w�A�� ~��7!���JƩ(���s������Da\x!~e<���+K>uņ�ڳ�:4V%E&�C����^����}/�`���i)�){k��愦o��UC�C5�td7å�a�G����X����g��p!2m����r�+�Ji�{f'\"���T1ퟱ0**���}�A���������Jh�2'�}�J�7#��T�F/۱V��B��8��N4�+s&Zu�� �scO�V�r�qx��5Ř�=�䜁S�|�>�J�X4,�ynM>o��N�p{�~l��b)��'�0�P�O�:�:_�F/�q3_Zd���){���gmr%��C!��ّ����Y�|��MO$���jz��dA�;�i�»���K}mF�2�2��C�8~$=��p�������N�"P��k��(����B�~͒@��+M�P�:�i�D�D��4����_�v�nq�V���_h�f�:r�dK��V>X�+Jii5s3iқ@�V����T�{X��	�U�"Zw����pH������k������N��Kp����0XNKO�X	0h�[EX,N�F:��`�]^��'�S{��F�M|�B�B�4
a�H>�~�g9���|mf�Ҙ���s��_�B4΁��q����8�Fڣ�7���1E����Z#���;�1��a��7�-.`��>ͯ���
��2r
~�c_	��!���sn����$ꇃ�/�K�f��*E^?�+#ƒ����z�\�Jq�[v���콭�\x]��9fJ��8��B܁=/2l��|�F��<������uE��	���@�yy6(��(_����s|��}���Й��rh�<m��W03���)"�(���<��#3�2��)w�NDX�5}a#<��j��d/�A�@1�y�*�[˷ �*�����',>�{]�I��~��W9w>4<WH�>Y���1�!�t\'F�( q�b�"J�&q��(��4�L�ӕ(��7ΐ�����Z��:��򡋱H:�����?7_b3�*Ǭ;>B�Z����1A��9ߖ��\Z�5��ϻ����N�n#&�5�i�0Bǅ��$���K�[T�Q.�b�z�b����a)�a���i���xݕ���Mܯ*���Q2\Rh
 �ɕ0�S�"d���ETW�)��c0s�3��}���ي
!j�&j�䱴�������.��lQ��v2��i8�)��	�)��b�.'���Ѻs�F����`ph�
Y2s����3ȆhK�y�w�#�OW^��_j�􋿏��F(�-�����E��Ρ&9��I!��pmS�*�͉{����I'p��~�A0�wb>X|i��#�յ�x�����si� ˡk@BB���ۺ"m!D�@�1�"Tt��#�IGL��|
PVI_`Й��f"�d �A�$�#�~5bJ�85τ��U��\ၔ�(L�x�������u/�/ F�a���h�5 <��𼖱�,���{c�9�,W�� ���\l��JER-�����۸��[�ݗ�g�]�)����* �]L�Zw����I�DhLjp��2|,��y�9P���Ҩ\!���l�!V�Ot�;NORԳ�Zy<?6X�?	[̺�������&�����4��&��'}��?��yT^�;�H|�!E^o�����LU�k�h_�n��5��[���0�C���7~��d5�\tx�[�*��IϠԵju��H�x�n����.rš<_��;�-�J�] �c����\����^�$B�)����G��f6?��b,�5I�앷����M�T��瞩�;���� �nX���T$�g������asƏ�|�	�:L��R���8�;6N^ؓp`]�AM��A�7i�>"V��TJn��+�Z�*�z���Q�,d8&�4�L\gt�x8��E�|��j�M�G�n��B1-Q��R.���l���8�k�t8�6_m��Q[�#��#p?z��^M�[2Z띐�E����.��
��/�(WkOn;�,'t��U"�gg`�q�-���>I7�<_B��Q⨚i���1VUs
۱|���U7��Ӷkh��ֻ�)�ƶ"�L����p͌VZZ-=bk&�Fr$I�CpÄ�{g
�7�&	$��'f[p��Z�4�?�W$3���5Iΐ����-pw�],�	c�K��p�Rs�S}J.��+5��4���![�Is`O���\�I�jV�5�M�*+��0����%|]N��*�`虡"��zV�~���wD�wH�������\��9>3)I������+#�=f�Bh��H��ASf��ny��pq���j�@paa�Kt!6V�/\f�н�8o.��x�P�2y���xȆ���A����W��\���]5 ��%���!=ޕ��ї�e�N s'�SC�K��|;�{pxHRXx�l�n[Pݵn�*vP�_�T6\&��L&�3���F��JvF��X��`P�Z$�~XHk���qI�W����C�7�tir���7�8Z���a&Ϗ@഻�@���ď�pc^@�I��M��T6�ܬ�y�<d��*��� �%_Jdj���f�G�-M�uS�V�~����]���Bd�ퟖ"|n��:� �'��)�Q:3Ll����je�	O��&Uh���eZ)W9^\�k�~Ԟqp�V��o<��$>���^�Z�+����8���2��k�[����F=�B�<oNn�$)�?�=H�Ot�	�2-���oTF%�d����D&���S�~8c!���k�4����4_����Xp���>���@��3��5=ȉHn�j�/	�#��Y�x_=jq�a�h��pwx�9;�됰������!H4
���E+%"�>����Ml�j����~���^�����⻟͝#��9n��#l�_*�;���1�����:L�ǸT�X��Cr���&�`cĩڷ,�;��!�?�8��Q��ּD�~�Ɗ�#�N�n(8x��w+��Hs\����\
���v��v�.�}�,=�6!<D�5��z{5�V�VY��ۂ`�@xc`�Q	����x�x�[�X<-���K��@���uK���:�W�?c�b�\�7/�����~��>�����hW`�!�s/����?�51�iO�h���m�OAK�j����5(���/l©�H���~��j*\ ]S��CY���f�Ps+�l��}�dx��x�+�\f��'L�`��p��C܀�G��^�T9u���}N�NZ���O����v�5*�d\	�I}�
Dʡ��Ѫ�.��r�r_�|�wкW�A�l&�?1��5���
�������-g(�GI^\,�7�0� K7)�8��VGf�O�c�j;�[���ϗ�~Xl p�\���7_���3�\?ls�=��4�|I����߂B҉츎H�T@�"��B\��xc���g�K� �t6�6��e�!�bz�榳�u�|�"T}��C(��aδ��Ӵ����-����T����Ζ�8
����	��.��;J���~Z��O?�[��6�zAegs�y����4����� y�
�V(qn�z�"�y�_�	��4�
��8�=hH�?5ٽ"�f��Lx�7T��b^�,>�<{&�&�a)+���#����cVW(1����y5���T@�;�:��=��o���.}VS�1t���@�jOv���@�t�W2���[4��(@t����%2��ʒ�>�eQ\S2!ք��c9XQDgs�pK��)����=�4e
�~8�0�s;*T��/�Wp��E�D��w�>�`^=/	�;�w�����>{����=�f�R�Zf���a#�T��~I�D���}�~���6I�C�׉�#�����x�xʲ,�*���?�Ϯ�1��L�m��\���I����d|���&�*��Y�r�(����+�����E���� ��iF�;@C���F=���C��͔W����A��zV���_��~���!Ο�օ�khb��͓H��	�)��m��w�M�e�B�BY�"��ͼC-�6�'���´��eɥW�w��;����tc�Ĵ6�B�Ů�� rE�O��E��ю����d|C0^c�֪Cic��&�����M��ăw,w"��/Q`D�	��Ҟ���v���&�F��dF�n���7�� 
=���vŮ$���{�!�9 �7�Ǻ�%)�3��X/��5�Ml0�+�LQe�C�dh�L�ܠ���:��.M]O�C쨺�L	�5���.?3��)��^%�YKD��_w�Bo_���^�\}yk�VdCV�l�����P�1@nǯ\`H�L[�-j*	ٔZ��2j����^���ᅺsWS�ɹ��R��a�9ArF��ذ�X�,��J;���=��8��ځ��V"��������s��$��/M���F�	�n���:j~�=\��?�`�k;���P�0#��)CRЉ��W�l*Ʋ� �!��.:ꃶ��m6��K��g�N4ׂ���Q-�Q|U�,������H�*9����fj�u� <չӄ������h�7j���.Yѷ��-��9/��Y�­g��L%ѥI��t���N<Ǿ5��Q��ɍ����|�˚RXawDDy���Y��FR�����j�{+�m�r4C��(l��
��U���<Lp��r+ۼ�b�QaʼrBF��Xa0Y�x�)�*]���H����-��'؂Z���ҩ�UHA~��"�����h��`�R]ˌ�O7�Of,CO�=�酊D�m������1�7fk8/��g,@���&|��d6_�s,H����t�D�D�f�o%�ݾ9��>�m�{!q�y%L��@���]�>�B�z^�HB�w�7B�c�\�ǝ���M�6��O�{��'7@��+�0[�ի��t���G8C�ԁL:yɆM<�@m����t�'���d)Ӌ^gp�r���c���U>��9�����T��%4W������R��}-���j��X�1�F{DԖ���/�T�	��
�F�:i��Lf[��(�[��t�U�:-�S$�d+/N0)�d����h|����
� �?^��/��E���d�,�D&�S��i�y�LW�{g22�3!��ў��z<�61����"��A'O;S�lWϟH�%0�������9���7e�n,��-ަ�÷���Ä!���LrXJG���2�(�N�%���v�����n�{1��.�_	غ��AP*��.o�Q�r�G��� ���#�1�;6n�p���{�/;��t��<r��S��O.�Nja��]{Q���r,��GS:57O:�&���*���A4/s�Y?�W���íHR[�׷<�_1xC��k��ܵl<ů����`��A�O7tzfA(����"�m��^~	�9Њ���Pk�pͮ>�2��Ĵ`/��﯅�j`�jU��8�ҾBK�ҹmx��3JWyT���������?6�����LC��(�]okA��x#��Ҭᦶ��cr�i���G�Ee&�6��K���6W�`���rQ)o���}��J1��<��/���R|(��P��*���7��s��c��X���|�뾊���.�����N�
9FrЈ��8���_s=X}{�/���&�{k�ڡ|�!�i3�$�#L,%��,�FAy.�P#��!������}J�Ht� \���L(dç�\1�0��� R�Z�tk���t�َ��S�PO�M�$�*�8_"������m5>i�����5����?�M����1<||#]f����7��׋�����5wN�l1����+�4���ePͥU��Ө
�iU�ʌH�q�uM࿍F�`���@t����F�J< w�I�r�z�^$��aK<�*M/�B�\�ם���=�T����[�ѢE<�k� �ns���qާ���U;U��u�J��ze��	������-c�鏕��-5���G. y�����A�ߐ��n�A�X��
�擞X�w�e�� [�
t�ƭ)�ё1Ƥ�p��<r��u�BIaA���=�����\�.�pQ(b2����Cg.�6*�6�B*ϗJ���2�q�@�>��&�"�򵌍x�~pe��g����1���0��>�0R��P��:��+��H�������ͻ�� � ��=S�$9I�?W���h�{��C����z�7,�}�x�)JG��
�j�u�����n&�wx6T�*
�G�xݙb+�������]<�֢�u�� �S�mfM�f��/eo�yb*ۚ
��WM��d�?��s�s�ˠ�+mna�֘�!21��EIbE�~����{�/j�h|�^��H���$�"�.�sDE��*8�j�w7�j�j��P�ܩt61ۗ�&o?�*p)�2(����c
�f���ђ4�OBv?���9��Xjn�WCe�E|�t?S L���VTrw�_��������e�\@'X�sͪܘn�����ȉ9�/�v����U�Z�ǠD���KU��w@���K0���?��`zJ�+��n�� Q97�*�~�qo�D�\�l�rAg��W	�^���9
*�0ߛ����n$�-��`
����lSD0ùR�ec���+_��	ƈ�3����񘊹nދX?��k�m��.T�R�2�<�6�j�{��p6��Q�dE�3絶�DU�MU*���{����6�!Gm�Pͯ_Z~U��pʷ�H-:4H���m�ǻ�ֵ�jn���i�9;J�@::{�3X���2��fC�v.�a?y�`:p��x��#���1$1I��w�,��P�N`t0�`���d����{���B���S�>����P�p|O����O���F�0P{c^�<;=ʐm��$�ۘ��ˊ�
�"o7c������X���d�4n�WA��9������S8�{����s�;@�T=8��M
�+�T뻎�,�f�,j�t�eF�����J���S@I�U��jkh7FN�A֏r��}k3N�)�)^�	E�ὀ���W� u�����v�==x��H���f\��i������u?��d>�l�I"x ��VjY���)Dp"�D��%��-�RFOIz�8;�Y���Y���x�J��;E�z�3?�ah,&pzՑ�0>�!�����8�x�o|Є߿afa�Y�~�����IH�+4�B�1}�Zi����_��aØR����-���az���'2/����b�H�@�1�o���%����X�i%�{5R�
�^5 ���������d�.8l
����'�CӚ����G����e�-�W~�u�L���t"�gⲫ�X���>w�ɨ�In&�SL��E/��n�+e�֨�x��}��F�#r�ƮD:ʤ�`�����\t�SIa�$!I�KS�B�o�sg�� �9�r�ǒ�����T^�~RcA�p���{�]<Ը���&z��S�k�����S�݊-'R��'NU��/�}���g]p�_*4��n���i��7����W�-뛯
;��;��bM�(L��񎎚H>��o!��3��M��K\��b��:�ۊkqi|�|�Y���= Ȕ����x���U����%ڮ�%��m�.��;�Qr���~�@F����(��������dy�&ҫ.�����(����ge^�(b��-� ���
�ģZ$P���B0��*�J4{--�_{yH|$D8Bg�F`�ap/Ф�u��>�I�� �@q/�b��^f��P�(�ﱥ��+~j��>�w.�`C����M�(8��F��2�="$p0��Q�n8�Έ���K[��{b�E.̩�ן^��[�֫��C9�?>q�&%�G������t�g*x�q��"2�P�`�N�=�7ʉ�:5;�x�ZCH�>�(�w��R	��]�(���z,�^�=��
 �vw�7��R㷑�gԙ��;���dj%�D�X39u�������
�����!��vs�*���y@t!Kb���/�^�ͤ��9�����Q��`tU|�d_/��D�'����Y��7'U²	���������_hOv�T��q���c����
��ΊX���?��±����L�z��
��y<��G(���I<5�G��;�١�l�����vv�jF�S~m�S`����W��K������{�����a�b���3{��4|�HcF-�ſ��pbڼP=�B��I"��󉻷,a0Ӿ��#�3��q|HSB�q�fhL��_!k��J.��`+*�]ީ�J���� ��������$��i#��Ks�� �)<�X���9��O��6F��uE��Z�2�����!;�M:���;��Oc����L�}aax�5���)N#�9�VK�6�$	"�nA&"3J���L0�cY���A��'�FuK57p铐ٕ�F��X��)`k�-I�X�~I�^NZE`�>��VNK�����mU!�ay��=���d�]�>O\���*��a��ȍ	t����m��̜hƱ�]�]�Y���q�&<���'��Z�%��!�/�������e Z�V_�~M���e�@��b�C�P[��9=��:W�5ƈ��Vt�C��O�Y(������2u����k�����i����;2�G����������!�Y�c� v]T�X��F�>��oO[/�%ר��ar7��M�gaxٰSIC5Ր ��^�4�Zq������(W{�-�'%�غ,�L� �=]���:���x#���@OZ¿P���S��������ׇ���]�����fwS��i����ۂ��!��:�`�yޅ��(�C��/��`>s�i�7US$y��-���E�Ar����y�\��9���zW�!��q�б�N���*�m�_\�8+y�\�:U�jQ�w��1r���mY�r��������m�e��_�H�jm�^��D����g�����[)&�2�fH��	�SЃ)V ��޲�A�-��ѽ/F���dF�D����a(!�ؖl�)��x �d��Zo8���zV2���ͳG��JW�1*�,Β����^n%�iQ2��8��x1R;T������ƚ�	[�hM�"R�'�s�[��dK@��ɗ�!}sh/I��\'t�A��@���-��M�Fw+������-�/%��Fe�.��5is�4z����3�f"��@E;7vN�����@7��$�ގ;�%cU���<E�NȔ�#�L�xl#��%N��Qj�q��j����N*�7�y	��&�ҵx���T��g.W�gIb���e����LY2�ŀ�7�Y� Q��=ш��65c���(P���&�& �oc09�j,S�`���v�DK-�gT����ڮۓ�Cr�@$�&�Mপ(VrG�X�+ؐD��3�(�fy>7��ߏJ52Fܢ:��J��xY����3D�y�)=������K���0�4�e�(P��n]�P��1��=��Ec��G�\@�hǟ$AD`����A�����R0�|���`����F�w�y%�㰨��{���v����n�����p��@���q9�{�]���|(S�s�NH�4׾v���y;���.{�Y�]�FYU���x!_�w)j��+B�;S�f+}�~�oY$b�6���{R;�$î0,����,�T(�^���Y/,����=�b���n��Wr,̏@���������O@���XP���O{�2,�3Q;Ѿv�9�~݊�J(�x@�oޞK�	���+��[y�
YN���x�<I|�;/ߔ��n1��A��d���^9�p�~]H��l7jェNF�"�W�l�.n{��D��j�W�l�aEbr7�Z���$%Em+^!������=��$ o��\�-Q:fZ�sB%,���¬;G�P��=l�k)Ծ��Sk��d���V��sū���\d����u4��p�jp�C䟟���ml
�Q�&k�@bu����'8��Y˽�K��{v�ڟ_�
\�++��;�J&m7E����o>�Y���6e��O�P&.��=]9��Cd0l��s��#�l�9�8z��{v�ؓ�����W���W�=��#H�<g�W8�2�f���˝�j��j?�\��{2��g��Ԗ��?_������Џ�ئRՁ�'��k�:F��T�I?���7�;协�ȍ�� q���x��R'�~���ɮ5-vͼ4�k��vOˋS����v'��\��ӗMo%�|`�n]{v���}�NR=�ac�������q��È'����p?���?ӺS	�������n���CM����G�J܏�з�����oPb�	��]�D|�~%�J�ȗ��8(4H �����������I&5]wȆ�.>�w�����A¶˒
�f�Ki���$r/�c�&-C<�<�����r �p��x�3/]��D��vMS�y��֠��:��qS��|B����ΔV2�jG2z꩐ig�n�$�	�s�R���Iei+��y%�	Hl�)�{�tɍ>޳er�bA}ZI
�,	S�=���Z��P闯�FY��md�A��^1	;��Ҵ%QS+�rX�&��I�݊�!C�)���Y��|ט+���XO�=̩}pA��=S�6�;�cQ7���b�k9�9g�わ2L���5g�)P=�ϣ��ٖwC������!eة�����a��ł��i��?�l�	^,�������?{#�FW�`$A����-�J��Jj��K�6G�z<���*^���w[�XݚI��QT�����a}�5��t�6�#��ʵ�50 ��i�P����	+{�d��S���U�gޔԹ
�o����<\PeI���5������´�f�2̺��-��9S|jP�>�M��w��̓U;��Ef_���]~|ulR�1�f?���^�
�[Q-�ȅ�%��o�Ӏ�c�����y����{��]P�S�����Dl:�D޳�8�4u��m�Ub�1�J?�D̄�W܆���a�g���\��\S�g�E�ْ�Pi�To�ޛ��7�d���^����Q$���D���/O��Xȿo��f��� GUڲ��%�h������\#�%u�3�YP|�W������DA
���3�yQx��Lj�#v7�um{J�OD�:z������jQ�w#=b��ʖ��ԑv��S�����MN�F�t� j��$hAxw\.3p�rq�%����Ve��33�TF��R���R'���#�\V*�8�j��ir���;}��$R[=|>ţ�7" �N�� �%�>S�����E��yU�Hς�f68�6���|�7�~�G��*�,�$����p�Z�����y[�B�~$K�bA)��O���i�#t�t�ȼ2@�gv�~A'F�3�h�tj��y�X��Ϟ��H��F�S]��[�H�K��3��ըq����c,�|-ʮ,O�,��$f�L���?"��<q��󝸋cV*����oU���ɲ�=����Z���V�hf+�Z�A�Vo��Y�\�KY����"����T7��9=v�e~>w�󢼱��A~�;�32��58��e�#r,��?52 =�p��y���'��F�������6	��L�`Y�@�wG�x�ǈy#�Z{Jy>�b�B��S��:u?�������V�)d���_ʈ7�{�����#�\�P�,��&Ɉ�B��)�58�Cu,�rH�����bj������F����k*r�.�F��M�Q�߷��v�D�7�[��n���S�G/9رꪏU^3l��Nt�S�,�jg�ѫ�˖u��W��W�&�8��+�l ��Co�n��7��v���2�a��M9�-���Q��C�����d�|1�p⩣O��ﷅ#��Y\p]��9���To�<�m��q#��gPl�E[��ް�z��d�E���(T��|<J����Ol���=�
"�U}}qs��X�GX�g�օ��H��.l�? ��7�i7��S�#2ҩA�Ԁ��샭��(��3�c�Şy�Ic���V��"��'.,j*շ1�F����!<+�❽_�	 _�dם8����<���l��k-�	�s郕`L��b����m��j$h����Y�f!?��X*����8M�л���9���ٟ�ꫜz�7�}�H�-$M�1�ξKi��|N���o?�~<[�l����TF�<My�h
��:�o��|hzD
�hr�j�_�k��j�Tkđ�|ח9J�)s@��B�9��$�������7g�f�3LC�S�H�c�_��<�w��Z+Y��}���  ���'1H�Y�MH���ɤ�}����,��~@���������Z|��E��D>*��c�sь�!�������D�2
��!����3�g�s%����?@��g��S�!<�܈�-Gm�u:��.燊!K�z�+�m� T�qM�_�uE��)���L/�/R �8���~:�RQ1��d� t�������NREm<8�4��Zɕ3h�%��G2u�/G�d8�������H�Ԕ,D�����a�w,�Ǆ4U_v Z�Z�΂z��|&���ke�q�vY���+>���ojE鑆���g��-�`��i19#mO-�����}]��бy��\v��%���}޹�M��˷���[s^m�GTGh�a��`]�?�Xo��Nq������*�a��9�1K�Ğ�[(f8\���݇�%�V��I��Rm�4P"���kH웚3W�c�kC8v@�!G>�ݕy�}��u�Rȃ����y��=w��1�~:�W��W�4��� �8Nh�����Q)X�_Ģ�0�K���	���Ađ�����|~=¿\��>4���=��{��A��&���%�A���N\�`�V2�yU+?p�"�
e�G�:`o�3�������/�R��Ⱥ/�p�,���Y_�Ds9֗�@d��V�X#������|�֢�#�qa`q�#���D?r�C�z`�Ef�ܡ�2Uuo�1&�!���2��0M3���Z9/�F]I�/'ﻷ�|� �P�V}A�}��Re�v��p��A����~����5f�>{I<�
-����M%�+����7�)�w����4�)�@Q����06Տ���k�wH��ޥ{���Y-Hm��e	
��]%�;PuwX�$��HM��Du��-#􉫶_Zf<h�.�W�������
�!y�����&lcm� Ӷ�+�3�B��J���'+$$fr��_NFf�K}gT[Bu,v8ױ�%�_ONyI$4l��|Y����`�'aSʥ���I�H.�s��E��ʟ�wA����Q3`	�X?�m�@����q���dMs7TC�lCT����:
��RA\#>�g}���s�Ma�mN$NCՉ5I�����F�e�(��=g�Q<1sH=�%�����l0M�=�P��	5Y�G!��&��Hj��[t�a���X��"�Q\���W���5���+Y[��h/-<c�����9�#�~U�agm�d(��ܦ�oE�H��;@]����E'�J����m��Oz�
tJr�Jx"�=�Y�G&��r��5�FN"�mF׫w��Å�*b�E�o��&RA�F����Usv�/��6�m�@���z*2?�F 6s����L��?��G�7vWO4;<��bn�/����� �Z����h"W�fu
Qރ��Hz��k�`��6y��U_��(uE��+b�E�nd���Vbc!r�.�[�K�T�Q���..����@Ru�N�+7,�A�CI�Q>,Y���yɾKS~�Y`
��rx��I/�o!t���<�:`�&����ȥ��n��>.��)ya�=PLԳ~�sU���C���Jݤ���k���Z�,ˎ�!���(��zx�W��	|��k��R�>r&���twp��q����D�L��B�a��������-�ƈ0��]}��#���U��v�<~NK��w����'f�n*�/Sh�!���2�J�H[[����[��8��T�?0���SyP0�!�5�x�2�6v��l�z�q|Vb���hJ�A�Uf��q������ x�*���n�OҊ[e�����TacL�h�:W?�E��՘:�|�WS[�c"���)ū�k��dE�MJ�1����vr�\�Y�Q{�\�x��0]�j8Xp=���cz����-�(;0g�=^�䳉t|PZ��m���ֳt2�� &��T~���-<����+-i���7���b�U�ٷ���s�>͞�?'e�L���Y�\rg׻M��|
Y�t�@����!���Yߺ�)d�upxT�ˉ��+(�d�>R���`����6-�L�S~b*z`˖R�es�N׈4pw�P�Tq�FEe���\�z~�����3��!K�u�@ �e]yG��?���䱊q���¶�X��:[8�Z��D�{�b�-Z,�Hij4F~R)�����ɞfY��:>Q��y'@�:�4�>P�>I:���uI.���~�6������]L�ԶN����U@��\�)rj���v��u`��%ϜD�&5�Sry����g�֤�W6��Q�!�6B��P�?����OD���}��tj_TQ�cXŠ�HƧ%����rA��Wu\pJ��d~D���F��Ő���5�E��n�)�AȞA't��j{���G'�R��v�Ճ�^���t��6�w�/d(n�
���]|�z4V���IMWN1��cL��^I�f�] �Ճd�1|�]�	��e��!��� �u�H�e�}����ez�6n�j�>.|�e[�U��N87�b�͛pV���0���K�"���m���̈�U�Z��F���5��t�3�^(�C%H8��E� ҕ�ꠌ�]��R?��[q��o6��]�e��'s�v*���{0�HR���T �+CU0���@Gt=p9�ҫ{�'� �u��-�*��Ec��	/P �L��<U�ɊB�����4�Ձ�ؖ�>��F\EsE��,�!4�Gn,����ӧӰ=T�_*����/9/5Vy�g��M�O���1�RH`�#�?�ٽ�wD��6���������.PvV�@�{AF��	ӥdڙqf��f[��1�Q.qУ�t�_]S��7T#MT�� ԉ3��I
�k�Ӯ#�^U=��~zu �=���Pzg��x8��ɗ�KG�=�A�ȡ��/|ʆ�3�t�Ȣw�����M2���v�{
=�`�4dD�~pIh��Ahz�os�}\��T�j�-��7�4(8�D��Q+k�2�끐WJU�O��rzԏG��\V8�$�bg� ��jh�ܓ����C:��>'�.��V��&���LG���XcL�\�������w��D�C<(����#���a�u�D��HEy��p�X�e�*�]h����3w��7�r���4��R�C�����]��x4��P��m����w\�Z�~��﵂�Ә-�93f.�:�]����6���ƹ]t/$��p�V�	9��Ƨ&t@��=���نf=�b�l8"�Жx��'!�9��j�_3��>��2Rz��ި2�*�5+�}��'"�x��P��L#b����o����LJȾI'!r�:���;o��T�h��I@�=�dP"���'���.��Q9�l�����������T�,��&��Dc��/��Ϸl�kb��1��:��GP�?l3�Xj��D�kH��'��C Z\<~'%��-e~�+��m�vߝ�c� �w��������Rk���
��B#��-��%�P���C�q��*��2�œ�:RQ��38��R��~��9�K^���5?������Ꮣ����z(���&i�X�	f�7��Qg�"���#�����'!��k�M�Ϟ�[]��B�]h?3��Rb��k�%��ss֧W=�]���em�EB��j>�C
}E�Nh\$&p�1M�Lq�q&nO��^�O��k͍[�͚�E�>L+	��mӭ���R�۴8�N�������'�ml�X�dïVtn6�QJ*yI��:�T\	Rq}��������9'���/�޴�ȷ� ��[��;6�:!�6���昮;:l:��M�M읖6���Cx̼ÒL�<��ӑ�Z#&�C��Ց��)������X�;�l��D+q�S��ӧh 
�J�L�%K���D/�k���W�
ބ�q�Sc�AM�lo�(�o���������"bz��}�	�d?�9��_F����Ko�=|�3� �-��w��`��]���K�<���'#���Od�E�Y��48�"x���2�9����N��H�/o.)�C�[ �(�*_J7?E~��Lx��:5��/��M�Ɉ��M��{�+i��C����j�G�����kW�W2!�Z��WS@d6A���5�6��^{������o��d&TSߩ�w*��1檉���H�5{��-��(�kP��4Ǘ�4��V��^��vp�kJ��P�(ݔc��1|J�/M���k
��\����ֱ�����m�ֵ�B�c3J,�*=�W�� nxf*�����e�J��ض�D�uge+C^����� �mp���]�^c���t��[z۷�Ay��>>�K�Sbxȅ��NwQ|��ku5�>"��>���L�
oVv�Ƨ��|�}��V柺���wz�b�7*��z١��OZ���F�7�ӫ9�6"đA{AI�h�t[k�_/l�d9�^�X8R)�4,Y?5p���?Ⱦ�#n6����3u+@8l�2�!N�R��L*j128ӿ�̴�Y_Ezd�4���:�읡�\
6�(��'�%��"����+z�Nk��!�g+-KE7ɀ��k.��h``]+VTG����4'��ѢlЈ��K�j$����Z� �<S�ՍZ�V��,y����a'��?������<~Ǡ<8���W�#h�Q�.����'y��vTI%�h�Y�s`	���Xt+�k��l@C�������,�,�Wz�L��?^�V�lS���g8�mU	9�h8e��(�X��	B~,F�&��˺��"��hχ���o��+��c)R*��ޱO��G�J�����+4�v�s����Gpb���\���4a5�������M�q)*1�}�&�-�w7�l�A0[i����]�EζM�Ff��k$z7"��L~��h�a􇢧�{��Qq���	�>�BF�"���� ����փE C�_!4C�� �_�X#[��S�N;w4	��v|Lw)���rMq����Y������p]w���݃��wt$�u~����p��L�_g�FTR�_z�\��BsT�mD#���w������(y�/i��M�B���1�;`��F'ﴟ�����J��pt�{�.O�d �"�p$V�猀a)��Z�PsR���&�WA���Ù'�-��AdNX�.A��ÙZ�6���^(�dH^��iEK7��}��*�Uj�b��=&�F�i�Ihb2ז$a�PJ�M�tIw�w�-�s�48�?�7�|�� ��!՗����!6j�@��x�~��#(���32|E�S3�_�.v�x�þ$9`，��@�X�t`�a�s�8"/W�Y'����%ED
���Yf*s	3��I:�:t��c���R�*��eM��{oK/u�W`�<�lc��/��@
G�.�1�I'�%�ݒ^$$�F��D</��i���D�֋�.�a�E"�g��dԦ��+�������"��kC�ji�$���#�jw����Yp��ƛ�7!
!�F�>����6���ugtx���,��w�>;]�� �kӶV�$,�m=1�x!l��1^�'��7�i�Ýs�e���1����򚫒6��O�1M�x �b*�o��]�	�����9�{�*�ׂob�=@sԯ��]9��"+����J^�kp9���mYq�&�IɁ��̋�@�*`�y�J��,�3#��*����L����9�nn�=5xY�\`�g����u� ��eu�E�<ޙ���_SPu��֓`��;h[%�d� ��[,��A�_N��;t`�i���$K��y�}�s/_-s��f�f�*�+��C)>R����&�Y9����^���?Ѽ��^H�_6#n�>u��6M��_]�Z�+/XĞ�稼�\�&�-�,,��mE:R���jF�B�s�*��\Cr��*쏨�gYE�aE����Z?�\ Q�3pbF�RxsF��!� �'�*���;I�����v��M���t�3�*�f�wd��W�\{���%0D��� q�(.h�!㹬�S1��;�kY�̢F�ZC��:>���^�^N1��6��0fj=��V�*��<�)�!�-���Т�� ��خ�r��� �k̜8Q�Q�x� ���.���슃x3�Z��q춤�P2(#�$O�J��a�R</�D���y_j�גbz'AP�!��pZ,z�wQi���p�-�K-˰�E&jn"=W� %@o���&R�a7ki�^���Mf?Ք��h�����zZ��e-\����N9]�z�*ew�yFhX�����?Ig�f���V��W�NGE��-{f���Z�._u�2��UԴݾ���m<gg^��l����"��W�3J��E�-�$
iFئ�j��۠�>W'b��A�Ɠ�;ڍ��;FVh�XO�\��@PMS�b�_�9�>x�{VH*� ����>�^FB�(��Q�0�{�m6�D��$$ݦ,3s��2҈�"����U�F�M6m��:�/�8�H����׼G�È�L���0���ſ�S�k�[H=���*ȝG��Ù�|uȆ�u�t�Y++�?s*T>ϯ�v��-	b�]�JFf����+˄k n��=�/�Q$V��ne&��{����Gv��'z�]�͉�Fh`�V��Pcr�N�|�<Vd�>��^�✫��o�Q�Z/��7�ʓcV�i��g�hM5oǲ8I?�e��Dm`*AQ4���mA�×��*�F���N��5�\೪F?�\�p�?t��Hb	���7m��u�v6_�d�91�*�jkY�}�IZ�Z����ՓĈ�Y$-�a1ڠRz��n���=ʹ<|)�*�32�FJ�_�H����L�(��2H���
��g���N�*5���t�P��pU+xڻ��R�I����|�(�D����>����>Dkn����ҫ=��+G+��������8'�jRtpR���*��j�}Q��i��mt�:&f���d�9��M�y#D��J~��`�;��s'3CR��P3�s&ԇ�m�fle�#Kƺ��x1�p;s��e�� ���e��J?��m�m@�e��o��m�4�u���!e����$�\��s����� 4��:�ۻ�o|P��d62;=mr�}`CԦ����<DH"۽��!j=r��&9��f���(
'6���=���#�����0"���o����M��)|��M���L�ر�J�6������Ԭ�\�	��`ڦ��ny���]�������S�I!O����H��� Gl5�����?5�ٔ�'�� {y����Fk��}�K.�~��*%���\\��tנs��Sk��4SFo�ۂ�q����V��v]�`X�f L5P�#��Dx�!�s���p#�td1�h?�7���*G�}�~q�!�W֕�Y;QY� �G�N���+��]�Ke)��0�s}��u^@��+i����V���>Y�jJ��ǈ]jRt��s�
�/��H���׿���ћ8n]X���KîsIɽ}B��}�U*��:�6.D�Z�Q|eab3���ӏ:��D}�߱�H�W�)�eO&�:	����D�U�4];�Qv�ګ���.ir��اʞ����o�SE}z>�|�X�8}���S��X`���z�u�oWㅓⓉ0p�	Y�����:��
K\�l4���w�|V<4�۠)�s�
:qQ�&Ysjc�du�i����.��k��c�]qAa�<�ΩUGȁ��π%�]}i�%�d0pO7��n䤘��F�<�DF��f���a�_�u�,m�P�w�����y�=��oW�l$��W,�v��=����j:�V�K�:���o����S1�f{���{Y��pj����e`,u��qj�`�G�깛.���͉��RSk��S�O2������&��ǃ�f�-G��$dF���y6)���U0���s	�lM{?P�ZpƟK�1�c��*\`��� W��Y�j�����p���~k�l�Ud��<O~]���%Z"����F|g5�g\�s����*����Y!����:�D.^�@XAKXe��Ԁ6\��-���l�[���4.� Q��qɻ��΍�p�9�r�9���:���#0�����܃�'^��H���lJۤ���A�c��ﳸ����74ԣ=9f$�tօ���2*I�y��lj�2W��W�	���OB_-j�Y����e@I���✸���0�[�I@��A��F�Gud�)��ks#&Y����逪�M���� �Pm�d�ࠗSCI���鰙�`5b�_�m|]66�&l���|�z��(�)gv�.�A�x[��1��5�_ �I�*K�|���%�g��6wc7
��"�w��9X�|SC���y��?4p%��uq}������2����]�Q�d�"}CF JXM����k2���Uj�wjí��:oW.Is
2x�{�H�S�raY瑡�_�7̆�(�#�'�H6�_˘&A�ǣ
�*�.��nIK�P&�)X�\�\ v�����w���H5P�~���&��+s&�</����'��EjT���%����w�*>����y4�Ԛa
@�A2J��P~�O���zg�y�]si��� �jӋ���� ]�îd�"Y�#�j1(��-�3ų�Q�[§�ξ�,��VB�3���[P>��ȫv�I�eT Q�l�M�{s��ҦRK��omЗ�tN��w�ÿ���૿�������mz1O=��[.u�X�2V�W��S*��}�N�����O�݊~ym�K��D'�c�3b���r���R5��[pW���3�i�I_��X/
��0%��ec�6���b�������1���rc�Twڟ6O�T	����Z*gZ}ʩ��?�;�ơ�ƣ��jk��I�����\����E�S�F��HŚj�ro
�g��Q�ժg�����F�������y"-�LeB���&K��J�Y� ��85+ډ�
u{x-Y7SBڏ��t���:u '�Bȅn&xIT1��q=�ܿȪ9]�Л���P�$g�L������\f��f���	`��3��E�@eT ���㒛�[����ӹF���إrݑ>���O����2�(��v�3|l��N9�|h�������e�,rYuO}�֏��%k]r� ��9A�U�a!�c�`˿���K,|�2���T�*��
�KI��źu#�D�`UiYf��N���T�f�wDb���S�����u�s��qbb�6-��ނK*���Q�D�[`��`��"��^���n;�kh@Za�Uxu^�⺣�����<��6����\�V.��b�a�Xdq!m���%Bi����n��|��8ӑ��yo�
�����`0��+)�O�_�
ߓ�=d�`܍'!㼸¬1݃��$u���N��Ϥ|D�4�'!o޸����+V�R��im��;t���z��qK�Ժ]�i��D��UlI���h�Tp��u,\�dPі�5IU�#>�9f�i�4W�c�ѻ�MO�y�{]�b<�4�,�}ʺ�)�d'��BTg���c��{H��xho�I/�o� �!	�n����DOx'� ^�0�<���"��2���?���h�t>�����j7N O��y�-�'����##�Nv�� �eD��uZ���~�5'8W���
��fϰDe,]�����^�B�x��Z!������t-Qː�]Hڸ�	��� �Ao�k(�9��,��j�Fj��q��s��� G�&W�]�N-'�4\VL�'dnͣ	����N������׈�̾���D���БhZ����V����
�]�:-���n���&���uTq0���c�#U9�{Pc��͘��x�VK�#z:lw�'�$��k���(܅g�<��ב�x(��6V"�3�U� P�(�ñ��,��RՍ���H5�)М��5Ia�
�mX�����, ��s܋}�װJ�0r@���ƛ��&�77��7����ٹ�5�5�~�w���%����=[k�(�)�3��#:��:�f�F�y�0{����E�ꍣe}=�7Kټ9�&���'f;�.6;��uZ�Ѩ�1���[�{�m����Z��
7U-ٱ�Z������p`+a��&��.ȭ�ei��9e:���ײ���r�L��8�ϔ���H��.���8�³���f,qy)�	_�`Y�2 �3�?���k��׆C�L�i��)��cUB_p� QG����Hx@H;�*.@]�$�����àż`�0��Μ�&�
<&}�H���F�L��p|��Ӣ�)�J�c�g�kJ+R�:�bO�.�P�푙�:��g���X���l3=�Ge�`RR  h�6[���e�8�A�8�ޱ�VcxZC�"=i:�d���-G�[u,��uvGvI�"-Ԗu%8:�������۠�A�k�yK}+<�,�=d�$D{LW(*Һ� ,;���+��$1�(����?��e&���� ������OjJ7�D��db��V��Gc_�*��A�3 ׸|SWE21�}�IѾ����ќ�Y��ū�Ϸ�uU�<���9+�*n���������Yϓ\w6��	���mxA=���C������\�yu9��F��r,У���� ��Kww�[��]�?��r�_M��u/�䗒�RET�9�BƭDC�ҥ��ץ6�YE`� Y�HAS���w�_ZU>��͐����z�����g�>���� �qM������Uq��Ο��C�Qz��H���R�
����A Zwr����J߃�$�̦�f�M�Մ���sD�\�4��� _mxTkw*zˌ_�`/
���ͳ�Ŏ䚽�L���J��(�₌���������2��󘵹H�&	R��;�c*�5��q�8ץ�\t��V�0M�E�1lV���L?�8�!�81%I�5�,"����h�q������i|Q���0���3O���H\��`�G˲���dZ:�.b��Z����w���ݴh�l��޶�:0�Q��$���8 �X���{?F)��
4#��"�RU΂e��X7	J�1]�@l�ǭ{֫<L���$l�� ����_�@�8Hw�o Sb�������Ŭ�Ck�i�#���ʬ%�iZ�} K�3��Q�&�����k�&�2���j�#5�uw�W�.��ɿ�b�y+w#�l���.�;��Ә�4Im�B'
�媳@_�T�)�`��B�*��s��҄��Ղ�
�R&I�52�©����Q���E���������|,�-�,����[dZ����g����ꊶ="�������z�<{_�=�@[]ArF.��s��4NS2�M>BB�O����~`�l}M5�#z�؊R=�_y�FHҲ&�-�:aރ�l�#B�4-Zߠ����c>R֡=g��ɉx=��F�|
�Pl�N�
���˧�G45�^�z�nZ���i�q~E����q�a�U��{��t^ �HMh��j�3��+|��)f�06+�]
�����I�=*AJ���lЕ�E�NA�".������j����g�xj�i\}J�������P_�$� �QF�Ac���d��9�C���N��6ͳ?�����������LWDh.$z���fRv�4?�CMk�ʛw6g!C<�0�{�,�s�u�E��&-w�h8d ��3�J�9�����Ф�l4{5/�,vۆ���	�Ts1]`��U��N\gw'���`�q{�h��ǭ����T�ȯ�P��pM���2�m�]������[v���n;��νWsa�޻�&���Q��)�ܷ��r��ג�惿�b�ʼ20������D��W�NW<�9�2��AK~��]vH�
�urh�YUÍkz����1F�MD�С(��ׅ�M���E�Ͼ�fo'�3e���<��(�WJݺ�f	q��P	��	M5�f��`T� ���5����y_C��.^GW&itD-�3�Z�:�[�,1xrp�6-A�s�jP�l�H�]��LK�i��G+��e�x@��W�n)��h]��~�f۩С9��zYij��!A��,�0�+�����ݦ�Pz��gߴ�h}^�;rn�ڪA�1�t}���F�0��&a�s3���û�[b1K����lЦ1A��7lL�6e��<8����5�1C���|��(ܙ4��Q�$؊��^q%���(I-����bR�q�2v[��M 0|Ox�j܇����O͟��ă��_ƶ&_��d�=v���ӱB��=�i,M��1ӠDW��Z�Ъ�u3�^���#��#��
�U|�g����;��ca"G��Iid:�)���H^����Ha�!�"����u����8bQ`l���/=,�K;:�
·bc�*�ہoŔ#���b�f�2�W�Q�W0��:��ޝ��2Y<zy�u�����6�����-;֗\
Z�藟Q��E ء8�)b����׺��¨�J�!�Fc��N�e�Ň��^�e�^��&�Fs4��Yҝ���TiZ�(��Y%2:g�pBO��6(v�Re����`g�H�;�;<=�T�_���y��#܁�vf�*�����@���}�c��l���#懵����Qv�"I�"D��h�v�)�B�'�g�*����
l,D��P,�{�H�f�o�8�8�T˾��B��(^�V�H�y���K[�J,N���- ���� �
��x��Ys�6��K7S2���&ƚ�ݕ-����T]�`����S�άeK��o&��O@�1����'Q����`��109r���X"1�!�L��,rx�V����φ���޵����5�<�(-�IBO��݅�D����6ͥt��aa췑Y���!���[W9Ʃ3X���D�֐Ҳz��i�����g4�(�]Τth=k��r3�d�ʰ�6�&c��� y�t�7�dz^ʎ^9=�,<�y��wrhvXhun�o���NcEL�ڲ.<����Ĝ���_� �I�F6-��*e�E�f��a�y>�bV<y�AZH]�4���@�����p�i�f��l��U���R�!�be9�>�ޤj�.X8s���nR�,56I���\ͨ?�ys8���٨~w!�7��Yx��o3:'h�'���փ㜤ؑ��/�0�12�4�,�p��J	����V�9�F�[���D���&`���6>:-�kq��$7���-����\�:S���5�.	�n�w�=ޤ�q�J�t�p�/l�<�Ӯ�:Q�c�����Ô�*����> �..N��Yt�`�䏘���G]��R����k�{��������?΄�hN�+���M4$�O�'�CTD��$z���Ǻja
Z�oy��_(C�\��z������Jm�&�l��d���i�$,Ë�SpG~+g�`ԓ���I8�0��g�~�MVT}�#j��':���:�|)Vv��R����]5��~ij��г��{d�i�<�R_�[C_և& �Ρ���������79� ���T���c���ȱ:���9.��$�(�]�qd��E=/�������|�!�Dz��q��1k�3� sTIO�u�H�^<o����{8�l�Y�ϐfs�g��V�n��ޏ]i@�D�Z9�KI;4�,�*�^��>T��'Kj;�l� ����M����v�Ԫ���^���r���Y�|yo*soYߨ�O���4��{��-i�c�.T�=�f촢�u� ��N1����M �Nqi�M>�s�Ͷ8P��%�鳯OTm�О�Ts���0T�9�j�տ��z�8�)�����r�0�@�~��tka�
��f���Q�N��=�e�\���F\�����.#or�z��Jz�sS��6w�,�-r�" ��Jϥ�a<
*M$T�����85��5ൟ�}�z��#��*z���5q��6�B�c�U_UH�|Bٹ�jY6�f�NIJ�.���{��[�"C��0��kNS�l���b���E��Q���L!�3t4�!��r��_��2ܢe�x��A ��yQ��c��R*�ƨ��ĭJ�ǋ?ɧ|��Gq'/t��&	��,�_.F��\
���\M��ɭY��t�������1wш�uI���W��mS�eVۑ�G��f������`m�e�
cD4���&'�-=|�ZH�L������-�t�;��O�UdlYUd*�M̏}�/h�ʈ����:���5��i;���#��#PPGN-D�K�u���Q��ɭ���Ffʠ�����nl�.�X�\���>�iw�욈��Ϩ�V�t�p=��ْW(e-?ݟ��Qu�_�e���9�+����9���R�͎7$�.?�9��������1�@��C�"^�SW�� =�Ye��e6�sg������2w��qM�m�Uݜ�$z�L��l?�+��n�6A|�����������J���$c�,� ��a����4;���A�^����`z��DlM5��3l��g_�|�.����f�(�/���e1�ax��{�V�T�'ߜ|�S�>H����'�oDa����bA�۽7�Q�KiG(BAv�#llM��e��d�0-�OgĐ ,r�a2E����h�T%$�gBO� ���;0O�7��Ss=P%�h�jb3�/��?�+qckN]�tBF`/&��R��C��� Y�#ͅV��	���+���p��v\?V�J���䗻˅�L�Ŭ���,OB?�~��[�7z����5q�0wv�{�.n�>jT�.�����N���\��q���rq����w�p�)d?�y�֗��8���%0ҤV���x����E��*��ܑK���а�x!rF9�3���n� ��PUB	�r+IX��[���6��K�-�������K�����R�r�E�f�I��|��?�'b���*vj J�{>�b�(`bgb�;�SW��l�ѱ���J��?���O��]Z��8"��N�)�o(;� `���nxU!>�MY�d�1:8��{��+���)�k�s��UۜԥI��V}�=ш\%"Xx3i5�߰�g�g������<��� dA�J/���׈�=���~�Hh1�$'xMH��?c��v7�$��dXH�)\���� �I4F����D�G��܌>
w�V����	=�:K����K����n����O�}��e��Y��.�-��Or�+��-����+���ort#T��bRКB56���D�L�SU�H�Y?檚�a��C����X�Z 1���Jx6�Bɱ;4eH� �o6����Oސ�d|���@����J@�n�<o�!�:�ˁF��<>#-��8T���"o%�G@{I�^�D�^5�#Fl��m�G�:O��i�T!R���%"k�h{޸A��6�(+�jDo��ZmM�t�S~'�O8�AI4���b;%W�[���-�z���4�g�?�����㙑�%D��R��C�I:�d����J���~�ܵ#�Z������f������6/�X��kkK�:�����<����a9W���[��:��
����BNņ�R�K]U̻=�-�
t�8bk�e��5��B�Q?y�zOw�l7�a,7i+8��t����|���� �s��CA%.Py�v`��<�`U�X�m���(��Zw�&"D���%�uI1�+��h�n����C���$���#�X2	
?��C�@��jZ��Թ��k���l�d)���
rl��$�Ӟ�ǡ�@�����t	w��$�)o$�Ԡ:E�W�R��c"u�k�����~�����`]^:IY������c�����/�K�NA�~7���e ����)v� CN����Պ�h-2�QW���6Q�>�9���;�r�C�X`���6\i� ?������GΛ��i=6�P�u�%�	=L���l�l#���N�	׍VH�ۗ>
G}�*�D*7v�9�ʍ���2�;5� ��Ky��S+�zm�l/X1B���R쥗afG�`� �-`D� ��~=�z�wp研O�6o~�����`QO��^�!�X���,i���s*-v�{���S�O��-���"Q�V�-�� &�م�4&N���ԩ����T:�a�qz�wr���u=�I붲���E�.!�������#��z仛�xd{=�J0��#<nG+�#�}�u9� ���#�J�V=�֞K݈��k�A9P���h!ml��ɫZ*�Px�����+�c�C}�:E��hFM���J�+��Bd�WN��)�{4Q�"޷Í)�J��{DC��Ͳ+��P�$5�}n[ؘ�#ir���1�)�=q��Q���S�	�}�Ip��G˂�Y1��FoI���ɋ"c�hy/�����nSp�C�up�D�c�4Գ�j�ZݑBh:u{�^Y�v���r7���K	 pU��ʕ���s����q�M?P�O�eƃ6Dه ����2���;�g)��k個p�WN����+�wI���|5���z�@�G�`�2:������ŧ+֞fn�".%��A��:{M2��'�|�u����:N�=��}$���E��T�1N<"g�
�B��������f鮴n��''���C�'�BV\g8��Q��� }A�����paY���t<�&R��_�Nu��Ñ�W��xq$F:�f������H�}�KE�u]�ݺř�gf�����/�.)gkDG[3���ϰ���>4 �j�L�cZ!ĩp�+00� �}�;5t� �t+1`�c���Y	q��8�l��:�>���'g�h��}l���Z,7d�ȟ�עy����!��h&������+��Th����rZ:�1�87���H
Dy��&�R���tJ1^l�������A!n�!�,��p$8���`���m�٨& �x��h�8�:{;f�a�d����-�&!�+��'�O��nO����S&�֏�w��?����tBˀӥ>N\��|;�SS-�Ǎc��$���~sA��G��^���R*�-z@e��s_�{-����x΀���QU�)�PD-nfv�W0�S,�q(�$pjB,��+LN�"�@w���N|�:W�4!��:�4I�ak����s�k�'�w��[��&��}���u�4z��^�HQl��hn*�-������v�AY *&��C>R{��P���'j���>@SCC�f��.��!�D]Ūf�f�4-0�d잶#�d�|���� ���@�|��o���,�:u1��BA�WJ�_�Ǟlv�����/��TgC׫wY9�����Oͥ�xے�f&[<�2]�������4O�:�H���{���2��,&|7�#��P Z}���D��^�-<ӑ�@y�%���+N��4z�{�o�}*��Y��":e
uc�9x����`
�O��M������u-��Ͻ�U�o�%~-+&;8?ψrJo~u�w<T3���P���K����mqg8��6�*�x�m�GXjF]\-�"�� 1�E�@.�[K�����%�����rh�����]���a�cU�8j��e���8�{���uU�X5��KP9��VRU*U����j����M��G����:�Ŧ}z3�[0��H����qd@�\*�/�M���ݑ��(��Qe.�#ؼO�aԟ��dag-N��?��xkR5���n̤y�\\�}3��������5��|�&D�u�P���B��	@�X���N��S�O�!�8�Sk�Y�O�{�}ښ�K5��A�Tb؞�<��a6uXvt�j!�
��"�xP�V���B`pǩη������T�YZ�F�t�U�󩘛ξ���`v�sӗr+
��/�Ὄ� �}N�y͇�]�ro���Q�S�7��>@0Pq�_t@�C�v��h�[�v�,��W@F�pԢ�e^��O�wz��5F1�����g�k�%JkZ����e�\�����A��e+}憧a|�[ס�X8�ql�گ��f�,��7m#�ef`�8�Ɂ����4�YD	]�]��GeȾ�'��=����A���cҺ5�IC�ym=j����%�)|��	��6ƣ�C�C�����);STuY�7�W88D�����l%:;��X�� V/*k��C�{uC�������X/�&3Q�o����]4�I�͊۰�6.���9U�K�?���Z&����t.�WKw>�p��(9�LScb�����S7l�IWz�%9@���
b�� �/�ٟ�M7����0:�4�i;Z��-�8�A�a��lp{ȆGsx��-.:@̆�w�*� ?7i����œ�{�N�-vMD��@��,�W� $�����X;nDxJK���6+ͱ����H������M�KXP����}�;�T��	��Њ+�W�6��l���S=X��S�+�Jqa��CB9�Z8moC���d���K�Ijd�X6�����s,M�!P\�,�"����BQ�M��0=EǞT���	$��-�+F��t����1�+<�]�@���j��YjP��qZ��2�j��t�����	Yd6�D,}� !�7q[���z&�6j� #1f�vx��#SO;oZ��dY���M�Z[4n��EO &!�fn��e��!��1z�U��׻�S�D������C/ϩg����('D��G�?Z�f�6��)��U{���j�Kb��ɶG��6,���{>�HAk�N9�:��8�W#^����1�F&����R\n/�.G�R�Z�>�F�;���M3��R[{i�wY���2"���+�U���dSǛ1������3���#�4�C�./��#�U����\��F1Wl6��|";K�\`���ٍLVeݱ����,g�	z��M���Tk�-����T���u��uZ���jk�
�R�̑tqUM���5.�Ц�m��c;E-�N�[�����^�a��+� ����@q>?	B�
=+�@:��5I󂏳`}�
X���c�lT��/��t���J�����YҜ�C{���;B!k�xX�zүr���/��z�����d�r���!2A��6�L��`�
e����ypY�m4K��ޞ�2����R��;̎�'t��X`6N�m*o2��eSsM苂A��h,x���uv��߅��|�8�X/�#�����х�Fn�Q��$�3<��� еΏ��hn����fÏ��Y��C$-���,�\�[�
��^���R6Hi�6mV�Bn�U�#l��=)�tB��t����ӭ(B��'��=k6�������Jlb-�� ��KJN��1/�
�+�)|�j��A�j�����ñ�v�Z"���U���G��!�/J���h�]I�$l�d������� � ��K�Š�/T9���Z�����6vp!��3�↡��Sd*O�.���Q���K_r��m\��K�^PI2I����f�;��Jkɺ��q���o�uH�s�V�Kg�F/�ÁJouG�Ƃ��"Jx)6F�����A��R��9�ŭ��;�$Si���C<՛���m�2���%����E�	�����"�o�#�������2@%�x��Gf2z�1ϔ�b�a��q�݅η�Ĵl-ƨ��fc�"��/	$貥�y��W�Ri�ԟ2v��NM��b]Vb3&,��ﷱ���xV�Q2�j�!�H��}�J!?��v����b3����vb�'�'a}6
�!J1���6��٠@���^�K�B��
�܅D����c@̸ci�(	d|�m]ț�ʜe�3 �+���h��`��ltIH��G;�b�s"���	���R5B�,��M�"7�]��V�͒4f��(��c/׮e�-Z��������(O�"K|� $r0Ɠ��NM�馉W��m1_�.���ԇ4[�\����I�kb�w{N3#/�yv�9�ԅ��� &U�Ҷ�Vvn<�7�8/� �h>���M&����
�yhbl~�x#�-�I!�����L���|ZDf�ń�'R�ֳ��\�6c��:gH9F}&x�ȁRd[sg|o�����m@�E�r��՜��)����R�˃Y��-�MY9;�f��IݎE�F]��N� r�!r�Qh�tK���vM�!��*��[x�c�IL���+���v��s`HL߱-t�o@>PY_k.����w�d-��J1��gG�����ǞV�E�:2�\%<`.��[�~`>����__�xI���ֻ�3wء�|c,t�穧G�؃�y�LX����ˏ}�}��%�9�͌��^�U�B���#�4G@�`��]�� B=T$.�<=��d���R�WI���c����\���Us:
_68Q�kW��V"���A�V��BJ�~�Y�B�������T��)��~�q���ҙ,�Ut���hFG:A�;>�F��O*#��N�"�i�\C@�"��
y7T�,�o�զN���0,Q���q��>�s 
���K���!?#0�H;�$��Ns���n�||�'"��;�<�*qZӼ����?L�����ֿ���4�=>��b�{�_˙f�G-��|���x��RɤE�7�~_|��w������a�R:4���V�^�x�XT����mz��$t�+B��L�R��qa]N�������p�U���J��!��H��e9��+I-�NDh.JNZ�~�-����ñgݰ��f��F���-=��G5�Jc�|������nת�y��G���������J���@�|Q2���ql �L!b�}�:5IƊw0L�)z(@C1�������e'���4WngFm��C	���b|�P&���[!�Ak���ٯ�U{U��i��j��Y�/��i&�j�C�"a��)\N��%�v0;�\�G��� 
� �SZrg힪&q� J���'�e��(c���/�P_��C��R��Q7��p�HS��G��/���W��zr��sڄ��]�U�:+�6��T7���F��GT/��6�ƴP���\�ʽҟ���V�����kJ$JN�̡�=�|��h�>��0z����;� �!�1���*�D�L(�����o��o�z�**Ȏ���s	�47�̑5-X9�Ne�����r�_�55kͥ?��;��0����Y��'m� �����p���s�����A-��~w�� �VHȓ�>6r�5igFgl��~aiNZD�6�b}�������,��~�\Ǒ��e�cG9>��#�]ܓ�FM�;�H G�VA/�v5�I�<ŵ)_4����:e5 �c+��s���nc��>�3��kt؏�:� ��
�<*Ɣ���-݌O9	���z�Q�1`�~�d1�ЋQ���\�~R(��t�L��y��EtM�<m��Η �.�W����J��h���2s�:�Uv#���NUD�@��[~�OF_��x�,9M��'G���2��5{��ϊ-8&���5�#C��{7��RIQ`k�qŋ�7����$W�@˷���i ��f��ʌ,��,�xrS$̼@;�C3y����a��I�o��l������tRFԗ��/f�{�[d�K�<$x�V���!!�����%���x�=mrTК�r����<v��e��؊8���P���u�]��xX3�����ygt�S�] H�<�M$����d���@)�s��e�E@�t�(���fb��<,\�czd����H����8A����b3������!������yu0_�'I33���AP�Iw.��x����1�C�!�vz�3�9+��=����
b`�
�zu�ټ\��mǙ�� ���!��'�L�t7]�m����fY�����I��y?y�~'��J�E����!��hX�g��ao�� 
��%T�7MzH=_��nu7宊�E���T'���;���Xy���·[�)�]����D0�Ӊ��E���ݪdښ
Ζ�v����E.:�s�b0���Jf�~oJ��ë�E�y!0��m��*Bx̄�3t�D,7ի�&�I�l ���_<K_<��'���������M�Q���k2x�U�.��9�9�Y���Z���u��EO"��5�/�3���J�sb�{�k�]H��&��q<��lm1F|(�6�
���D�e�K�&EA�&P��ƏGe JD|�+��t���^u>�+K|8P� �R9������R[��ѭ�z#%��0�v�ݙ�5d<�s�6""�'��Wu&���4g9V~�EәE8ΟW��T�b��cS,*�?�PTFaD��FY�?t+q���$��_��wY�H"�Exѕ�7���N�]��b~B�a���ê����7^�+-E��jSq���*��9s�mJ��ӫ�,�n2�Q{@� ���s"y@vN��4C&�QK��O���xgP+�a�yo�356�rf�p��:��V�h��I��wT�DW��Yl���
�W9�RC��p1~�~:��D����GX���|j��ϫ�Z��Pv�]�=�?;���� #��O3Z��bL��(JgՓ�G�
X�s	�H
5����u���$��㖝���U@�R*y�_���N���_�}O��/�ʨ��H_�R��<1U*G�����Cy�H�?��ɏD�99!��
��bZW׋�Om�!��FHg�KҪu�>H�剚�\u��w�fˏ]��^��c�S��}��'Zj�O�.<{H���d{[��9xN����������iS�{91�k�+H�kJF�s	�ka:"A��!Q�5g"{м���'
N�8�&�g��uJi2/��.4>��@�G�����آ��/�ݥ�����(U�}C|����'�R�W��B��(N:�IX'��~5$z몴k���!�I�r$�Oy^h��(w��[�k9+���Vn�����U��}d�������%����@���ψg�q��F��zi*1�n�Yڦ � ���H/�Ǣ|y��K��E��/JG�$M�����;Iɻ��	R�3@�?�.�{��`��5U�+���r�����Q�QcMZ]H,�J(������m!W�;+��`s'��n�ƨ�k�,C;�+��J�O� CM�s�9��Ϋ-�OQL˼y��~��fM0�(���u
��!!hqn��O��#���k�$g4�/C{�I���zg�q�.����(Ұ%1@@��O�.�Y��z�oʐB�@c�e� �5djPtg�D����������=B�,(��G��2�>�u&܀��!P ��-�Z�����7;�(�ǜ�3��T�à5h�7��~�j��E�f�/�������V�ä�i%R���2�SC�n���i�̌��im�"kX�q��ʜ�C	A���>I_��Gz�_�oH|�MD7�~��I&F��;�OHr��"�r����,dh;|��Y5}��A��O��&�!HS��w�)��ȧP����n� �.&e����Y��K�sʽ*����2��Mc���Z 98i��=���Msk]Z��}�Y2.�GL�`9+~�HE�,�q9�z.��m�$�ƐN���>sg)t0��a���ݺ�J6�I�vte��E���lȳ­Ն��G�mP��Y}�N9�;�)��#c�Yz�,�Y�Ӥ��5��L����JS�����'s���BaC�ݸh���ɾf�h�>����.0�.���{�*�m�����p����F��P��q�� ����AC?zGW�Ӳ��m\%�fޮ)�N3k��W�Bd��e���X��@���{r���x�Z����v�1�~�^z�L��L��ku!��PxN�9~h��խ9������M�)}�Ց!l�
�����jy��l�R��bQ��T�az?9��^���^L�&�O�xj��@XQ؄y�#W75W��GMtg$��:�^ɪ�kn���nw�17�K~�tY��_���[S�4Uu	4y܃l���&�ץTW|ɘ��+�Et��=��a|�ɖ����n��F�B����������z*gH+��҉�TW�i)>=v�O����C�s������_�=I'3�F�e:��������uw�"}��p�Шza�k�R�$�6�t��39eĎ��(�d��AX~_j���ݙ�]o��ԏ��=��Đ���\~^W���>�ʷG���HЩ��d(���ΈO�2K���	���F��(-%���@���-��11��ܨ���ܱ�v����{���WWi�w�^D�@�Lt�����K��Sr�f��hM�f��:�+�����|v�B��a\$a�<o����Ÿ�ǋ[�+��'�]�t�e;����ޢ���cߙ�<���q2�I.]��AH���j���Mн��� QcY�%:��aH�/I�	iCj�x�l��e�,����Ia���$�`]��n�LaL?ֻ�:[�2Ƴ��o��ԉA/­B��tp���Hb%����"��!l?|�NR�m��DA�K��JqǤvO���R9�d�R��T��H�C�s�=!�5D�d�3C?b޵�ahh�!Zj81[�!ąu����I
��O
���a�H�X����BU��c�2Uf�_Żkjj:�T�O5���1A���^�2��S��sM��M�ŜgN$�-[I���2���lB�1Z��6��⪞���*N�|�x�ㅹ���[C��Sf�-�N1��^���f���=���]*�MP}ɑ�+KV̠dY�91�s3�M�Y����65 ]~yd0|�7�����!�S���q�ܸA�>��I�����g�wb�Ő�G��Z�f�-��F.H���
�N`j��p�r0�E�b� `�7=k/}���N�^�&�gnI�:U��.O)M���_�
����2a�����"&#+��5(s��7L��a�ۈ�hp�2��X:�� >�S�����z�sה�[@��K &��}����et!�҂߄���M��ԏ�Y�n�t*�#�x�<��0���l-{6��M��h�ہNZ!�ζ��Y���8���Y�4x^�\L��ڀp�-�E��S�b6#(�ωd�B�| ���{�f:��W_�������uml��ѭ����R!Z����ȯ��،���9a�P&D�o⣛�J\b�:�aYǄ��ׅ�d�z]&!�0p@M�Qx�pO׆?����r�bH�MTw��H8�V�9��Ȝ�=�cF95�v�0�'1S��u�������ɪ.{��@�Eߪ�!	P����V�!Vq��Kv�ê���@<���Ųg
�iw��l�!xu���vU�E��I�w#�-X��ہL�wu>��M�d*��Fm�+�}d	���,��ٌ�!��O���i�Q����G��8�"���������'�0o�V��>P������-�J���x�p�u�8�S��2��[��<����O��/颺�N��B�v��7^6��7z!S��E���5s�|�����k�������R�>���������0(�r�����)i�ӻ��� Q��ZZq֑�5B<Aܟ�(��.O!�V^r�c���It�g��8/c��q��$[��-��M&�5ם��X7az"�H����Z��`�V4p4Pu�?l�l��QZ�a��)"d���^Y� �Fk�߶֣$<ҕ��c�7�����l/�R�2Y��p���_���^te�ѥ�`�.q����O쌜�� �T�/[����T���������M��@�u���0�s�d/�0�淒/��Gذ��).0������q1�	UK��cҗ7��W�Jb��ߟD�G��nO��o��ɛ�T_�'9���=��?�6V��5�!~��~�4�?�$�9aL�@ 2��q��jp�m���kS���*8�@!?�W�C��ׁ�k\-\�����7�����W�ڢL�X�֟�]�L���^D�.�r3]�$P� �.>?8*�&#vyTlwy��T��c9��2_�T��8�]*%�蔺d���A� �A�=ވ����#[�#�$����	@W0��+���N�N�?�ħ�U�9�:�aQe�
>���o�*K��#�W&��gS�^f�QA�t�d,[!�R:N�1VY��bBV3�9Հ�[�z�!G&fU��R��i�7��7������x���g�1x�!�F�����Vr��:@Md���M5y4�m����z.Yg�K���x���(^�MK�d*>��]g��߰pv�鲵���;}�
e��j������Ĳ��/d4ʕr� Z�@�i��k1��.��󛮼|��,�ٴ�-�����s�<L\p6%��|�3ۣ��za������*K`�MΞ�|�@�.߉?d�<���z]M�������ne��P��ۥnz3:�g�n[@�b�������u����������m���u���K�W� �yAq�dL�;D��V������ഋ�S�3̗P7�"�?K������f��Ln��Bge���,ʘ���}�8�����c�M$�� J$3�{��֡RooM����X�C��}�JP3|�ehr�F�/�VE�r��|PҹT�@[�������O�7p����`��]�����l�M�5�?w(���D�!�2����Ôrƛ,��M'�������<�I�^sӬ;K���E`��n��Ɓ΃q�߫W�p�6��0�ɱ�eَi����շ��s�s�$��gEq6�x�>d�0����z�@�3NՔS)�w�b�M�V[z&~���{~=2��U�9���`���Ed�)�կ3=�í�Kb���H7�̷�e��(�g��i꣩9AE�C���r��br�:�G�
 ��ۡm�gQ��P�_���_uxM�/[WK�<:S���:��� �ˣ�܇
��r�n�;>�]�:�z��H��r��I�^F���K����8��׿#nLl-�Q=�D_t�I�Ln�#{1��U�{�p��LH�x����Z�����z�v�??�Y��%��	۳$�rL�ی�W�k�.��!�:r�_����\����(8����%���ۧ=iy0��\/W'z{5Z�9�-w|��+i�r�i �tG8Mw-w3�i��[��\b�a��P[x1����$P�$!&b�G�}F�q��[��o)>u��d8��d�v�I;�rKæQ�z�Х�#O0*D"C��C�o���?�z�˱*՚W�`Gs��/�9�y�2v[��>1���C�X�� S�[H�����:Cv�
�G\ �W�p�l%b��G��=U��|��%����&�KHy� [�ޕ:#T��,�=��Ad+A�C\A'��[Jո�GM���kuT�����Bo�0s�s�1����lv���0�������jd�k�U��!�|XT�.�ҹu�%3�Ԅ����M�|A��\E�N�X�>i�i�1��r����s[p�E���+��L-@3"�fð��
%��L^'���ӕ�u h9/i���.~-i1�]�����:�z��6ej�f�6y��,�C[�YB��(�J��T��iLScÂ�����գ�a���Z�T_W����{�����!�Nc֥�A�/�8�P���J<��~W�iɪ�[�VD9^*����{ڍ.��y�2�Ӂ��P����/���)��9�>M�����eM�����y��D3J^�I }��"n�;��*�;���k��O�tV�6�b�z=	���-�8$��p�Ƴ�_<E�}[�s灣7�/D��I,��b+�xژ��Ccr������{��+����i����P���ڎ{O���SZ)(��ﴢ2���-�	l\Ô�h��[��kw�ٶ���y-���\r?}��H��
i�����5ʣQE9춴|)Lŏ�Nh�G�π��::4�jW������\cG��|4�4�������Y$c��	�3��a��[ńAm�7�U��C=aVO�R����K9�X$L r+�ű~"�e+[ۥW%������k�`g����z��y��R����>��+��/hԽ�l��Q9�.p�����)�{��x\���;a'I���4�R��U5+��ZX9X�g�8�}��[��E�'�/����6��U�����R>R��W�|��X���Ѳg�6)_��˲s)�h��ҨiQ}��.���%���g��ICX��-D�?�I�};x�����"F/�i�&8JX�W�.W��57����0��5�R�ҊI'JfO
`����A� j?O�秿�z����'��	Ff>q���=�0M(��f��
�����hX ���&�H�}����]'�p�@m��O^E����ە��g�4��đd�qb?A����ę���y4mE���sf�fp��r#�U� �Q����	¡��J�%��7�w[^�r��c�����8]�B|Mr�U���/m��`3��ۺ��p�-wD�� ��4k�p�݋�����w�Hו�!�8b���ȱ�t��?�y�����?��
7-M;}{�p"���x"玻?�S\��K���@Ʉ�'ց︜��ef%|g~�*��^�!����hȕa��6yh-���m�JB~�n��;lBY=я�|Dd�6�q�@(+s�m�`Y�(�������J�����?`��"��2�D�͂y��`��,��:�·p�2|���P���NZ.�SK����K����Ն%	��{�������^�I
����,껽�V�3��Ĳڭ̋21�<Q�B;[Z��[	:��S���%�B7�I�݇�i��/��� 6��v�H�\JR^F3�4Q�D�@�r�-��A�ƕ� �KI�L��1^2�D�B��R+�Zm��>�iM��Ť"w6���O[�^��3���\�'�*�K5�����ҁ����8�C=�"c�02�ødG~�(M%<(9�6�ϡh��'�ln��p��5��5��D�(#W��2d׃���w��� ��'��C���{��[*!�!Y/!��w*�K��tT�ƅ��Fi�C8T��T��`��Bƣ�jR����9_�|>z����X�(����iZ����g� �o@�}�ד�A:�v�hI/�/s��%��h�#�����\2����S�_��=gE��Ǜ8ề ��h�"(�!~��v��N�25e�j�KSg���B�t���r0�r.��,�<�z�F)��Z*��[	,�īx�/�"n�l�o4�r�Z����w볫]�W!���b�8�/Qy��(���*j5�1�O��	��-���0�Y*�����rV!X�Q�����.���_qĽ�sY���A��(g6�r��2P�D6%������J��:�\��>����O�g�暱�@l'���JCP�x/}z�J��	��q'�L�3=���a�._��Y1�ͩʑ�O�`�!/"H�[>!=���_�1�;����\�[�v�.xB����
H��x)�g���f�mb�6�)'d��Fב�B?w�y\B4�=F`��7n���$ e]�x�F�9��&`��95�^�~[D�y�A�nf���ҧ�=Ց"c� �t���8ij	��m��d�P���'��5���I�5:�2��a �#����@"l� ��6�e��L��3!��8P3処<'�< 2	�'ޘ�����m�l0U~���_E�~oO�H)�EQ����B������YAl�)�,����K�֎��jb�\��j,q�5�ή X�Q��J��=���
P-e���P�e���WxM����'>���v������c�;�:Y�z��:\$���|���=���,���įB�)� ��PfKn��W��MIY\ʐW�e�ѿT�p���^�M��fI�R�W���,���.�˕�Z����c)Df�{�]���%^��>���C+�������j�*�:sX?�Z|1WW0:�pD<���e�i�`=}l�V��WI�&I5R=�d�M��Q"�|�}֢����ض�O?� $6a�U�k�=�0wC��J'���n�B�]����/�tu��K1F��y�4�ޅ՟DnhL����0�ɚ�{��~8�9����w����wx�-���l��F��uu�.��gv=��}��Ŷ��L�LPq�Ɩ][п� ���� J��U&�B��n��'sC�������h���gI��Q�� s|i����~�]��^}6��K;���D����;W��z|�țzeD�6؇�|z����?[��EŊ>�´�P߱(�	�����P7���>$�Z��QP�?�:`g�b�����1�v*ۮ\�1A^Re!i���K��hFqn�`�����ܷ��z4�= iJ��"Re�kq>�Cq�F/,r�;�#"��S���^����~*ݚ�=.Kb��
g�<k�'Rl����xZA������e�y��U�5װ���5}�8�=4��q^m�"�Ȝ�$�o�c>���M6����1�������������<�&��7%YL^�[�����ǹL��.�.�^v��/�l,�b�v8�65��°����cr����:�ղP=:��l�ܙYG��K�T'��������j?���`�j:0���� ѻ�}{0�9����Ñ�7O�3��-�G�<���%�����Q"]�S͑a��z$�Lp�i�P��c�_��2NcX�9�x���H��
�g�F�Ĉ{�ЀT(K��
ph;��U���=)�w�����+�t51iC�h|���¥�Y�Ӹ�;������wH`��@dr�����d�`�=��^�F��R�HM9mŊE��Z���PYr��/CH0o�q����#[i��ROIa�8+=(�ޙx����U��r����Kv��\]_'��P�w	��o)8X�z}�`���M�QGS9n�}��\��@��q��U~�C�j{�+35���{���wZ��ꕲJ�Z[c���y.�F"[��ڳ���hHz�+z@�m�*c�0VۊjJ��RK���y�"��^x�p�7�������4AD���k��-���c�H��^�Wt���kNg�4����u㺝(�'ͲVG�:���ʲ䳸�m����z֦��o�߅H]twJ5�4�8���9�g1���75.�N:7͠ ���TL�Ɣ��v��;��%O���zۨ� 0j�t���uYe�WrB劾C��ŕ��02ɍ�LJ-�n�������"�"\:A����$fZ�xh��侶߄��0h&� o���#볏f��k�Ֆ��L�
�eN��R�������q�H���,KTz��LLl�x�ۤ]	גP�-�:P�E���cӑ}���S��՟�*k�$k;VF������*�׬���kKQ���VAv��|���<��K�H�\'�� C+�|:`D j�'�-{�^>�B�[�g5g3I\��nG|z��eț���%҇��"@tC7|�+D�L�	�����"�Z��P(�[�)��k@XO�3��'i�v/�L:}(���ogT�]�UՃmh��#�zK4�߭S�?9U^$�Ƕ��;-*�>��=���F5މ��7���.�?��[~����LƋ4[DZ��jE�D/�����&�S��j�
D����1;l����$/!/�.p���uK��Z���Ym�y���T�Gq�#�m>�h����P��"��Q��2Hyh��eL2l�۹�f�ed;�d���|�g�s����.�r�u�O��l2 ���D�6w�TR5�m�H9Cs�Yn�'7���
%pߝ�N.�a�Z�y�]��.G3���Ʊ��BK��Ҋ�y�Q;d�p��-8������WN��1� :d@�o�I��*�7D�<ګ^j��n[�c�O�eiL������H�".g��ɕ`����iC�VZk�������������3w�ݜ,$���1k�P诬��&�ݖ�Ā�el<����Qn��9�	�n&�T�%��D�	PR�� ��G����,5s�L3��<^|ZM�veԬV%�c��2�0�jY8�h/�T�T�0�}tVvEUqR�m�~Ҿ�&��NרQi�������VFb��C�R��;��y15���u������,�x�C�V�~Z$�7nL!P-�) ۯ���yA-���x���-�=����&�р�u:.[����i&dj�b"�^]�N�V#�4D*�_�(Pv2�ð�E_�7[4�3*�t�ig�)�3~"7$S��i���[��p��� �+a��5C��Qf��k ��4X^/?R�����ӊ���eNn2C~�mi"������_k�U��!ŕؚ��M�$'B�F���+l��"�?$ۓ�]�M�[�v��Xu Z}$��d@2��a2oP~�%�P�7p�b��:��"�{�rC�c����SSx����#�B��;�$�z Y��Zav�7�t2M2�*X�5�j���ѓt�`�������4��)�?�=t����d��ϗ4�m����n��DRn��(�i�%N�����'s��ɝ{�|�6��Dxˢ�6��˨b���v��^��e�xé��z����yA�}�2�(98�~�����\w�g��#�Z�s�w�TIX(y��v~RR>xf�r䃛�(>�"��7�CB3#�nv�Hr��+�U��6����3Q.�׮����u��,,}^�l��Ɔc�T��� �ǈ㓀^��i~�5�� )+Zہ������� `��5�Y����-��=]eFn�r�
�\�q\k�B' k�ZC�"N6��������@hVq�a�����-�2E(�%�
�Ph,މ���T���M5t�6sJ����+����ú�zX����Ԣ\Q����*p��t5��Z�O����mQ�6?��>��s���T��/;����rQ�#�4"���Ճ�����h�|�'�͎��H�k���ߕ��e�`̎p��-a�H�j����j�R�q���"+Q�cz��7 $%��癁�ɼ�_���պ�)e0�����m~��iT��Imm_F�`s<��E|�!��H�n������O����)QO9d���%FQ}6g�
�V^&�;�a����<��Փ*�l��@�D�|E���]��}�Nix�Yo�O[@X�p���	��7���(0:���6�W�j�����x�F�<�6�8��:l�Ў�:*�p��(��FA����vpl�9�?8�ם���8������(K�����w��܁�Cl�-�Gf��L4D�+/S#��#�lg����s�1-� �K�k(:�h�X�j"]����pi_����F?հ
/�j�i�*�C�:�E2}.����0ey�a\F�CN�Yp߲��$�V�t��h�!L<!_��4�	X������z���~a8aģ�1!}�Ru웍��7e�$��V�S�r�T�)ZE��y	
%M���̐�*5\���u��tH���	�^�7�r���Q�S�d5����p^s	���\��	�[@�}�e���\��/?�|ϜAh��O��2?�)%J�\��-QJi��К.ٿ �gd�9b���a�7V��D�!Y�w�o<���{G��6����u1�b�/dL�6��E��մ,����I,B�G�^a���k��z$�M�BP;(M֓���]r�"����76h�Z唹�ܦ@9�x�5U'ոxRScN�'en]9�kuS�]�I���߈�<�mW�hGW�uL���\��5P!�CK+���=���Ѯ��w8�Z����L��Ҹ��	W�nX�K��@|!�i���}c��N4�Dh��#����C���T��p�diAxկ_ K�<�����u�����3���M����6��:���ϗh��{�z�Oa(�
en�Re�R��'��A�a��5�b��}�b*�s��^���r^�[���n�� e"F�q�̝��L��݅ �M�n�2�К�~=8@�'m�ӘP]�|��;�4��4��T��&5a�X	�?��?��
����i$[��:9x1��q���nJ��Yڇ�ϛ�j�����	��Az�N�@
�oAۜHv���}2IԒ�S01"|F�[gn��a:R/&l�|I�+���Z�Q0�Lؑ�Շ>�KI�D2d��W
`������$���B[p	��;ՌI��/x@Q�2�J�5y����읛Dy]2F{�ɺ����w�5��ߒ[�~�~���j�K�z\�����\��8Kp`?�:X�J��\,�)K[[<�QN��2�~�q��A����n,�7R���ź�)"���'P��A�N��T�u�1]���Z����L��r�-&�\����6$���&	��Im0m�C%��5-=��x&6��O�63�@l�X���k�2�⻨��@�����V7:�&��	@�P��k���&��ߢ��lZSe�e����ش��Z���|����S�e���' ���K���bcA?�A�('.�~b������� %.)���҃�(�:�WB�2^fa?���C��ؐ�F�i��y�Z�6R�k{�'>�3��L��r��I���X��+$/�l	�Ʌ�J	��W&U=�9�b�ɴ'��b):��x�~@�����)�T.��m=�J
�zޅ���fa*rp��>�����y`
h6���Z��@����kf,$��������e��7s����('����e�`��CB���d1�p�K(]���ޓ�ho���L�'a��}G0eD������-� 
�!u[M���������Lʽ�P�Q��O|q7�0W�@�������x�4��_^@�0����F�MB#zo�L�R%����]�Ԥ;h[cBt��j,θ�|��ˡG��T�)?�,o�}Cgyd�&b.T&��jT�����=3���z�U[�Nb%#����Id/r��(M����f("^/�ڨ�[P�I��M>n��7��l�1�k[���=��G?��OV.E4����8�v�{��YG�-�gk�}�!./�չ��}����.�@�Ԙ'��3�[ �j�7�*?����������n��|\b�#�7����}QC�Q{�H+*D��Pw�f:K�5�Y�`��$U�R�\��ڤ2�%Z��n����
ӛ��jn�u�<�l��"�A�{�c>���@���:���8�K3�K`���.�P�CVz�� ��%��$;�1d����b�u�-ס\�����%���������e�P��'���*�̗�T�v���X�l��5{�a�u���[<���� �����a鑟_��r�z����6�����П&�K���Vpfh��:�Z�)"��Ș�j�q��}MpiT/I�t1�U�i��A,w��"���PD��U o�#	�`���ݟ�Fb�QA��t�����w��iS,�m�*���1��o1�N+�v����8(	���N?�^�b�����{��|g�����3���u;d6���̌HH�"��b��V�Ab4x�]đhC�~2+4��ɴCxêVb�o.	Z�T��u?=>��&%�������=1�WM&`��j�-�L���"u�8�~��*�ה>2�Si�����TJf5�E��p��1!I��=�b-�hy��O�Ɣm%o��i;�*��x3�et�nR�`�U���C��bCc �U�&n�r���6�;����s	T�:~��X��|����x���6u�:L8!5��E֣�00�E��|R�����3�	��.�&.�#�z�P�M�����f��	U�n0L�#���_�����Ӏ61��y�]%N�>e��KqK'� �%E�g �7�u�};tn:����E�sp��̺���mi-Jpt`A"E���a�(k��+�ޚ���������d;�3�#PB�-��Q�`鋕઎GiO�)F�hg}���lͫ?U�g��7�T�	�2�Y��~ �(p-'�4�p�_����d���A!Z���z@p�k��L��w��0����\Y�Ef�6%��N%>l�Gl�N��f-wx(���b��M.���G{�2��`Z}T !���Ë����B�/O���ݏ-��&��[�	9䪖-	��QVwl~�Al���߾�boN�Q�	ή���A���l�\P�6tD�(.�`�ԧ���/a�cyN���D�^)Y<�q8�YIH�̿<U�ylJb��q�j2�*6�Fo�2**9��"r����+�}�8��`U�ҋO	�'�F���TK�4���r$G��l<�c �q��b���d�P����n n��3��)J7�[&I�C�O�R�?��k�LZ7�aN6k-��WCAm d���������s̻Ϲ	F)H��C�Z�p'�Wx����_:��7H��B�\G���A-f75W����р�¬�q!�Q�86�m:�i�H�}�:�e_�״�jW�ԸZ����ON�i�C�D��w�����W�֩0
��}t"�}���ǲ�j.�'kc�]�r����.瀔/�80Kt!��Sl�K���1���]�iȴ��i�q�@�c�@m���	g9R�pl�X��A�5n ܬ��9H��y�����ԭ�*u|L�*�=͌�Y��r̯�%�!h\W6	y���ݩs��\���<�~3�N���e;�6��U]��Lb�>�g����ŧ�Y��C���̂KܐA���c�����6m���fA���q��ʙ��Sx�<��[��6 >O�/L��s�u�Le��Z�@�҆m_S���911M�'Ĭ¿�]tE �>>�b��!̵���?�z��2~X�{v���V��S��Pzs�.�ѥO��+�����}I�����fc����Zo���;
�^&���������[~;�9��R�?�q�xu8� �ee�e�p�a0�׺���/���bi�-��������u,�mP���B�#.�E�� ���k�������m�I�'q���J�W��r���>�9���ƣ�/����c2�=��0�F&��Z�2S+1�N�*էq��[��$��h�6������o�Փ����Q"6̝�0ߞf;@M�\/��?�ǆ�8�\�Z�'"<�O�����Ӓ�O����O�+�����r/&�ñS7�����A���x0(*�22��GI&�}�C=���t�)�3H���BR ��Í����!���&t4ǱO���mBrdK��O�V#�+�5q�{��é
z`����Q�\6
�[�n����6&ѝ�!��n��5^��S>�a����`.
SF���H��� �mֻ֢�ij�@�ժJ���5b�D0�+�Ү$�s?>=��)��7WEfK�?���i1t�;�6IqVs��&��D"�H���c4�����~q�X�nY��4�;���F�p�;��%�d��{%>�;�������@>��M�)�p 8z���?@�'B>�,��g�}F�H��ޏfZ�H�Wx��q�x�D���d2Z�����X9�f��R����`�Ĳ%�������D��*�&5��V":we�(�f�0�C(vM�� �
$O{V;'�
��g-rIzq?���g�8Ê��{��t!��n�^����fxj�~�!�����if��W�[�]�g�H�s,�ܧz�4]�g�O{�E�#ⴓ�����8�5��vn����~�c��ι��BO�F�)��W�YX0��L���S6�vI������ԯ��d�������?7r�!�|����}%4�lN��(�p�P�g��ﲇ����{�aĉ����|R�E$���7�܃�,
��V��&�_���hª���s�����j�S( ����]�X�|d�s�bm���}s(}���VϘjGڊ�� _K!� ��P�
�M�����i��y�Zd��t�'|�2��ɾ��r��v�Z��r\��|��L~9��i�h.��g�8f�<5�`��g�Ϊ�u���A�t�|�A{f�ze%�.WB��c�b0�����E&�u�k�r{3�z�j��(Is����Ɛ�����-�D�.���<��N����9g賨��:h� 
�5"=��JM��"{���N6�?z���&œd�_S�+9l2����)��Z��J[�4z �1�b��$.0@�2v���J�l�=i\�뽒R������.@��&J���ӫ��Τ�M��W�x�,�P�'w�%�I>T1�<�`#������U����.D�K}�9�P���^UQאK�cK�U+ P�`��A�!P��2M�Zm�[��uE&���:��CBƙϸ'䜓m,�&��߅�&@5����@�4��w��C��ö͙�ן�2c��T��U����|��`�ޝ��"e�ݍ��6��v$�����ϒ��jlr����J�)\ �0�
2�o���SC	���y)�L�S[�Z�;Q�/��ס�+6ΰ��j�;^��O�y������p���L(����ۃ���ld���LSDy!񽓵��c�!�;z���@8=:�q�?q���Q
"ޭ׉�֠av�R�q����G$2�DVA�� p���:#�%eD��B��1��y���w���[��#'�,��M���,�`U{�4W�'J�2b\�9��L�@�s��?��2plW�'a��6�ӿ:t����x�.2�V��5��}��Ezur��қ���[��֚^��U)�F@2|7��'��t��_X�m~z��OV�4U����n���좏��%����Z� n#3�W��Z��X��P�X,�g��s��]9�V�r�����,j0H!�4�G��:�����燐zU�~���� =����*����d�� �T��1<�^ߌ��)tJ���r�����|��Z���d!��ZX����<��j���)�����ٴ��#T�~]$�nI�O����j6�zI���Ԉ}s�Z�<镔�����c]��h�f��0ǧ��K�H�JƎ�{t0rv2�M��8�(�Y�Ç�76�/��̃����v����1Of��H<����|�i��'#���`���:��y�'�G��yMJ��`�v�(��D2��h�nO�����贋��A�_��P�����N��E����_2X��w�礠>	��'��Ns0U�g�,���_S>�+6؟�Go�Zn�flR����r��� ��O8��YL�v�8�H�C���6l� ^��ܷpb�0c_s��$�;S��T+J�k:_�g���ń��P�GN��o
�R��j���+*b��$���B�s�E� ��>��%�"�2�
w

�N�m�[ڱD6JF��Ϋ�����CW�E��v#��0Vy�־y`@�Vyا��\�/�
��y9Vp6�A��B��ῇw�X�7]].E��D�l�AkI��!Sb��ۥ��cB��`�,�k��W��74}F<l���[=�u8�ƣ����^\@��T�:�x�i���l�͑�^�<��)Q��^�S�>��0FMZpc�ֶ�n����I�%�`k�hm�� +�͔�~���f�Z���LEf��?p�i��u'ʸ9��W嵻V�7�+�)m �����1�d�b�n���b��B=s6��3��� �%[�;�E��Q��ȪrS/"3�|v�*sJ�ݶ$�3�VLO�������2���U^���v�:�P������4����N�읤�f�^NH�Z<���k?��|CSE7228��{���^�#�젒㱉{�jGF`�I\�8����d� d�P�h"��*n�,Sy�)Et���9�m���GRk��Uг��h ���2,ܭ�3 ��t~I�[q��1�����M@��E_r���[�$@�0,{��_|�D���c��Z�#g+�B.�J���ӱ��E�E����sG�o��<Q�PW�T1�jjg�e��b���)��ӣ���8@X5���"$��q�\ت˙x�i�斧��0i8ٗ�^m��^��	7b�:|�`�x���)Wy��TXܼ�*>3�Oh�g�p{��j����$t�!j�����I;�S�IA��#/�IǴ�ΌV�8&B/�����=���k8 �ש�x畈.�� -3N�KGHQ�R�0_����d�ٳ���m"��U���3�K�.`���Y���q3.���f��#�&�q�;���?X����MY�KAE�D��rV��5&N%����d.��	�p���'�Y���c�?���k�~���9�ӄ5B
�WsZ`�����D=�����;+���4�t���97i�=�*�<G� ���L�\�f�yeQj�!�T�-��z��y n����_?�/�>�j����ܐ��(>P0��ӰK�d�SĨn#3���ϊ+��������h��+p���`� ���w�l���m��qq�v�l�趻�?���G_Λ:�M�a��Q<w�I&AX�&
eeQv7�s�yT�r����4�Uc�MҾ��qB��o��k��*&U�ܴ�g ϕ��RgB�y�Mi�.Ā����oD0��Z�ܜ����E���k�
��� 1���x��qt�/
J�Q��b�-��Δ=�>�ȯZ�Ki�}*믕��?x4O���^��Y���n�6�%�Bu��]qO:����Fo'�)���W�s�B�էra���7�
�>�a�+
�6a7�ECnܪ��y!��/%-���߉�"���/���gx����Hp�?���@�k[2iŲ:m���Xh���F�����J.�d�1�Y��M�y�q\x�;U[�E:R�A���)+��Y��o�7N+�~=�Fh��d92����`d����U1�(����Dƍ�H`s�LX���ʆ��چu�>9�"�B{��Q!,���(��L�]D�D�E`&JJj�}�����e���k���� ͢L�(�_�	�| $�[��{_����{��ѹQ.ߛsm�sv�P��c>�Y4�F@���Q&���iv��i|3,�EYb��}>-�5-�i]���&F��Ύ� �3K��U��A���)�NKq��]W�r��,��gJM�j�r�a��h'�Gtd���sF�a�CqcN1=ey�M�a����xs��)����4ZO)������P�8��������"ϖ�j����󏩗��s�r
(]��aO�<�1)�A�b�T��d�f��q%P�.g��]h_F��4�֎)_�^@�V�w�y�mnrP�T����6ڧ����u8o)1�3��vFBv=/U����g]�R������R4v���u�S1D�;�k"�g��E�,��B�A0
��ݦZ
��CY�5��噏����*�D`+]NќA�e6u_7���+��J=Y\֚�f[+�i��wV���H�	�R��*���9��Π`:F��Kd�G�h�V�y�#�uT@W�#��>��8�K�|wF
��=-G��k1JYk��-g;Vg����2�(��6����U\2���d�	]�)�*�k�k�r���49N ��[�*tb�=����vK��V��דʉ�s�nG �װ2e�OXo�7�L�M}uZn͐�qxW��¤o���-�C�:	�GI�z�VvC�d:��-��Z���ʴ8(��2���y��3��I>��#Y��j��Ӄ�����y��	�Jl]ӱg����䓫�! �����^Źhg=�A�J!��h�?��q0�j/W4�7���V,X%*6ce���C��{�d��A�J��Y����Y?����V,ì�Z1��.`v/jh�ͧi�3��[=���1�Ϩ��F�*���:�KEс���yS$���Ml�ׅ��J?�ÎN4Q��9nZ'�I�p)�-�)E2���P3/�X_^�1�7v����{�W���A�6Yz�����g�(�,��H��F�ۭR$���g���O�'��G���l�2����㷑;�"!9,%g��!ؽ�1E�[�Dv0�-��F��_���R���B@��2�4_A����m��,����l��&�|��J��┗��i����w蕊FuY���q�3�ބH:��06�X3�/p��:�D�iQ��A�>/�7�鵄l3��e���9�Fv�D44�S�Ñz՝��N4�Hi}B�	�������~W��<���RoG�Րz��Y�'�� w��^V#	����k���'?Iz��lvi�Qz�Op]+���P٦��!%(�)5XXD�M΅=~	���y�����i��"�S�&M��@����4t��U���]�el^�Yw����E�܇�i��
ɡJwn�%���R1�l��e�oM�f�_��tCl�]�ٔ�����Q|�$�����2�4?�g��j�-�z�P�%�ԑ~�+t���.HJ�.T�f)���a 
�k�+Qqd�=慶���]�r�щ.
��/ߟm.W�᪼-k�Ѯh�F��>Y�ȗ��eU�4��֨��&+�E�&X��Oy�3�'���ӎpF�_��~$!�D5_DeuO�X���ADD��������ֵ �3�y؉weC���sT_�����r�&�D�_V~տ�Lr)Y���I�<���N�dgn6���x�7h=�6Eh�I!�'@Z��+N17pm�Ra2�<�d�"�4��aOSMI��H�K�P����7�s�����7�����ד�r�-�ܜ���E�h�X����(� b�դ%�,z������,���x�(�#W��?�txc�գ���߿��ɦdu�x��d1�?&�Ks� @�&��+���.f�����],��Y��C��mڬC�\���GE,DY�O����$H�)�C��v�BM���z�{C�,��|�2���%9�v��]�Tړ�L���)�Qo��]�:qT7��`'(M��ߤ��Z ���=�: ���B�%+�ک^"ͼ%B9e�Ⓜ"�4Q�������Jq����0��s�	�
uѵG������NF#Ũ���P���� E�c�#-���9�M]u�w*�����~Q�����a�Wu��9�/�F̽^��NYS�~���v�1]�o����]뎽=,rruI37��rx~'��B�-8{쿥���05��N�ޓ�y�y�u_Л�̹�ʙbj��Ӳ&�4rE>�I��:��,�� �fƳL$d�z�rݓ�[x��9��C�ͨ|����#lZ:	�s��IL�l�Q�3�Q@��p:5cPơXT *4�}���m��w�	��ᕧ���e��L�c+�����l���n��:�5���QX��$����e�R�̄,u�c1��	�Pah���]E|3 ���W��AE�1���]��2�m2U�L�q|��C����f;2�C�����s�f9n�Z�D���C����Ml a����GN �c~���񄹆�Q�1H�S�KZ:[F{��Z̄ѫ��nt�8�4,��z�=,��%d������)�sH>zB�r��xY-G�i戻 �N�J���:٧��������n��P�܄�7�J\i{R񦭨W��½�u9�V��(DR�kJ��S �IgX��ψ����~U��s�<��|��V��8k�RgP������y�]�|�4(3���˂��{]z�?�B?��(#��$�b�jZ�������-�L�G�g�77�c	��$o`�\H�}�t�J
���lR][9`s|��	n��_��ZN	}�yb(�
�2v��0)�J����"���o�Ψ��^�mmx[��P�z:���K�\p���W^�V�k�(>N��}"��_@��]*�H�MLcf�tRWLIϻ׶�_+vA've����_��x\���J�]��'#�VO<�PGN��=���^!+3��z�:i��!@A�'�e��j;5l� �aӄ��Q&)HƢ��G�|V'QZC[��"��犞��z��.^���I/~��h������9)kݨw�_9��G����#{B�կ��zKa�5���V^�^9K�t���]�:M���ͳ#{�C��@Wd4����8�+��q�@9����}vIuU�� ����5�QS*�w��b��/���MVʐ�_n�m�O͸*J-aXr�L,S,�d݊>{�5+c^yi�T��(;(!�+�.��ǉ�;,��G߬<���7�Z1�I*�dX���L��ȱ��s>�3��Q����
tY��'����D�Z�P�����ӭ�zro<���q7M9H�x�5��=@!��oX1���e{n�Qqwd���ls�1����ߘ =7^E��sѹ��x9$���fu6}n0Sx�h�ɚ��p[�im��<_��/�V��Ȝ�N�F�Q?%�D?-�%�H���Vco��׮��/�=Ӵx�Gh�uo^��|�Z�J�_�U�W%n�8�����:H8�M�9��� �$8�ۋ�D�MS���i8l�1%ΐ�]�n8���ɬEA�1Ӗd���	w��X�d�m�Ն���
�3����,��##�?D��ѺC��U��E�1�oҘ�L��.d�n��I�iX��{~g�:�m����{ C�������%�lO^��S#K�k�	,�LV	r@�%���Xn?	(x��*x,�=�N�jN����xF���}���V�c�*1X�B-�I6��3=�@Uk������/mmk���m��	���ږ�jo��+�Z�&~T@�C��Py%��R��ӄ䨍 !���#�n"vG�4��o���f�Ϛ9�5!Xݨ=H�!�s��xs_��+aS� �����ʑ�e7L߯Sk����b��Gc���顫R����%�ÀEə��~V�KQՖ2�]?�٭�J�#Ț�(SM,�yT@�.�Vl6��ޓ>�-(~�����ER4F��7
�I��z79x
��!Q�i�^�T�v,�@��;�O4�P�

�q o|���2�v�4����%s���-�G}]�E��'ЮN���w��%�����]���b"�M唬����}�sp�,||��//��C�u�*',������L'�ͯ�}�'�����o��8�4�w�}w�"�~���tPJά9��m��>�c����D�F�ԏ�]�ڵ��Gʩ���U�<.�f���V�:���C[����d,3��U?��)@bx���歯A��o���b3��S�ӕ��k��  �����P63��A��/��r"��]n���^��n�r�1v���8
����
�ZtQ�.7.����.�4{ g��x|Ko��/�(v�#,���o�
�5ٙ@�H��� ����}'�_��.<�6�t�
�(T`��}Ƚ�y�j��#�Uܖa2�ȉْ���x������t�߹%y*�D��b��Z��D[�~�O��>�L�Ňʮ e���u Q�w������P0�8���OO7�	���q5���5�Y�'@������u���>���G8fq�����[���B*9�Ή�;{]L���`�\����(��2�|/�����H�=�(&B?V�{����v^�/��"�R�X�, յ;��2#��a{"�qE���jՠH4�NP%���TID�|
��w?�#Z��f�T���9��x�Kj��܊6 �;g�'��C�VO�^�`�w|��lб�5͌ �
G��(%_|��U�:��B�e��d�͍�X�¼���	�R|�ip^�\-����V`)G12���ʷ��>i&ZBbL�x�j;d��%@�B��"<2 ��
�X��^$Pz/W��]�k��=�%�W��e�oJ��-�"���`5�j���龇Ŝ8b��V���ܑۈ�}��"�ԌR�Sd�}���4���աȱ[0��[�ax�go÷4��U��3�`�_ȡߥ�`�`a�"��}!�/G'jn��Ԛ����R)�L��<����*!)�p
%��"�[���4lu����pS�d6Y^t��&��@x�_%�}� z�S�TnO��r=�g������?���������۶�]|Ÿ��8Y�r�ص��	y�I� �����ug�*���'�i�ȋ����q�֢JwW֑���ߊ�h>�nҫXGn4/�;�����)�c�8�D�+����oi�y7�%)�����=��q~D��C^\�8���_�պC!�X�k��~�BIR.�[����ܾ6=�� аZrM��}
��|�M����@j���jbP���w�� ���O�ҏͳܱJ�L��Z�m II����q����QB�V�p�U @"�}YF��)�0Y��M�B�beW�9���	�H�'P��L��=Z�,���v K��TW� "/���Ђ&�b�gڻM�y�u�	�o脟)���wg%�;�m�����&PX�vl<��&$&�.��'���'�����n�t�cQk/%���pf�*��p n�mBf7\O����}nZ�s!4jY��q�,.t#t����b�S^��_i�l�kW.��6����x;���.\�_�����X����Ip���qݻ����c�褥x�1�a�:���&�䷱/��__)�^��2E�>qh�
���!������W 9y��e��/��qcfL:��8��Q���nj4Q��?�t�s^p>�M!��Am�g@�6����_���*�݄\+ i��I/�tm����)�	ľհBm��<� (��1�{�_���i��L���X޵��쫟R+�C{�'b:ӇQ,�=���:��J9��ɢ��'e�+W������e|]�ơ�8��E(1�\�z���[᪥��3�ߓI�O<</�0���m�/L�tY��ﴥr0�b�œ�h�	��`f����@Y.�r�q��FQ�S�kN/�1�(F�ɘ�v����7c��k���;�ߡhf���;���u,#�吟i�����|-�|�f���7���өuU����KC�*G��Sg ڰR\��
�3��-��X���.�\�dj6�����־wb<��z�T0��@�������I�/2"�w�E�a��V�Z�k쥄�mU}6ߘk���.ڗ;D�O	��B��\�������n����Ci
��������$"�F��������w<��B�x�����`��58��@�sF�o�Pn؜��xz��LW����<(Щ������	]E9#mR��;Wn1��F�o��o�.G�2�B�~,�h/T�����.�3�>Z��;���.}��l+��1��;�Ht�[o��8���@MlB�"���}���v�F����%��N̊�+�q7��k@>�CK���
b'�n6�zњ���k�8�ل��y>P���I� �l��o?��QKw]��2�M��ݦ�#�N����(n[��#`�EY^Z:�J��_������|+�H��P���TR\���4��`k.[~p�g[�Gf�1_���c7j֒1��ŷ���eJ	�.5�.KB�=9�kz(����R���l��)I���,�b�~/�rݺW�l�b9-�Kl��o��sf���ks����`~uW�,&��΋�+mk�_;(�&3
�|M��g<ĉ\���5F/��I'���?˟�W��2� �M˜l�H��oX��uV�K·[�+��1�L�p�%�$<�~�!0`�к����%9��Zl�<Ƹ��>c��@T�m��1�?+�&P�R��L��c4S����L*?M�0B��<�E�Q�W����)�>�LC�M���Ey�O�� �v|�/�o�!Ge"ˣ;E��X�_aK�޿���/e�G��g��}yJqT�>yq�E��#�{mX�s$~	F�t���Ȃ�}�y��m���f�O��8�JI"t-n"ɽ�lq;�	�_d4j ^Z�"-��Q˄���w�)���?�G�'M.����"G� ��v�idk�D�{iMڄ�K���6q�=:�\���@%�دK�Z;@eL!�7��q5՝��~B�ad�t�
�9`(��ʦ�S���P� �{Kxy���$�	�f7��3�`�Cd�����8�g,�8��!�����庢�)1�g��!����(��ӗ+qSt�Ͳz�sǫ�_	��ʪ�1V��xZ` ��S��r7o5T�q�DuN< +��GY�-�=���d�O���X�g_̏�2%�\��s��\�Ė��`=`W��Fnְ��l�[Ad��V����"�7'K�O�)!s �`9{w��~�ڋ�����M���Y?P�`N�;~ج��+0M��@~o��t�ė:	�22��V�f�X6�>��:����[���ߗi,u��d���/!���ϼ��� �b�GS�M�*���VQ(����[{�`[���3���6I���YG���A��Q`������/���ݤC����{~���{�5��Ke���y��w<6���H���_=v'8Ͳ/�Ǩt��*���}��H~��GʩJ9���Zz��S�jTK�����|W��B�mTe�i���ǻ��� #.�����OP�m�mƨ������/�f��+��WW��Ʉެq�ko��JA�w|-��<K	`8/!���XN�4n�)�u�9:&�s�w3�<rB�|�q?6^F�e<O�:�yq�[:k���$��@䔱�U�4�i�CW� ��n�tUp(P<ٗ)�H��}/��ݥd;c�\HSt��7r��-����frS4=m�W���2�e����$�[��%a�!:X��n8KC�WM^ḱ�"}Hf\%X�4�b-�H��V1�H C]���~nSqv�g�dS)f�t�?�V������L,L���`���
���C�kǩ��8L��2�а!��H�IRۖ��K�d�����L��&`TQ"��W��9�sp��7ȚO�9��ԑ��T�4��ʂG�#["��{�1ɖ� Bq��$ۻ���,���{�,����3C���!�J�Q��~Za���Z��t�t�v,��$����;:<�Kϖ�`/��]�7����L��uf�G����L1so��'�w.�P�~�5=lW��.��:�xh4��F��x�F=گ2@q��ع\�|O��hK{��ى[���'��.o㚂�=j"���':�ϩ�Q��F�(.}兓m�L�2'�q��_A���x�8��:�_�|���B�r����n�g�6�b܌��p��h7��C� �Z4|Dbș�!I���.���<i�BrY={��'�_����b)�G@�L�.�+4�Q���[ ������ςrF8�Z]�'m�ZmA����uS�%���K׊�ň�L�63��A*)�E��U�<�6T;�$cɦ t�����ȭ��L�zØ�� ��U�(��4��U�-N�^1�~���-���df���'���\��}�3�F�x���� 8(�ȉ�폭i�b�����2�-����3b�~�|��v�&�����:c&�\nc�+��'�8��1	�E�Yh�,?�h�5���,����=���N�����@JvEuN�AE�Ռ����P�hz����x=NK��z��U��bE���q��::q)'�<"D@��U��|������1:�����j8�Um�4r�c�!���j)��j�5��f��P���.E+O��!G$���#��yǟN�� b � ��j;K�r+��i703@��4L�rB|0D���1��OVY<�����q�m�36�h\ό/�:8�
�L��F�����R��MW��%x>%��f%�g�m���v暪�[�}~o7�I�U�^x�|F��8�'V�v��aO:�gӭ����%V�nI^��"��yK�VyN\��L+n#w�E^��%�������bQ*S}�w�hb_mCqY�L.�C��LZ�`x�pNf�!��b�gEcA9�3hj�J��ij��QV�<��c��(=����x1��<��8��a�g1�C>�(��޳����9Le(��e'�A�M�m��h/�Y�oؓP�;����I�����5��y�M��ػ>t����	��{�|���}q˴LI75^�e�l��@�
�����c�y��9ܽ�v��V]_�|	�#=�C@����]��`#���@\M,�$��P�b5w[C������^��r��2�6mtl/���|6Y^�")�������1�xK��8�<�b b���8
I�5��֤kK����Ժ�#W D᰾	G���6̄���{���u�!�Q�֝�f/�At����_4��J���4F���]~���MH>�jw��j�O��bz=OW|�ُV�R���Zc�o�l�Ζ�-��s��F�?c-�~W�N��Y��'���bƲ����������.@���ׅ�wȋH�CjB���_�::ع.�l^^�`u_�~�꫍l_�B�B}
�{)��oK 7����O�(QZ�*q��N`D�*N<P0w�)�/���N�Ày�N���G��[���?�{�����$���#��_ʺ1�g���BQ���N�x�����w�VD�U�2������fx�%�8x7f7/`�o�.	FP��9]D]h%�gT>�˕��a����,;%E�)���y���gTl�`���vk4�A�}��E]�n���O#��pN=���� Cﺧl��r�&��턄˅M��=��fa���j���W��t��Z�[�8,W[�p�KB3!f��L�#�����"m�,eY�3��{�� Q~�J<���n���5�)�c �w6���C�xI�bÏ�V4t:����i�d�oO�a�W+�_֒�SW!03��T����u�'�ʣb˅]�5�-�����HQ3���R�<x��9�Z}az�'J@j����,"nxo�3���MQ~(��;xϊhU3g���&�j��m�_C u2���?��\�1�,���s �-�w�piC��%q��~{���ls��C6Xr�vv�ڐL%W��W�[-1<�2,~B�)���$��cG^X��~팥t�@9�2��_�s?(�\<&<�\��?����Ƴ�l�!��K�]���`v	F.�ֶ��#����It^���bQ������,l)/�B#�~(\�$�d�%)��r�{Q�NB����۫�#C�~R~�Su�AU�| �3��Zm5E�pS���Ŀ��T���m�V#��@�У-����|�.�P4j:2ĳ�ȡ����ե����E!��1�1�0��*�獯&%�ۚ����/BZX� aK�W��W�j��9�٭�mm�ʑ	t���qQ˒n2#[�DpA{�e�,��z�ׯ4��!�}�]����#[7��|�)P���*��L���?�
?V5�r���l�?ĦV�-� �qx[J�b4v����:�|��k6��#�b6U/��ߜ`jP9��=Wc�_SB9<+���<����K�N�B`t�5�&���k�]^/��1U�nO�E�����c 5��"Յ+�'���g�@"���}�/t�����5�%�n;Z�8Zڱ#��N2Zi��èW ;��;��G\�c��i�O���W�(V�� Ѳ�����e�W�9�6d�p_7bT���}ඝ��spR_�PE��ٜ�g9A�:#�i�- ���݄:�)2���`ޛ*e~�|�ט�T�h-�6�AhE"�~�>��J��<I=IS�L.�;����th��ƉU�G;�����bRN�^Q��Cmݬƽ6�??h���6ZJ_���a��f��?�}�u �k�y��HM\���W 
Z����8�(�G,�̈́bV5�%��n]���
.�s��FV8��_}��ei��`�B�Wky�
�!]�,�>�f<Iۆ��bdX��
�noQx��K�\��ޤ0@� ٛ��+������,��D-$��-ѓ���|���*tV'�}RߠB��^� �����a���O��0io�ݘ�Ti(<+�X	�v���pVRX�B�NEL!>d|:C��J�G��y9� ��%�*L4���m��F��EKM���r0/	2���؛mzv���.�׃�=&�"� B��f��U$n=�>��v��5�E"�T��`T��F� mP����0'z;�/'Na�(���\�g�p�A5�a�p��Pl���\�J���h����G�+c��ͮ�3���s��+�2��:������0Ԅ���T��<�G?�Pm���okr~���'��g�k��i�H`9��b7����B/~��l��b���w�	���)�����F  ��@1��{De���9*��V���i�rK�F��Yw�73�`*C�魡D)��U�/r��t(���]Ҡ�9� Lq��[��kg脔�/�HIY����CL�V-o|"*��0��� ��S�n��v�:�;f&�}'`��l�ġ�m��_C�������x��.��cH!�O$���f����W��?�k&M�|	��bt��f��cpk���%���5f�Npߔl8o���rY�_��,'�ܘtĹ|����w�[���a�(�����Ί�廅\L��@�����@�v�,*�CV�B�k��vG�-Ͷ���b�Z���r*��wg�e��G�U^ސWMGvDw��턡=�m��"L��<���wy���4a͓��������ڒ�D��P�mqI�I��o�5>vI"�_�F���5�k�4yaG8?�Эó{"�)M���.v�J�ڢ?\�3�м�w!��~9���'�UD�p�76��{$ă?�߸A�)���ScɄs4�n���H�7�ФoG$Ӌ�����ʂq8�<�On�?7�r�#+4��ՈvU���y����Q�J �h��CP��[eV�*�2�d��XlE�W�O+R��`�H�>5�Ʃd��G�)��o4�	a%�_K��L����M2rm�e;۸�5�4#I�j��B$ި3k&��U��R�^|�7�v4]�Ȁ'���'jL�x���ٛh�D���B��OO���zi=�c�	%��#|�	���N�m�N��H��E��x{)}e
Р}�z�1��it� V�H#�j�>�� ���������K���:<h��v S*'ܲ��-��p����r6}%g�z/�liAfWH��,9S�r����ʹ���`���+dAkV����*�0�ED�O�Af+�-�iS�o�Y�d�k�Z-����@:�)��T�n�KPdt^�|U�ܸ\/�1� ���1��(���QteY]8D��1X�b�02�!�$ַw�m�`Eg��������P�dg��4:Ɛfn���6���e�Q��s�X�Y[�iī"���H�+��^=���8a
$���A�l����{&U���@3�� �ôh$�߇���9�D�	�V%�P�Ȕ'��Ƭ3pYO&�7,,��Ӟ�2<�@fΔEZ2��|��z��\l3hoE
�ō`�1��f�}^+�*R[_��^Du͏�Hy�J��ߊ�+2�/�dkv�t-3Ղ!?��ť�&�
���ٜ?�����\�aJ�M�ZL���!<'�O�VB���ڪ�bh��9��U[킉�J�6m�m~z�JwLl@q��ϱ���5r��<�[�TL��J#>`N�kv���@�3���MW}��y�Ё)��DOrU֌��S��pO�һ	\B7zLJ~�o��J}��jD��74��$,,�+�V����f=c=��u�C�`O2--�����
K��/(oUk<1 �W���+�$,��/v����k�*�m1�ҹEm�|���,��0-�$IΡ�NC�O��+�fȷxPќ�J�����w�CӦ�X5/xQ��zZ�㫃p��l�~��1cps�Od�D�O.�g��>ꌪ���в)C/�[�� F/��q����k�������|L�IEVXc�<'k��zU�^6z)�<wR��#����~���#�&��E<Ć�&N-�])�R���g4I��Z���Ia6�u�!0y��?q���:���8�L���i���*�ʥ�H�W�ϛ(vgOҝd�+��q�د��˳�kr�xp�N����3]���G�8s�-(�T#���ð���5L��0\�QEKs
j��{�������L�ג��a�{r��pOu����]�����Z��vd�����g�1N����ύ�����81����N�Ej}� vW�}���<5��p&�h80�F����{W���xj�`�v�]lnLx��_B9pX���I]|�.3��`�M뜭;J#0�-��,Z�>�����w�<s��H�3�JM+���%� "��3�Jw!u%)�:�:��Q��%h�	'��C,�S��~J7ү×U����|�Ķ���ד��9�:	�;=ɭ�830���=9��J��/E3� ٥�g|B��\\�T�c�u�!������d���?�'���4����45\�2��=5����UJ3(�T�#9��<S��t��7 �t�Mv��bgcPz&�����;@��&߰��m������K��?�M� �9�����[$��_���g�oP/��"B��+]��AN���E)0;����[rvfR��66��Z�/�d:�UMɱ3�1"���RGc2 ;$��X܀=,�u�bw�!��ό�x�F#�o�"A�h�
<,��Q��>�M<\|saq���΢��`���zB�=dn4y�9��r�s�E�n.y_j�Z%��(�-�A�m�˛����n^/$�Р��?��������������m*�m4��rLv�T��mGD>8B�C��B8����Ɏb��J��ED@3أK�����3��C

P�H"duvw�u�BX�/���� �ZΦXz�c�����oz0���M�^������T����D][yGg�٩IVKMAʚ�1��dA@��f�J�4���i�6 �ʔ&�/����kn�!� �@�(��c��.b���}���d� �J9�"�e�g������;cSSd�8��O�� a�O�8:2��0�lb+t�?�ѕ��6/	��+C�L�y��A\�w��)N�����N@�Gs'^�vW�����+�"B5XK��T��]s� �c�yp�	A��c>�S5t�� ���i��q�LsоBh?�J<�h�j�"�ڨ	��v�����'�A�����6Y��,w{'`��˼yˬ�^J@ݙ0��F��tx�\jHd��x���pwk^���`P�.�\��)���y��2�� ʿ}!� m���ƕY�/�K��5�M�fhձ|]5�r3w��톷���ЛK��Pr<���#�� ��E4;\ۺ�������rZ�K��Bm)N�f�>����})�m���0�+�������	N�h0bJMԥ�ӃTξ����,,Y�?��GD-�҉��Ei��-K�$"HFI�/׳W�qw������K�.'幹\���.��SY�K��年3>���fpa)�{IR�i��_Ԥhz��v]6C�o�NN`�L�Ź�3-�?Ȍ��j#LS��)C�ש��L��~��n[jq�T+�5��$��tC���m�/U��Q�~��4_�ʻH�PWs@6�e=��R���~\�Qv�~_Cl��41&�j#�J��D��kY�������>p�W1)����%g�H��B�{�Ӿ'�H��J�j�i=��8��J$�jT�H��b�u`����	�3fr[����M[�8�ъ7�	"���G�����н�w>�ɒ�Ѳ�}3ܑ0̿�D����"�[0��{&��ňr&P]��W�v��w�?e�"~��ro=bK��S~�}�5�#�+)�f��ܼ�uy���}�_*�l:�+@oAfW�^�G5*gֺL����vv�X�2�H��]�a�#`[&��x}�P0ȅx��W�?7�C��a-��V�獍�o�fQ�������t��+:h�[2�5��O��,N�[�n��[2���(�p�����czg���?�*r~�N1�z_-b�ƪ9${p?�e�u���g�׷�Jr(�G��OOV2A�.�F�ğb�s;d�t�ww���n�&ZǪ�2��#b=�I�����CI侀��]=/y�����%��G;>��rC�@7k�盙�'CqI*����3�x��c{����AE�K<�0��PJv�@/MS���茤�����V'!���-�%��W�LXn�M�j]�}���_�&�%ɪ�����!6=�LGZw�M!�1����ԨC�I�|!�8n����]-�SH�.+4n鯑.��a�z�Q�PwK�8�Z7��Ai���>�m�=b�*0R�A�;vrb,����%�	�j��fyk}���Ӆ�i��g�b�TeIX6��;�]B9\�~�n���隂��ӭ*��t./�����$IQ0�h�R��4�'�Y-���[�CTTd���CL~>X\rO�E�f��A��e� �pJKоR��QN���B�Є��0������Zq䟀ᑖ�Rѧ��2d�@�����s�y]6�q	�)0�9$ũ���
����������\��;r6��3�)�7l���=�=��ܨR��wu1Jw��6�<���~�ǰ�}'����p���@'Pԇ��,Ѥ!GnD�(GT��c��T�ݶ���U�
�G�r��|{�u�!�i~��b��sxox�eI���Vk)�*K�:��CBY$c>^n5���~����^��˚��x��r��&'� ���� ���`��^�=�McbM�Ag J�ٜ�z�P�������Ӵ=�O�0����#�Fe~�<�P��=����6!�V��)Uy��]����%��ЃȎ������ߡ^E���
{
��EB�NȐ�Ω+�Y�#1Q�%srC�M�^B�5��қR����R�=G��%�
Q��oM��>@��w9ei��	��,%�,uO�lfZ����z�ݬWɳD	!�W՘��kp%Y`6(C~����LK�]�>�&�9$�ic1�X���c�y��v�?�	x�0w���r&�I���M3@�y�����}XI3���ȨJY���I�s�;D:E�O���4A�:�j�,��N,��Zpcj0C���Wf4Q��\	��B��a)�����n���9�����g6���J0���O�k��i�R	�;t�~�����u�οM�,�����5Q�]�nW���N��-���<�t�K�H<�r��>^C=	�M��g\�<N��ԯ�繾L'PH��REt��o�<�6v��8�O�:�"���`%����~פ����Δ�Q<Kx{N�t]�(��ww>��d��B���*�@�����x���Ԋ)u�>���{�i��J���K��̞�mͼ��-HŻԻ�)�9d�7j,l[s፿+��޾UB޴����+F�ֈ�T�l�kE R�Ю��;�m�VJ]H �¡M��Z��މD��c]�Io�6������U�htٔ�h����6q�e�����P�> RNV�	�唎�pf�[6U�5����,.��y���aP�$l�����L��	�Y���*�?2]��G�=̘��#�?qe�z�7�)b+� �C��Ƭ	�8F�z��Y{"�g2�w�� S��\k~��{7�M1��d�fw*�{8F¸[�{Vl�'A�q����h��}T�c_4M���!+7T5E�tE����<
�ۗ����+yx�����wW{d@2Wzo<J���]1l7��ŞBT�R���a\��M�M�i�('��}^}���e�s0�(�w���V��,�
��S��V�g��<���*$��m�go�K�`��jk�Hy��ϸ�Q�2S��sB�MSK���ߜȄ���I�X�~��t���0�
n�S�˕��?�v�r����+�1&y;��(j<A��T�@���ڟ2��.�D�r������0�]nr�cPs�����Q���pL�ǵ28����V�z*��_�O� ��W�"Gp��P��;��=N;9$q�o��ǓH��Ρ��w[ٗ������gYuBH�b�K�Є�����6K`�u���Q�k��}����������.�i�<h$�%�0��ˊ� �Z:9R.��"�:��#�����-:��o @�e�i�e1(�#��'���&�D����wM+���?ɊU��I{��C-�	�ǄO�c]�v!����K�+���#�Dr�z�`��i6�M��|,/��H�O���ߡ*=�$.Z���!h*�~1���CEcG\G��@^�2ʵhC�o�z�o�������2��F�w�m�Ŗ�PMn�)ʈ="��&�T}�JC~�K��B?�*�c����~Џ���b��QKiĖ�']b�t�1Y%��+�?��O��ʔ6���$z�>tJ�Z����߹?�RL���2�c�����:���i�U�b{��sg	�3`oq ?k���gS%�op��x����׼��e�x�^�Ӵ*GK�ғ˵�Rw���*ߠ�3�E!�`�B�P���{R���ȝlذ����n���On�v��!���a'���	���`�g��iGG�,rؓ6�] ��v:*��P��xv/�}j��K�}��^%������C����r�����h�bNv.>�H�8ѧ�ȓv�vY���#ouTO�CV����\ɳ|�M���(*ɢ�"v���1<����ŏ�CW�@ w�.T:����ns(�^��ڋ>>�n!UˤK�=b�(��BR�Tqh��(�{���Q8
7$��<Н�^�o��7�G��h������H%*�iz�����vΨ�Ͽy�ΊVlPU8p9*�TS
x��5��-����5�SC�2��t����W���'~�IP�����ar;%�x4���'H	��&+6Y�'e���h�o�$��������;��m���&w���B��O�W8��LB��]���<��k����<ᒡ�-*�3D���3�g��O<��d��,MO�s��>+�=��=�C���a6ę�v���Q�rczk�_o�Eo�`onix�Kg���x�G�P�9�H�kRe�y���\�%���F�k� &i��G_�vWȅ�|d'aW�y�l��n��覮�s������Y��,:���'׋-W+TV�6�%�9���`=;}���dá�S����>�� �d���`Yk����E�d�OH�=��Mj:B�TA&p���I4�+'کU�6H�#�`	����Ҩ��¦��f E��'���FcoC.��� .ɑI	�!��ϛ�~�8i��ޗ0��M��Y^���%�.l��ڦ�\�>�C�Ol\P[�/���A�	!Ŧ�,�ORe�HT񨈭�]�U���v)�˂��Go��O�q��u[S=��ѱ�6�\_���}67l���={�,zu*�ǐ�:����)"5β�*:O��ϱ�Bh[��&����;�\	p�3e�d&�6�C`��[[!�8j��',b�1�n��*��(����뾃I��Z�b@L�O�Z���h�^���I�;����ry�2��1�5�Q��x7���q�W��H+J��-�U;����~VP	�HB���;L�������U.{"��`;vP��hN�@,��̣��ٳ5S���[�&v��n�Z�1�kŤ�td{n]�:�H%S����1%'����J佦z�Mi#5N��԰�y��;�DeT�S����}���#�|2�z^�O��y_3�u"��r��{N���z7{��C�·{5�Q}����'XY���'��
Aߒ�/�XV�k�W�������E7�7���4�:���VZC�"-�Ϙ��4�q�}�ƛ�E�7�Y
.�	�$G���5�H �R�pi9G$TNJ;g סl 0���(R��1�d���.f*Ů%�����t�|		X�@����9	�<��E�]��o����Z�z��,z�!�e�a�J�]��KC�-�T���[�L.�!����<^��y�9T36��K�f��>6�9GFE��ߥ����}���o�W5{IS�\ )����r�×j����Rƍ��D�LQ�u$(��0�G�\4Gy�m�� �u���Y��F��� e��8�8
�m��DeV�[U�����Ś�����y���J��ｐkCe3�Fbj����NRDq,-�@~h�D"NaOu��/��ݤ��G>s&_[���9���-�G|fF1�F��j�g�=��FGG8,<�S����g���M�$���Ǌ�Gm;�(���f��������Zs_��$���7��F a&q�ǸC�b��J��!s�X�sf#���\ ~�d5Y�%Ck�3,1�	���ţG�|P�� '�!�9PQ[���~{TV{��@1�m�;z�>y$��$���?R�
��>�D���W���2W��o��vJ�V��sm�
 �V�ץ�{�D��#s�.�Ⱥ~".�=�5�],��.���f���w>�<����^�������{l[Na��醗g��
�� .`�꺩�=�e���xΩ����9ʼDV�
�4�r��Ot��I\n�Ჲ�.߿�A]Qj򔒋�
�����a���Sí�T�¬�}�K��%)⥓Q:Ef�����Q=6�C�ω�߰η��͵���	+/z�
��7P�X	��Pnm�E]���F)��=�-󰵟4�������p�_�a�-p �敺6|��A�doF��|�]��Y������1*s�\a�!�rs0P3x��E��beYs~f/^�0b_D��P'�@�Hv�!���l\�*�\K!^2�@�����B��A|x��1o�S�N�^䇶',������B3��M�0������J�чCM}­��v���̭|ѕ���$w>����$��5
z I:BT�4qpWp��]�q�P#4��T�b�45�3�e|SFuk[��,�s+W��a!y�L7��ה�лň���:��J�k�:yi2>��Q ���L�Cp���������o�P������KÖ*�����q�O�H�e�6?k��;YšH?o�f䌣O�Q�Dm��")��T���AO�!�$�p�7�öV�l:�k~��'"�@2�-���Nv�R�f�����!��~h�y�/�X���������n�-�ǲ�[��G"����ʎ�j�����5�Fq�}Z��kj�5�9h���J��dK�i��橯��ꭄ�C�e�
��i�)|va<:�qóB���t�F�OZ�BEe(q(bhs1F�*�h�(тK��o9w����:���>�?Lr��k�$�v|	��j��:���2��S���"`����p7Il�. $I��E��O���G��k�_(ϕP��M�WxK�-� /	�@���JR@.SMs����凷i���\&��|�)p-�-��M�}5�أE�m|aYU�ˊ��BWx�E�+=� H��&K���ҡ��r6l��QD-��W�FQl�)#v�>�2��o�������&�!�@��Y�t�K�Iʿg����3�p��v׎6A���u�܍�kf�,��I��i����쮮��?�	��+R%E�sԸa .���&���4�g�<���h�C�����9�u�� T�"��Pqî.>ܫ��i�s�~�t'��?#q���pOF�ۢ�O�����{;? �Mnq)-��a�h.#�����\
^k}@�4&��$N�[��D#"�d�ZF8�¨Q>b-�S�[ ������O�9�͜6���'i��<W�L�g5N{ҾMg��N"Ɵ������!�(���UFc΋�&J�3oVē8#|A����F!-{��v(���m�<�`!�q9�cf�@���!}���j w�}�1�ui���b�wÄ�t��!�� >As�'7a,�ܤ���Ԇ���5[��g�zV�WS�ψ  ��D�@������ �Ѕ�h=1��Z�#K)�XوZ0�����
Հ.0�3�,�s��$�KnH�ܗ۸�~+�{�H�:_�ݳ�$��>:����#��K�^�K!���^;�~��N��M���]�\�ۊ��pʹ�A 
�] =O��blp@Yqګ/�'���R.��2;�b�xr�@ʊ�Fᶠ���Ȗ��W#��B �g�H�)|��T�a?�Gl z���1�k<"T���j���i����!���P#�3>9�HBY(#m����?ib<k���4j혥Wd&a�`��m�Pٕ3�|�J�7����]q�ә�D �Y�#-X]�������ūWZ�#� 1��	B�q�sr	�`\K�/�Z�"G�t%7�)�ICUK:�� r��el1�&�d[��&�a8BR<��D��<ӂ�ʣ�ގ��w��iˊ����ꝗ���D�J�O�MDS�"�aզ������IaƓ� $d*y��P��<��3v���*1�/͸Ñ#��W�:�����F�DD�TM�ˀn88	�iv�����0��e ���>`�Fk�V�X��q�\ �X7rI|O@v�r��ث�R��_�#�m@��jM��G)���'��x#����7�ˁ؍wQH�E�[(_����x&�0��SQ��+M�W
N�%?�����È�؂`Z]^����3�_��55�iAdj��f�V�1�VKkjF���=�W��>�o6nsiutC��+	SF��+0*����VҖH�FY6��l�-?/T{�ה{dGH�_��)ވ���_}��ݝ$D71�}
sfµ��JFm��� �&U�G�^6L�bdr���T%zg�}�[Er����e���S��-��KW�]Ayp8���:�*����J[��n�*�����/�$�`>!�$�i�
����e�Xj�	cɜN(A�;���(]$뻝��:�lo�EMC���Q(��ܗ5dR?�b��o	��Aj��$�I�r��+�}�P�V^�~Oۺn�X�ՔL�����)xS����t�����=�/}����j��V&�0�ԛ�>v�?�0ଂ�U�H#CƛD '%�U/dm�����EQSWG&l|J:���t}U���V��H�f��a���2R�@q����'G� U� ��&c͏fwЬ4.q����z]�c>IUqё��6��a1����$��ầ��2U7Z����;�TM~�!�p��Q� sy�@-=�U�Lj���K��gRoF��Ӝ�sC�r`�4��o��To�3�r��>h����6���E��_�_�B��y��x{:T�A�<s	���l1�7�nf� ���^	т-d��0tkoq���a��.� ����	��~�ڝ[0K���?e���:
Ś:E����\)��x��D����X�$�e	|�P�n�rU&a�@�����dy�e�{%�2���jj���ɭX�Y��z���_��#}mn�+�YYJ�����a����'h�р�&�+���-����i{2�1S4ƹ�C�'��[W�j��5=v�ͼ�����1�RVo:���-���7�Aߕ\�~�{�R�k�q�������s~׾�ߊ;���/�N�Qj���2��)�/i+�H9JM�
���
(��}�t�ګ��'�\��_H<��S����_�'�h���0��/ˢ,yo��uV3KN���-��T�=������@�K�НW��P�_�Uد�
��,۔�� T$i�.���)壃i���1��zōU�b��@�<����Yɦv��Xdp�2�q�̵ �����F"^e
���LϬc�m��,��m5:�i`Tϻ���($QBye!��
�ɘZ�xq�l�$.W��'�U�Ps#N��X�E�U7�5��L$�jQ���)V�`����&yn!G��{��h��q��?�h�M� �?�Ȉ�:y�������X�u���ǡV��@}�S��E�@�	��hK�Oim�[��סok�U��7�q�7e�<�5P|uja�Լc;��)�����V#�aZ���iu������%��������>-��L* �:n9��l���μHf�IV�'�A�-l���{�i�ڠ���g2o%�@L�<ql� ��kB?^nl	Y�a��r�y��à!�\�Y45�;:VM���g�[sgC@׎�K���uc��ɡ����ٗ��gs{7G>�;̅K����E�~#q�Bi[�s{́�X(g�0�ڗ�>���5B4ͽܰ����	1s���k��x�#�PM�1Be�Y�Rp~�71��!�T��*Kϫ�F�/��B�Hwt��,�GC�0J��Yr�*0o������E���WD+���Vb:����nqsųa:7�U�Q D�%ۮ|ڭ`�r[iӱ{��� o��n� tFU)ЊDqq���/��_: >�:�N��5o�S�{�f��c�'j���S��+�4F���_��\��G�`٪唓>T�Y�Nk��3-�R�����Sr��,���$A�=�3<�"^F,���@*���y��#�*bT�?%ܖ�u�
�;%��(��p�WTY��MP��Nc�ʱ�rj�N4lyu���5��lOو	��V��&���Bݡ�#\�[��3���8#)�'/g�:��A8���8���z5�F�,] s ]�#>��6T��kOI�d�-N��8=$�����%�,�,���?$�V���>l�!�S�bj����^��v3é�	|n���y��ZT	�J��g�2̆aE.��6�5��W�b���5��8�Ms��u:"�΀{�"�Wx��J�m���Yi��f��f���O]�"�v[���ne*�!�?ܴ�P0rf!I���kS�ԝc�'j��L�����w	�f<_17��U��O�%�W��6�
��4ctH���q�ne��`H ��9<䇖���E��1�L�mz��b۝x5�`�v ?�URd8<CE��@N6Uz{������5y�0��oĖ�Va����P>y�Y�no�c-�#�$Fۆ����rK�|?S����zM�rٺ�M������N�����>mj��.�����2ߺ�a������66�g\�آ��0�FT�I�!�l��Bz����5y�Eom�Ķ�W���e���7~�wn�t��,v�-��f�-�4�)�X���u�B.�����ǟ�b���}&�PX�/.vx+�H�P")p!��M�Of�:.F� ��2�4��ƹ�9۔\��,�Ueu�We��z�D �4�d�)9vV_e�'���ReD
��v7�y�M��	T���������z(�դ���g�}�P��>� �lۀPEҔ04����߼����/��wo�k|��Q�e�ĵ⮜�����;,�{��h�d������$��8	��pr��__�w��֠��eLM���%M��q�C�4΄�I��9�<���ӻ��w���1Pw������&a��L�vP�&>H*������!2i���-�j�t+|�� �f��+������-/y|ea�+�$��E1^K������M�����2�{d��T�n�t

��❌�2�Ճʉ�	�7�T�AN���)��`r�~4��OB<b��f��"�0�n�����qT����+¬*�y\(^��=9W���&�u�]V<຀R{���u�>�����{`-	&��2�@���d�N�ְ�i�뼯�0Y����W&�2�y�"T�I'O炥[�O����~#��&�[������<���t]g���u���O���F����T��ީNz���VQ��9��n�Xnk�n�����~tF=��~Z�A��:�7lU�q�o�xV��6���#t�+q�3�D����~�!K����J��K��~\�ǧ2��A��ݳ��5�,������\�x�Q�&�Ϡb�CƓ��0'3}���#��^Jo��Vs��5|��z����v�:3��N���,��L�S�T��L�hQhѯڐ��Y�����������t>�
\�L"[\���+Rb}�
��$_l`:��¢y�D�¬ ��*���n��O���y�(uY�m�j`�� �s`�?�p	4	OJ_d/�\U$<�
*9���P%�]�+�����(7�0[��K��9��M��~�(>7� N��G�Zb-Z����Sd�F���C�'�K�MF����2��,i?�{�4$�I��S	�h��Up�h��y0ߩ2��Ď�
��MJ�D����]R�ܱ�L�j�nYn�o#�%��hj��Ȼv����=�EU�T#^8�r�Pp�f]���=8�='��S����FY����n �ˤ��E9��Z�?5cοM*��j��pn��"L��೤����[� #{�	����������RHPc�ߘ+�Oy����IS��R^�/���]�2���l����B�֬�-gYI,ꨡq��X���*}<*���i9� 7a��|5��������3���.������\e&����L����|��LIBy?��"R�.�Q��w�E��D�q��L���E@�鰌v��g�L����(��M����L�p���Txm>�8Y�����;�D�g���+����V��F!�RWr�UzRU��P[��iC�;�)����� ͐�j�邻���tAq���L��Wl�.E&�_A����;��,�'ϐ�a�E��[G�К�1�����
�T,�����VB,<fX�D"�@W�����a'HﱍmW�����?�ڶ�C��e�z,�[��(��-�#'��4p�W�ȴ,%3��':8.Fv�Qc ���d�$�Jrb�_����e�S�|�dVf�w�F�!�)�j�	7>�v�=cE�ԔK؞&�^"I�힝qf����m�TH��O��5#4��۬�.eԑy�|��&�Z��Z���B��\x!m3FL1���r&5��SE&���&]��-K�J����O.��)y�c�P�}uK�w")�����v��?�>��}�(�˼�+6�eS~��#�ꯣ��i���2c,�� 5���̇2���êg~�b���M�Ҁ�h����Ʞ��"6��EH.%`Re�%aK�Ho#i����l�j�j��rlh�~5�nm�ޓ�N�U�
/T�$�p�er���5K&��F�;��yhp�]���<_z�X��{���"�dQu8u�}�x�nգ����Q�X�j�Y�i�C�����f�UE$�'FR��X
hD&{Q-�/$"̽k�E�FEH��:��Y'g}Me��������ve��EMoa�I�o�̩�촜�>s�!�n�Q�z�o�:�+��gcD�d�}�)����p��Ŕt95�`�mY]qu?d<�lȸ��C�9*,�0jyBzb���o�E&��������臀CI��k��CcrV��Cs��C9m�9������o��'\=�2j�'��M�0v+u����D���U8����v+T��Dp��N ����=�>�6�3��*FϬ����J�����<�o�.���+6۾H��">�b��Z͞&����x�D��W�J����8��[��]2L��V,�}��0��xT��?����ĝƭ���<�J���T��5��M���[p)OuԆC��M3�(#�C�o�s�p��j�ډ����XI��B$Y���4xi���W����@�b		/7��]�}�2c�~�9�o��7�eǝ>R�@���Vi��<����+��S_R�(S��<��B��v>H�*���Xa2�D�^>����&R=�b�WB��J�:�� �c�I5��5�2����nQA�AG�����eh�z�`ԁ�٭�C��|X�M-�:��4�b�o���܃-�f��տ������%�l�s,�c�T�I�9J`�.G<z��*�g��ieB`�I������lO��E�1��r��ﶱ�K$o���`�=�\ٹC��Ƭf�
.k�\-��u�BhJq��Ea�Ɏ��х��M�ޔ2�|r�i!$=�r.�rnz��0��_�>��N���hI�s�*�4|WY�L������p�Q.�B�59�ޥ!%�Z�#mŉA�gb�8��䎊��C7�ׂ���^h�����5��Vm��L+�����[[r�	��4���#���[��J��Bb��5;��h���.���c�M.᭰�,SL�R��B�ꭆ[�K�r��p-h�l}�.��+��^�=9���`hb��R�k��%��,�yfV>bV]��NH���2��,FG`�M)�C�"&7�
�v�h��~p���g��3:f���g�RA��������Bw{E|��K�,jU���kj먙ɇ\!7ѵ�ܾ�,�'���,0}�|��B���<x��� 3!�j���pg/G���	D�ƻ�tڱ0�a�R/\>��ק�Gz����݃��F�s-cH_V��Z>m)Bi��߈\3'ȷBZC�ze���?!T���)dZ�1��<�otFB�w�0� ��0�2�"Kƛ��o���N>cL��Y��-�[G������<������Ry��-^l1��c?�F-w�@�{[$#Ή�)7P�O_]�Ls
�+X2��E�v��۳�?#���<�ݖ�G�'%� �'��kz$��)�*6�N��Fl Y�������J ��x�[����}�%���$��8�r�E�w�^P2sZ�DM�u�v3��Ʉ(��ۃ6��{�E�X�=c � ��@����&%��]?*^�XI��[��^k\;�O�i	���B��z�(��a����>�ĩ�լ�$��=@�O�A��CNЉ��/��|k���,�t�0��#I���rĻ�E �o��n彜yi!;ᗼ}��׮l�>h��W#G�Fb>Yb��CVB�$���pY��F6$[�k�wx�8a�p�`�y����
��2�ʣ����x"��ׯ���PP�Y��/���{B��>>��	:�M.~L$'���p#S�C�R�Ԅ���-CXp��-CyIϽ�����H�7@W5v2�=xm9�	ɢ�]}�?�?�C�(@6�Y�R�7��Jb�rA�q�)=նꉁ�w�Ar;�l()i��DTe	�&]�Z�𬊚O16X�� py��AWw�_l��҉r��p�*[���ϗBIJw���G!�׬(�Gx?�P�zŷC�;sD�M��a �Wo!��yc�;�a��=p�'�k����il_u��q��L�ۃ)��I���R��N�����b|c�M5T�����a�	�,��U*����ǥ��?���gCz���,����n2���j��H��l�����|K�'�X��z��e��mj�=|��r��A��YXnd�M��G�n=�1:�S|��T�蠺��Ogp�K�g��ƥnHU��v
��rѲ�b8�^n�>^�ɋ���+�u�x�z�:v2I�O<r?�Pт#����4��r����Y,��P��0� �Z~�"f3}ܣ4���$	��7����c����,ҟd�;�a��ԩ�7(���[��TX2�Ӊ����!�B�EWV������D(�l�|)
;��6�����u��X�\ņ��蚼��"IP��B��+ZdǑᘐ�d��3�� ���C�4E�\�I�m��4#
�^VI�&�c��c�c�K��ǲ��=�m���q��$s`�@h�y �>+�u	Y(Wn��'�C�;9��ә�����'��vĀ2��G��p����]J|��+�XO�{�t��r��.��z?ؤ�kr�V���N85X�d��9X��$���6�#����®����8�Xf�Y��±�0~.ӹE|��� ����2��T���SwZ\��O*�V�\��x���1�iL"��&ePQ�ɳ�y���Q,��[#�N|v@n\����%�*?��1˹�-^�uL�8Rn��L��Ā��-q��}�
K���\���Z���.�4|��j��g�6f�U�H���A(��=�&���D��ҫ�c�8����Gˉ�=���~��gm��I�������ÈU﯌����l�cb9�O6^K���FH�Oʯۮʢ �h��S�ߐ��\�hkm#�i� �Ol�,=���T����m��j�Nu4��Z���|?��X��_��<�n�=�tWqk�(���O�0��������Ox���@��|�J2�+��ڹ��x��R���B��H��x�9-�j�"�����!7�ob��kᅱ��:5��
kuZ?�Pc��)��o������M`�:��F��q�,���R�'�&~��Cv�>uR6�[��p��D7����W�s����)�G�.k��_���dRc��\�yA���.+X!���Cb�����X:�k�C�B�NBWqf��ڴ(P�JӅ:q� $N5��a5�o#t<0Ij�v�"4#`�ù��w��O��rH�aN�ry�ux��������$�$��������w_g�(�7f�N��lz��vs��$c?�u��D�̕=�5�H|���B�b_A+,�� Q"&���2ҟU�A����]�yO6��r ��of�T�AĂ�u�F�Lao7泹��e]]^=�����4`�8�Ш0���������R�=��$�yPʬ�t&\���iA4$铞��s�thh�v�cD�l�B��z�_��!�I�Z��<�+�Bi���tl" ����4�l/OT�̘���0���X�?$Zȿ�B��u󟝼&��|Φ�\v/@�k�X*��[X�!�����n-��M�E,���; l�w���l!�'�p��P���Ev+�c*�I'dԽ�g34�@�E_��QSt0��7;�Ō#%�$�O�����p2�UY��9|�YIL�]���˼��{\��D �W�ֶ޽���.�:�s%�+���F)хz^K�=}!j��B�m���>�G�1`i���ZT'���԰]��׏8_����v����n���{B���awf�L�Gg����)7�~qR+�>��Z�|7W��ƥZ�V�橳 � � N�kV���:^��ew̭��)�>h��&h�����%���Ft�d�8Xm����ܐ���@p�8k�}�_]�K�0���i��e�gj�<��@�����wK��%{�Q#�0>�V�t1fN�����xK 4DT�uQ{�+����f3>LHQ�������Ow�ǔ��X�X����\��]��=J�h>�A�pޚsbkU4�C��<A�h�J����+s�D�/����:�(��a$-17/��� �G�jP�k�B�ά!�L6'|�f�s�T�'�^�oژ7�͕�j$!{P�xm���"�)$�񖣲˃H3
��GDˁo�:� �����gZ���6��O'���lѣ2\SC��n�V^M�M���O�Y�VK ���K����oi[�?]���o"�~ف�6A@N�.�,}�3���8T��1�G��I�B�/�)/IV��b��փ�����e��٢~s�v"�T�}%��"tX`���5M�^Z��Rº��X��8��`��l����Ka����C��Z�hL"�Z5�Th���N��K���-���3F�_����[��d�[t莛�$��G��eԱdu7	�[xPLTj��� �ʜU�]����S�ƽ�\ȗ6��&i43�3��~Lsh��v�y4-e��o�V<j.�ٛ�1����.E^�\^.K�U=���L!%1�G��#<8/zR���H�����aa�)��(��jih�L��Dd{����\U�	-#g�v~r"\��
|sj�:��x���f�FL�,P��|���+;��+��v��{�]�x��ʐNlHq��г���^ST7�5�[�LI��t퉥ud�>�ٙ$m�LB'3�N�o�zWM}��L�K	�Y~%���[6�]����F�'��e��<�]����E�Ij�qg�[T�#Xa��8���j�Cn�J�#į ����e�Dr�4�ًK�㹠@h��Y�����`�-�����'���	θ����U�t�hi-��pp��v�*K�e������h>|��H�v?� ْs������ k���Ss����,���Tg��9	����!���/���!i
�;x�]J����)��6��KR���m�p�˝����7�s��}DB�m�k^�}���^�ʩ�d��P%ǋ�$��p�/�g}̧�*�a���;ܸ��S�z�9�����Xs����j�@ĖwZ1���疤�7���G�v1�tp{`d�IJ8;��R�����MM�[Wcg����4dW�I"�G&� ��ր�i��\�������Re"��������ΰ�9�L�̄��5�D�N"^���z������q�����<c�=��x3A�*��r支MF���O��l�g�;��ʓrI�n+%ծ����X���B��>sm7���33� �� �li�t�����M�U� �c���7�����_��4����ƫ�����孟u�AOa3������Y�y~*�
��|A���`R�S2P�J�W���4Q��Cm�}�No%F���+�p�1R%��_�	�K��5��u?��yC+�������k�)�ta�Iʕ���ͽF#�N�]F��s9�A<m���lM���	��ru߀�������Gxt�)�Ȱ�*ǰJN7py�3&w4A�Ce�&p�/����zC�i=�K�-轨v�+��]|���1�37N�y��T���]�2=����6M���l�8��	������.-q�5ܶ��J��[�Ǌ�ow���o[���W&���U���W�ן3�� �]���Yo�9@n�K�"W@��Q��;W���)��� �5�!�]�V��L�J!�)d��r��2�y%\�E�_���]�C�=�s��x���k"4z�>A���-�@qV:��0HoY��;�E������L1����߀T'�"I���XN)X'\��;�$�-������8�?��n�	>d6G�3�8�aWe��E�~1��J���I6�E��/7a�:���+�k��+/���ɦ� ��%���#U����4�	wQ3�8� �)�[	VbZZ+�ȭ�S}b�[b�+.����Mc(�["]LvFɵ��}O�\�� ��o��4�ߑ]�O=�����]��q�ôfX`ڨ����!�.]���k���| �(�e�X�R�8�Ro��\6�6�
}�-�&{�C�L��/�W���ש�.��A3o�>�EVXx���-+P��F<�O8S:�;פ��vbq�e�چ}�Wέ2Sh�%𑛋�QD.���:T�@z��6�1�R��NR�Z�J��s4:�5_4	�zL��zr,Ub_{�i�,*�L�0����X㧶��O�n��ӵ�Հ���v���"�[*W0�..�I�:$��+9VL��Kx�&�*?��[�SÇ~���!��+�o6��x�`��<G�������{�*}���A^-��!�Y���*L���5zx�*irf?�`���v�`�
���Zz�T-��[Mx��Q��C/R?
C�TB<�P)⪺R.<�Ϋ�G�kE+B�Yp�Q���,*Q@�{ qj/�,N�V�{|���D)2f-i�B�IK5NI��<c���B~�< .�(X/%|ί�&t{��.:]�a'�H8�-�[!�<��3[R,A7[�@$B�䥘RK��?��f0s������|6�.��'v�w�1Ұ�S��U�xo�8Ǩ�K��"̟^�z���[�#��kW8��������;z��e3�D��T�b�r� gR-�]V���B�?�����C��t���į��U���M6Ń�`����W/���~hʙ���V��oEЗ����2�ɽXA$����7d�xu:%ƌ�Be\�ЍB��� %��բ#�A�M��c��g���.,gR�T0|�&��t&�w��mU��B%����q�Sɸ4u���^�~�D��۵__,���q��X��w�V}��f&����Ġ(L E����ʟNma}�HA�}�J�������_V�r�t���ؙ^����$���0����{�ì�l{�F�}�^|a������C�]��8�C��&�������!�7�`�p9w�	m���fk�v$�MA�uΪW�������֍�s�����2?�1o �!�̪��5'vŁ��V��m��ȼ�->���P5�L����TE-�1J��چL��x�9�X���w��c���~�0��p�!j�"�����چ#�D�F�~N�Z�8��#
���Ol�щ
���`��(}4�Z>�/0wl�8���� ���Òٛ�<
U�Uc�7�4���=c����rb+�Jn�-Ѻ���\�a9U7�����>1jK:�~�[K�;�ʤ�}+cĊ�DTX���x����' '&�)/���< J%�������<�|�9_PiJ �� {�{�q��@M �5q�\�Xۂ���$~⥾k�~�$�tD*�ke�!��H]?e�9���G,�OP�:��zߎ`�h}l><���d"��	U��`6&��ܠlC�r�B����VKs�<1%�gt꽗��)��[%� �]\v�{�;��?~5�B-������<��3Wdn�)��\w�ؔ+b&��D�hݙ��_"�����'»iz�������[%��=�ͯ��Gx �����'7�G
�o<�Z����ҏF��pG���>�������Wri&�66������iw�6*�'�P'k�5�z�i�2>_���n��Z;Z�^�,]��?Q�2��!?�m�2�Ş�G�'uL�^NOf��b�KP�����̲�C��0����C�<[��`'��� �KF���`cG:�#Ӆ���s��;�s0�o�	 s�>a��u��^c($��3�ۗ_���9���9U�1BE�����C\m����6DpY�\�{e�Z�/ҡ��
Ub��%�#"��o߬�.x���
�F�=��^��l$��NJ�PT#h�-���s%%u���X��b��s�^��B@�t�"*����O�ţ��&��_����9����J�U
��mvg��Kk���"��e�r�j�G�b=��2���b[02o�rpV�=\"�Y�|�	 R3��#���K|���+�g9��tM�E��+����-�{���J��I��YRxyfpB��6����srm�ʟ��Ra�A#|�lq�8�F���)��m���w�ߨ�����_<r6C�J�Cc5ɪ4`pg5�8	�&���Ew�^ �����ݝ��K;����mj���\��tP
 -$���,����Xy�ڷ\������w(�q��L/Ӭ@ŗR�� j5ƹ�l<Xj�X�'�-��<KG��?�L���8����C�)1�����K���mt.��~�M�@A_�EC�?-�����H/�J~��5�5t/Ms�.pwb?�.Y�.���֯A���D��i����\("�4���A�e�U��DP4a��hEx�Xi���_}x�6>k�`4i�6s���w��8����F��6��:����ֽS�
zŹQ���J��Kڹ��n��2:���4�' �~:T~y>3�<(��}�U�J.�B�M��%���u��"J�����╍�����B�Zs���x1�ƷGo/�T��f� ��a����(vT���T7?�6�i���y˰A��8-�f��d*��*5u�����wHϚ!A��$�g�Å4�F���m��.�ڶ�ثlo�;A�o)B+������ͺ���v�:� ����2�a��ȷru�(1xԩ�9�>�#6I��;+�����8*��("�ܚu�MbZ���V[�Z$�V�)¢|�l����;�C�]�(�Gy�J�q戡�P�}���j���\D=u8Td�m�_ŝgb?!�H�&7���γƷ.+Q0��&32�s~T�6o��� �j�xΤS[���<�z�Yn��Q�N�|�i�P	�/zﺜ�R����V^��.Z~��5��~��<��B��e��^\d1U����5��i�	٫��=u
�:c�CԖ��x2��sa��(�s���x�c��1C�0�Ou�=G)o?�j0�+��1�[�K��Xk̑!��
��H��q)I���@9��=lʉ ����?>Z�=,��e��" GX����@��0s����Hk�O���ū�	�=���)~Ԛe� �D5��_W��^�ud[S|X��c��G�!���Bl�,�2�A�Ҍ�E�A�Q�>-� �>q���ϯg<����	�L��ǀ:�_�ދZHH|�tMӤN��%�V���_.���O�ۚA�V[Hm��p���Ct0{1x�"/�+�V�6]<%�����{��[U1X�D�$L���v�b�N�x|�������^�`#H����Ok �Ȥ�0�Rħ�v�
�eߢ=�U��C �3Q��[#����LII�R��tBp���>�,<3�t�v��6Ӹ;���~�P��G,_1~��H��+�ɛG���J�d��-���V�W��X�1y�������^b-�����DIN�x(T����+��B��`�X���'�$=[��b�v�P��N�M����wE�缁P9-��>��㞙���7-=����(3�<��ù,o�<\�:"��c��ۨw�!���k�?�<�ug'����4�(�><�PwE憣�b�?ޝLV�դ����zF��t�!��,�4���.e3�<�P�j����1�.c���Ԇ�$��.m��ҹ�PVf��jū�a��Cf` .���E�'�E�,�����>����?r�}��/�"�3K�v6Ƹ��yp�����p?w�������%�=��
��݆�7��E <آJGX1��bvw��[�HG�f���_��j�q��v���V��$%.\z����8��3�W`k!�wOm��Ӏ�7���6(��C�K�Fd�5$O�nI	{�_i�	1� e����+�j57��O�|�鱪۔�,Y
�K��t)���K9r�*_k�2 �Vs������E�[F��Z���!�P�� ���O2��7�wU,,�E_G���¹�&�w8���[0�K�A��-��3/yyc,Ș�]��K�P�x�M%�'�zx~ds�l�j�G;��7�aɕb�wqC�po������

�M��P&1������K��ɋ�ҹg��I#]Ug�Fwk�Qd��hIɢ��A�q�v"��p�Q��D*͕5G<���"|j<��d/\xw���-�*��p�M�o~y0�ު[O�������u�$��p�q4V�qg e!Js!������ d����fwF�z�*�S=�KM�`Ϲ�ը����3�S�oI�������m���Sf�ԻՊ��C#��)Iq(i���
�Vy�*����fV��ܟbݩ�.��Z��-���dO�0D��FܢD�?;��J���%L+/
�Ţ�`����S����լ͔g� |�>S~L`Ѽ��/9�1��K�Q�?�+?�V�m]qWط&`��k_��᭰�@�t��.&�����D����}2�!{�H���O�~��*����Uw^�X�����Y֙�@<���&�s}dEH���:�^:�c��,��%������<�QVykN��\)F��>�(���~�zZ�iz>�0��u=B�͚�~���p��$J�1��Y7��U�;�@Q���㼚�u�;\	�H�%Z���U���CW�&`LQ|M�a61&2��?�1���?,�:�
���>)�kP�(a�@?8b�B����uQ���X�\jz����׭#����]Q��s7x;�#�Ě~����a�B���+S�j��I�_��}�k�jdXbo��~�c�,�:V�Y�0���K����C�i?��*T�m�DI��I:諲*��Y��ᮆ�>�Nn�/R2Vr�/We/mj^_H�ke4C�W��G�T:r`V�v�Tu��:W+m��K��E��D�!oE*�ʘ�_~���]TJzԶ�� ;�J�]�v	R��z�0�T�m���Ծ7O���M;u!��8�	��Ġ~��P;�H��e��4���))����#Ц�JG��Id�,��w��!#]�-�Nx��cYR�%>�&�Y|�8f5����p�$�f@=<������"-=�!c�a6q���GM0��C��2��HA��P�Q��9�\�b+���;L[,�5WI~��H%1��lͿp8�V-�Pֵڷl��>[ ��T�,�=FG��#��x�Fe��:�֕o�k��;$�<�5x��z1���)*�V�Vr�:Sbt����"V�|5�������a�������� 4�]2t⟿ Ym6��3m��9%�7���+�Z�Az�x�.�$t���c�
��d�+q�z���f��*��*��i/v���i���TL���x2�2�2qr�o�
H�λ>�����u�1ٔ�'�V?��7�j��$`�[+�)���vS*Ċ{Q��E�?��aZb\����e�0� � O�-����u�H��ý���M���bS�>�8 ͥ�r<���Vhg�-�OدV!QϢ��6�=�u�S>R$�2�$��2;�:�۬7`kn��
����U2(�N�M�d��@�]2Ԁ�Sr��<�3q
-'���d��82,0�LW����Bg<P~a���DU���}6]� 1�L�
T_}�G��E���*,#�%����Ί��n;!�$���e�eM[�Q�)��n�p,/��s�55��a�T�db��=�㐈n��4Ό�J�쮰 J- �������G�p-s��~6��l*��P[����Kc/e���⎃l��Z��/Z1(O�_��b*��Z?�Ѳ�8��,�^�_X��jj�ls�͊ӹ<�&�ڂ�Y�@���E7OS��{�	��Y�AŮk�����G{1Ă��p��j2ߞ��s���bM�_t�T'd�������6A�/��iN�7��k�m@�2��J�(L�$�-�+��%t
HjV�C��&K� �I�%ޮ��Y�LÖ�L%@��z��e{ϸ�ݤ��J/���-�]WI�q�L:	�db��՗�q��o{�e�W���-ͯ���E�wU��[�PH{<ʄ[o울5v���*���P�E"�5o�q����/-z��ľ��$�{�I��w}h)�De���Y�����JN:�Us��Bo�����+�Q�&����s�X��VB񢹅3Y8�E��]�>�W��ƫ��={���P�Gn��KM������������I�w�Ρ�v�@�m"i�;�LJ��ī�ȳ��k�a`f�c��%�����\�_�(D��ft"7C���w�O�c���oְ���Y9��d&�D�r/<���P@h��sa\sd������]�W��n�4�n�����Ma���"[
&H�{`C�:s���7��ߦ���9�s$�7��1�B�c�Z��o����h�,1�W
K�L,1�� 1�1�6�ޗ�IIgy+�4��N���!��AWCX�y3�$�ʿ��a���([18�5���Y���##�fr=>K	a=�Gj}��L��q�V<޸�_)@x�lmW�f��#8 ��gI��;�K0:��D�%+��G���2Sq?��->� ��es�&@��h������ay�$���θ��o�%d��c�ca����,#Q
3�lxjv������4u7׹�eC�_q@J�Z��F��zx#E~�>��a�����a�!�r)6z*�?����z5�E.4��~A���x8�w@%(*��$� �4��M��*��/� d�blL��)u�"���#��1�ʤ�HDL�VW$����_m֥c�Б�X�j�L�Y��ۡ�V7II�_�pe�|֕D�)�C=��S�����ߐ�����F�\@qM�Vb#�փ�2�ƣ�F>���T՛8�USC���,�g��������sc�7��3�3]��l����6.됛j-<�_��V�B��I'��褉���V�6�qB���Rg̀���k{�� ��o�#��r�$00�߿�sM�أX$'d��tvƫ��c5G��+.${u�|'�5�'	��/����ְ���:��#i�<a��1 O`]�Vd�(�qLK�pҀ����;oYœ��kWa�����o�C@)���eF����/S�=�A� j�+R�Q�ɔN��zT�+4I ��*�����M��B�u��y�<���	�s�ܔ���pz�7Q��1,�q��%�{���vL�ݾ��j@����1s������$Xz"W���arb�m�) ���W�������� JS;ǜ�P*)�%�M�#'@0#۽޼��6牸~�c�6�=�{O1i��;γ�DGJ��6H�!Y=�"� ����w��?�\�?��=j`������p�b�±:����k�q��h�2��i!�L#�'w'��4PK�٭���ia�����\�?*�J�1�y~������WR��Y�-x� s�_�i��hw��e�4�鿣q��t�]��H)�@�723�}����&
n@�yԥ���&��K���ӎ�d� �(U6IJv�X|�8�P?�!L�k\؁��/�*U��t78���У�.f:0�=�Oj����X�.b�&YL%h����9En:k֋!b��	���3ޅ����R���u侘��瓆�ÉxN�����B�6v *=���%�j��\-ͬ����eau�ۗC�v۫R[s������ǩ�z^���<.�1KYXO��X�y$�b;z�j�qWH������q�E5�D�r�].�KӀhh�������<�|(��QT^:���q�U�?�;���A7��֤�pPN�+�O>��D�l�nF����؅�`
l�!�N�)�§�٬��;�4���F��Aj� "���n�:��:�0�>1���4<���]���aaw�gH�z`GӒ�c��Ұi/|�����%釀$΁���$�XCǠ�]WD���5̻9�K=� �3�e��YU�M�ڗ��Yh��*�?��ꥑ�O�<{�1��9��v������	���/�o����F;�b&�@9#����y'$RZ�chE$�vǩ������X��:�=)n��jp��Bj���b +�M����ì)<H(>��"z�s;2�����rMvl��j����U.h��e���Ҽ�q��w��:3<�i�F�����%�Ɗ���m!)�I��K��C��ɧ|�mQJOυ)_l9o�|d��"ET���e�Dc��FfDg5%�/�O��sN,���f~f�.���GHӯ���I�~$��|Y�r�r*�RDI���S>�R��v ���+X�^��U�Խ���8������oL~����Odϣ�⾄����Xr��p-�胐�d���-к�Y�rʞ4��/�R������K�i�x4�_(ph��8+%s���V�j�q�`�5�P2�\oc���湞�+ �P1��j�fEav��H��<�@��#d�m��n�6^��4:�=��ٛ�1aS�Jc���&,J�=�fo�w�4Ә	 Vnm�B�t1�xP������?�	>6^�h���\�Ωhs�X��s��0��n� �J<���E*��K��HP����!�.�ǜ�;cr� �1z�ׅ�F�˿�Ǫ�x1��n`%���I߫E���ͬ�m"5�J��� �d�l�Wr��R�Vఁ�J1� ݾ�;�/{K�+�y�_BS�U��������?���,~�w���;ޣ�K��)��w������������0�#� �9Ib��6C������S�e�Z���@`�l��ρpRvǸ�`���;�����ɘʩ���w�)��Au�K��b����;�0�1K�z�E���L'9K��G)�#�R����e�Z��|jP[��8�j�1E�R�ƞHΓT�
ì�[�eg�I�U\d�v��v%=5�����3W��7:G�-9��_��¾k�)�QT�<���|��lUF̰QW���l%�����;O�
	���)��� '�͓^[�,)<R�U�[Da��	x%���%���~�/vv.e�+��8�%Jh��
��\R���,�χ"�@I��d�
�(��i��zZ���^44|����c@�����KgX"�~(��Gە�,���_�k5��P��{H�y�����+������t�pKM�˪W� ۔,k�3�5��d���½z��5���=�$�$�ڻ�f�F���������؛�8b��>yu�YZ�zz���*�9�~a��	�3�|:式7u?-�kN*a����|ήG���Zl�`Aj�V�o���E ��G��I��먟ڱ�ד�>[�����X��?��e";-�s�:�EF`Н�w�J֐0���"JO�ו ��~�Lb��4WAEr�	�f�6��M# v��E��"�����i�	���c΀PЯ!b칖�q��|�c�c���nn��7���T�&$#�@���$��Qauĳ�H78#���
�?��Υ�ב��Ө�B��Vҋ�#���r���e^%V*Ʉ���B����X���^�](]P�VW�V�FT��8�򌝞�����NyF��Bh�g�#���os��^�(I�\"���Ƃ�y"5����"�,��:F�x�;�n/�1��g��=�<W���Qm��D��J�.s��X�T4��Y�����P�"��"ѷq9�����i���~�)����@L<W�q!zx�i��Xؓ�;���ЇK�~�w��
�G3�^
"�H���
��g��p;�<��bF�����{l��t}� �q@])��e���-��$�&i��r��+�g	e�9�g��9�ƨ�5��F�@뿎m�F��� L��72��O=&��}Z����Ro��s�}�*Cɭe��n�220qQfW��[
Br�%���۶y��b������vd�w[��:h�,�^!�{���'eH��H�F.'fm�V��u�����a�WՉ����"j!P{0S;�?��^0�B��*F�G�1���¾ dۅ�4&�L/(�#�G�{���U�1R +�ؙ��m���������1Y���j��W�Q�gTtG����i{t:���=6%<ll�Tk݃G����̜��?�Uum��F��*Sx:\�Z�{K�EP��G-�8O�\g8J����:����I[��mi�����]߱3,���^�,����ؽ�أ^��*a���6޾������k�P;��.���R>=��_B��y�x�
�C���o���FlBh���A��j%��}��h|�?�b;���jЇ�<�|ȟ��'�­4����}�V �^w{�a��\*�<jW��r�o��JQ�k��D&�	�[�i*�HUb8�Q�'H.�N/��~�5��&��)�I��7Тkk�
��w�^���$�8�^��.�K.�,y�>��[�1����%.�}�p��$�V��6�n�!���c�D�F����x�����8ـ�Y�z
��\X���Nl�G��Q@@��G�8h7�3���C�0��x�۷2�F�,�Y~+�B��������)~�#��tS��L�_�;-��Q�3���G�pك��A��H����9	��]�P��8�L�<H��p5�{d(�D�M��%�����U"&US��g���F�~�������o��!�}̉z)�"Gح�[2EM���:_�����vQ�0#�	XYꚄ�Q:���5>��J�w9(�Z����s�PM��z�U�F���)
�mJ_�ju�"g�L��K�����Dm+�䑗�by�3~��CgM{�#?�īJ�e�-"��1Y㿼��6��^��䭃\st�Lb0�pȹ&�\�+b��v���>�c\s�`�X�O�c����U������c� T�.BZݵ�Rl��-���x���<8 ��
�ć��XA=s�d8&�β��D�R��9$��i%-�o�+�t�
2�e��o�t�9^~+��n�${_�<�"�5<ނ�w��U��׭�D���U1���$���{;)S�W��g�!LU���ǅמ�'���.��䨠�w�R�����]qB6YE������}����W�����*��T^� �C?g!�E
���/w p¹�"0B@�#�:8�%<�l��J6�)�۸$��(e7_���)�8�8��6C���{`��%Dn��ip��K�Kg�g���xd���@^�X�3#�_���ŷ����b:��7�]��I�mپ#����G�ܕ���,�b5; ���4��߭:�~@=�b���`}<vG��E�]#���03���0I��	��,P��P��3��/���x�{qc^�����U�f�T��Q.�N�jp�k����I[ӊ��v�����ad=�ܢj1�4 �����7�+�~z��pQ�~ �j+�����CC�V�F����W�K���]��9**�/$�e�B�x<$�iAQ����O���伶�2Pm}��G��N��{Gtw�2��DWOJ+d���I�p+�/�����㖕?��?�;���#�7^� |�c\���bu���d?/f�WS�����T8�`�T�h	�{`
zP���� �x�睲�ʣ	�?Xsg�D���i��F+�B��K�(��h�7���Y$.Up5��5�5��1]L/�rz�hbq�uM��ى����C(����pc�<4+!p��>�k�F�Hs��?����$�_��f^q��<o\�א��_ڳ�"�J�oEEd�������&Pi�V<b1R�	w=�,�?�U���JRC���sy�q3�% ��捤CK*���5�{rw
�1E��\�rY���1��6g�����Rh�p��NC6��g=�R���BG&�_N�sP�	p4v0.� ?�E����l2�K⢶�����);�
���d��v�ojEZ�C�B���X����$��SwX?/-��%����EN�����e��.X�J?#�}'����7j�RY�[6�s��g�-j�����^(آ��(Lv��+!$`����~��T�����EW�9�OHvtX|�:��
����t/7bb��ַ�L7�'xs1C�R�S���Rr<����3P>�4.�ҽ���g��^:ˋ�����Il(��Iȡˠch���\��
��[t�:�`��:Ԑ2_n;�I{�Q���u�ҫ���Ry��z��P�]�颃`�������d�v�����D�(��D(y��K���w�����#N���o�L=�������N\w���� �z��g�iIһt����<����C����n�Ns�ep�U��.8��'�'�Dy\[ݟ=��NcqU�k�ܽ:|O��yDf�������\C?٠\�Mtk��M����M�����L���0Lab�?3:�vi������Ƨ�&�|���^�ClD�|jX<k>�EMKL�~�#t�4#疟�w�1�$��",ᄭ/;�Ѷ�Y4� ��%�4@*$ˀ���ًiIK��w���;�f��$
�SE���|��,�,�;���)N��`.���E��䶫�$��eĵqf��v�o)��Q�8�?�����P &$���6�nm��e7��DɃ���	1.�i�.R�XѪ:@շΠ%7�{:��4NO�x��>�p瘧��=K�[��v�� �y� 0�Y�R�B��� D��;���F*;�����AV������N6k�E�����9T����\�\AE�,���Lj ����D5�#ܓ=ޘ����+�yܽ�Ж�qX���ҽ���͆KNi<p���4�������m�$1@�&��](>' �:n��Ee<7-�!������Lb�D��4"�*
��m�&3u�w�ԁ;���As^��J���.m<.�7�)�<��QJod�y�M++ي?Qt���x�n���V�Ǟ�C��_��;3 �'[�`S���P�f&�rk�� J���kZ��,M%�W�u�^/�<ݯ�H_ӏk�|:$���q�	髇0��oSٱf�?'��N�er{ �dИW��&��3-jY�1o����o���L��R��)�߀8]�_�O�C��m4���,e�^�]��ղ0̱���B,��z\�z\�ˁ�떃�2��bo��:�h��G��0P�:�q���4��~ٖ�a���Z�Wf|��'`^cp� �\����O��k�����N5�&�Lc��Ւ�ө�i��\���)���5����t��X��^M�j��v�`pk�]a�#�Z�E��*����Z钺������|L���������7X	�yH���؟�Q}��ĚP��
CS E�32ڭ:���=� hB(��x_JJ�2�0ڨ=�qH2�j�U���`\�b��k�6l�u��E����I��l��H����8�A$�6
����6<�g/�,&�]c��cr�I�,�����@��$ �>ٱj�6W����+�U����<(s���L	�.:�c7�����g���"��� �{VN˘5������������MH٦�u�9��}`�<G�	�t������4՚��ֆ����Bo��wl���:����oҒ_g��E��c	U�j�^j訪+��XD��{�!��O��3Ā�F�Ԭ����F������X�K���OZ�ӓ^�������%5ACC��G:�俌h�A���qXIso�ֺ���w�e�����P��W-�����Y�Z����]8�\Y�̭��G��F�B�$�`�p�"�V_8э���߇Fo�<{f���dYi�g?T�_�X_���C]�To����� ��W 4����-�V�J�K��4�,��V;���$�292t'� �L�~?�������./Ri�,�mT���u (�@W�r�K�X�tHx��J�V�a�б	��� 5'�M��J���K��z��͒�P��'WS���̿�]Y�6?�9۱������/�J'`˦l}��7l1W�/�&��~蠪O�@��ً�����_:����Ae ���8�<%u��V۠�K*I"y�f�ӱ"IU�6?��	�ņR_Z�;$_]�C����˥06���U�a�X�c���3Ӡ�,q=ɋt�V�>|�-r�}Q��p�-�b��go&�N?�]ԁF���%h����5�{���!�'Ӧyj~�� $A��(k��e����=4���3�!dN/+���/���n�oE�}}=�#�c7{�z=��4`Ŧ��Fz�j!k�xċ�
�b5|m�E4��|mVA��	��kYk�(��Ǝ�4xk��[јTB2Y�C˜b�ei۴�A��8�^���Ai�7�M��)�����uT��w)�S���������S�z[�z�?[s/ϧOħ�kڍ���.֚dJ^�cbvD�uw9��^�!���#|��ͷ� ��6���6�����A�#R�_���Ħ}	pdJ�u��?�E��tV��;E������B#�H�p��=R8���$/��f��������h�d�k��������/�;��L!#8�EG������w|M��+�]Wh���a°�a�FR�[u��<�t��Di2�����E�_Ԅ���O̈́ y� �~��vs��g� ��XE�gA�[L' �� ;,81B�'��.�ET6��n,�T/��kwii�Ӛ8��H� �<1���7���E�CW��2�3%���a�)s6&R�i-m���_lQ4t����ܫ�y��H'v�5d�0�ԉ�su��ԟ��``��RT����2�h�&Y0�m��,�v����ڟ+q�����+/� ���o���X��pfz*��Ss�y��Ք��ܙY��K	�K�@�4k"	*��S�]�~s�O�l��`aq��DV�i�nn��x���a
Ee��������{���m��o``$����}+��]�Vn�ҷ)���B�I	@?1��Y�+A.�g�-:���>����;��4܄R�e�I
Z�i1�j���ZG��y�yi��ϭ��Nx�f�ўt��w��g�\�ʆn��HLSd8���t� �b�����g?��4��p���bZO���rWc��z�f� �Ȗp�n(�kf3w�K/���'���+J�깡��"��'��$%�ڦ7���z��D����0[N\�[�����[�IV&�"���Ι��%tё
ic
����m�C+)��Q[����=*�P����0I��.��yKQ�@���'�s�nP���0�V[�yx��g�lьg5~N��$5�\��̓>�B�n��C�g���k�ڃ�`_I1�1	�F����ڜ��~z��d���~���!�k͸�6���� <�;-k,s��zJ� �5��f՟K���)ϰ����$ˎ�.�H�ђP���zgѸ�����Z+��Lփ�����8�vК����紲z���8C����\��aIZ�w,`K�{�#U�VoF��r�ۘ�9����p''G�G�
Ap�ɛ��h���M<���:��T��G_��m��k�����f��=���d$��Bh3��Qp6���73�Ec =��B��ÛM]<CM�A|�3}8\�/%���̊=۳-�����܅����������F����ہ�8�~�м��Wߍ���A���G��j�7 ���9�x�H����.F�=�cch����5]�b���;9��A�魀�ʿ`^G)�������_h^k����I�N��l�+����I�5fq�*�J�m{�����^?�l�l�#��Á�4�S��5k6�,���9��Lb� 1Dv2�|6�}�Yx�>�yD�H6:O����� �8��'4���ŏ��,T��I)���C=�)!�-���Ovd�>U��>+ae���9)�T���'�(�}�� tb�^�t�;�{&��+�ds��ɘ���V�6eF���$t�	p7�c0կw��B3�.��I���&�kss���u?�E�Y݋ʆ�8���ٻ=�dX36��.�H���{$���G��U���ʙ����pK�l
���븭�Z�ضS��M�`��`�������N�p��y�=���:h=͘��xu�\�������􄰛�ńG����h�+�䴢P8��ި?��W�� ��6�8L��[G!��X���P6�0�/���e�k���w����#OD�y�Y��54�1��v�@6�C/� |�HeI���Hg��>��(�F���Kg�V�|kף���3u���7İ��7x[��t��Z��ɨ��������n� ��w�<;-XE�#��-b���S��+އd�����x��p�����_�a@�W=�ˈ����q$

�4�sԅ����w�kO�V`�mz���fe+\�?�r}� =3@n��D
�ĸS��MD���;]�R$�������Ln����F�~��n�ꂍ�b�EY�ׅ4ɂ��s�hC�̞U�f}��z�Wm����g�
��
i�`a֙^�ִ�6ɖ��^�0%r-޺��qb�Nb]WpF94ߚP�z^�2Ǌץ1��B]r��ķ.nG
����r�k������a�eH�dH�+�C��^Q����	0wV�5�����p���Or�}X�ׄ��H�^�;��6`�h�:�v����N�a�͖� 4���7���,�����/�͠T�	�r�{�;�a�'�5#M"��6��h�� �+"�d�)nҫ��o�{�:���A��*(��E ���P�2�uc��V���C�(!,���P3��~��)A�Bhq�k�	��(���b�$��i���
o� ����)��ɻ�xֿpӂ�yXX��Dp��
T/Z����Z��٣��j��?+m�<N�>N��D�w��ͯ��(O�#�T�F�ø�J�Jn�����=r��r�/���.�sc7�b�� "�]ug�%k������n������l:��Pqd3Kgn:8�}̋�R%U�)��c�	x�=3�� e�wN0�Ma�I��Ii&�;}LfAOƭ;�]�_����s�I�w��"k�	���z��+�Nt?UKYK!D.�|qdc~��[���1�Td��r��v��ŵZ�N�<C��dHR$j��)��F�u��d��D}':�����j��e�\^Ռ�9O��j�

W�+t��*^*�dd�E��V����_���+�W�����C���>�Lk��Y��
b��Q�<;��ʾ�s������տ!9�կ�م�Df�e$�h)>��n�"� �Y��;K>�Q���Mv��
X���m��y�=m�>��Wwh�� �W&�;ۏ;,U��q�W�n���H�W�'���H,�R�3ߣ�B�}!�^�\N����Y�N�`� ���l�z������"�P�
��U�&'f7�֡-U��f�ޛ
PI����U��	4o�D�BRVc�Wh����>�C��;<���?a��X*kÓ����� �,p�\<��v�ޚ=�W�+G�`v���t�pF~˨)eg����%gw�F(�tu��h��H��_�ih����	�������1���^�$�_�K+(�$�	��hK!f%:���4�#/��X���^õ�Q����%N$��b�������2l �o�'��gɱ�Kn�V�֙S1��t�p�h�������܅�G)*C,ׯ��m<��|y�س���!�e}� 7tc�LX�ӷ5r��v��^�lh`9����I@�\�_?��1���铁ۀF�M���B��	������g��{<�������yXM�B���5��qa������ ���C�YL��dd�_7�����a'6I���"�C�^��9h���Qn��p6r���K"s܀eCI�%�a�fX���gi��<
��/�|$�}���_:��
z��8ޖ��Q���Ɣ]��Upv�$�����;D��,���A�H{�8�Tp��H��p�<��|WiY;�e4���X-�����U\۟�/ȣ^	���U��39W�Ϥ�l(�gq gK"����}
Á�#�!K�4Z�N.��� jQ����#��	<ʐX��1��x�K=�틳[��X�H<��N�)�?��K:�H��<X=a(s�|]��j_�@�U��c��i"��d8�$̨�������1�(���ර�,nΠ��_x���V���2/�L�M��*�����P����p���1tm���d���,�k�a �%ZW�p��mwͥ���t�1{�����5�U3"�-�3
�&֬zS�t�͉�l
�"�j�y�R�D�?ա�R�'����U�9�pe�=k�L��	4���姓9�}É�j+���pӕ�]t�q�0L�CT`��
|�@ItQHhY������mX8��;��7�=�����nd���vX5��:�q �=�����O�ÕC���t�a4���z�?�+�r�E�̸v����c���_&�
��k��)�ۣ�!9J�6K�'����3?�$�;����<}��51�2�7����C��F}!uR�iwC��X�w�����e"�=*_�񭾽-���֓g`�����Q�p�`��jC����К�������e�q�2Kl[>\�ܯ݊�S_��"���R�;�.p���X �l��+�Cq��QX�`W�(n�����-�g�3��)��'��nu�ODu2
�T�\�d�˸yfw>j�Րt�ѥ�����M�x�O{[xH'��sp�ȍݤ�����.��?����>vD��<"�~&8�J�,����6-��gr>"��;�,?#�ʥk�S�Q	w���;��X�@$�贱�2@d���A�,dK�s>uZ1��q/LO]�MZO���i�h��X$k��w�2&�<���Ef1C}k��Ι�%��F�}����B�k�������_��$lFZBBl���b��y
9-�:�i��a�7�W"l�q�w�@U��Ş��Y��� C��mayD҄fT͊,$���spS��>i���H_nX�&K\S���������L��Mf��s�s�^�}/��g_���L�x����i�L���(J�( ^R��R�c�fWJ����]���*����`�/QL�6V1
'�� )&����p�2 f��7{� �w|�F�/�
�����a���x������ ���g��@�b�O~�6����h&���w�Vk\�\ꇱ�����{R7p���[��G����:�FF9�)�Md��K �E�aΫ���pY>7��:j�e�����%	_Hi����5����m �G�#kI8�P՞C��^�_�i�ڳ���;��������g�� �V�!.ӱ�%s�K��#����F�4��~�3�UW}����#��@�!Ed�^����洞YPƕ�$���9�t�<��*�ӛ0�1Dq��������o��Tw8!��/"D����^�f�V
A@J_,^7���[9y���y����r\qN�.��/x��<Lq��.3�`C�OH��)̨�x�2�q-�g�ׅ�ԻO/�@��-c?kb�2D@���.��E�HX!�n�ĵ5�mq�9��Ŗ�ˍX7@��y��[x�U�쒻�vP;�&ɹvg�s�C�K��y=1��1g��&1��]=�.�5�?��P���V~��O�>*�׿n8�,s������sv��y]n���b7�U���vr�(`�',X��.=�T�)Bc�Z�r-=�wd����>��*$d��Y`�,�e%��O,������'А���)�q���S3)��`Ě-�Ѭ��ҌRr�3��ó��bd���G9�&�{%�*��ܶ����X�a���'"n��ZQ���0�}�¾�ő�lz"e�������;C����έ�H� ���j&���SИ��L'Ȋ�y���|�g�#_��W�>����*�QN��;uIG�.qkC/m-�N<)$���j��S.6��w J>����tC�TU��WvHG&G�[H����8ƒzk㍇�Di
N0._�j�U��U�a�%��H�oQ�"څ���������7�G�fA�/��ef�!x1M5�pKE�˨5��b��i6[���[Q�b�c�_P�(y�tv�����%�LShT�=����5~%�g�]��ڢ3��^�U ��<���d5��C�Lϑ�V�	�ώ����J�T"h��8,aC�J LӶ�)ŵ��ϯ
���+rQ�:�4=��3Z BK��s��mJ��Ҷ��a%?#�Nh�Whl���%�!��`������N_��&��|�GŰ��ঢ�a;WO��fWa��:�R_�?dE4������yNd��P<v����x�?�˚�ZK��]t�m�u�7	i��rI,��y���+�Z0�V�o�>��*�(Pg�4O�r?�G�P����[}'�h�Kh7��թ:OeP��\]-�9YdBHݿ��,K���Mļ�E?�2�3}�:G�����P���<�ƴ�};I�µK4���,4pr.��&jYF���!υ+`q�c{�����XIM0kX/U'���]\:@S���B$I�&(bk]߿���W�eH@���	V�e���U�,r��g!t�\:s�p�2�~����E�|0�HD2%�T�5#b��Hb�]9���%���4x@h'�JVn�E����ʏH���y�M�)��;_��R1;s���G��`�M ��T�1:{n���>1V��CB=Ɍ�B�w�2��}��5)�>����W��x���d��w[3z\�X���1B^t3S���Ԙճ3��vK����y���mɬ��ӿ�1U��}*���-��(�!5�� �)[K���f��[�+uZ�"����x��(�̈́����ot�u����Y_u�`����P&��|����󑴡* �K�h��gń������wz�|�l؟T\2#8��w�Y�w�K�۸ī��K,��6YC:���I��������Ra5�gU��%���8I�!)�w%8Pw	_�RJ�/���?���dW�ۑ���%f	L	4w�TL�G][#ݸ����v����ţ����(c���

�1�A���r���H��lu|�_h�bx?��a!awR+�^�,� {^��7�	UJ����ϙ�j5oShn�@k�!OY #�
��`[!"7�J¢�'j�Ò.pA�0�9y�ҿ`x�����à�8@�ŀjV���Q��#�
��bQ��~%#p���ʰ�����c�O�ʒM 䓼k�v]!�E���{��w!�7q�~��b�,n�F�?-Ux��d��(Am�3-�����>�諭��병"�>�_oE������E aO���fo�1ž�`�a�!�9������F�x�������)C��~O���"���"�)AB�����eŹ5o���O�0��9E�xz�^�{�HMp���=k_S	��*�I��)W�VG^����i����^{K7�y"���iޡ�/cπ9F�D�ק���E���b���Ie�8%;�!�Ƨ�݃圝iiJL�X�!>�sݼ�Cx���Z�"��!7�I���x,\���QS�&
���|?4���8	k��o ��[c�%�E-��Gˀ���lX�������e=t�n5;�|V����⣎���A�s쵶��!���ݍ��03s�=���Y��j�T��a��릵gJ��N���U�e@�Z��❣C�|꣞�`֗�-��6�����7���� ��ً��|l0-'f�|�x��z���[-�_ʲ����&4b�w�h��ń(q*`�����0�u��iNw��B$�0޵��;/Dͷ@�S����.CI	p�)�)��*������c^��u���9o��$dKG��59�`�����G�JmpT�<<��O-u�@��ۺ0a=��B�b���I���#0[���s�x!Ó��k�+3_�M8�/Ƈ=<��?�	�6�y$��SmHY����o�zz*`�)�����^��ݘ�^pSvò�u�?�~r^<�?,�Ŕ��Χ�,: ̡�T�����o%�����G�}^˯Y�h���2���Q��Ƃ:I@)�$�C5*�yM?"e�]���]doJ�uiJ5?{d�4R�nd�Q��y�^5(���70�0m���a�>�G��qDK�{�����T�4 1�4�F�=���K\��t��
��ѥ��p>�#L�ǅ�&�?�ABU���/w�iR��D"�h��?%��M�v�����QzOنu����2п"E
��س�ި��i5?�E'��p"���p3s���s�~��c1����k�w�3�*�ա��m���Ү�9��$d_��`��`��e#�/��>e�:g���$��F�8��{z�J꙰�k���z����*���]J���kZ�d�ԟ��"����N��a��^<!Kk���#�+��=[ZSiW`�O$\�Z��w�|�m�A�#��A�Ns?,����@]}o��M�#����K������)����I�ə�d���wea't�)�yYT	m0 8_�e!s�=9��\��4`�fԋ�9[�)�!�K��s[mGy/s(>Kv6m�vJ��3܊�[	��9�����9 �=H�	.S(�J����oV�o�xP��z)�a(����mH ���B*GR�(��[r�/�N�g\�OZ�cf��8+�|���og�cG����f��u�$GWc�v�wF̸�M�������:����a���֓�!�����f�>w+�3��/!/��Ͻ�c1Ν92�&B��Y�j�L_�%/��|��F�}͇��.#Ӏ���p^P��_eAq���H=D4���:}��`��>l`K�p^��!�nųNO$��n!�2��@�?��7a�]��T;�X�k����Z
�[9��e��ƇJ�0���\F���g�����/N�p}j�6x~��&z��=?�Zk$D��1�W�Kz|������y���晟�m�+A���s��`��ls�jܭ��b�c����ǡ��d�����|�q�Иf�P��V�su�oD8ה�OrK �$�{ �-&�viM5�d9�ݧ��AZ2�O������Ј�mL�
������
�F�n�[����.]b�~�LI�6m��%��:	�N�r�*aF�K릑G�AӒ�3Ґ� ��Qc)m�3W������uJ,{' �&��ئ�lg�N]���/Ɋ�~�<����tyL�*�Ti�_�t�J���L��	�h�R�vF�G��Mܣw�၅����ހʃ|"��	����ڜ+����:Ri����ئ`zVj-�H��;��[)5�{I�Fa.�����<_`�D�v=�Ż%�`��3r'nn:�A(���Φ��KNB�D��2y�K�.���E�����H�ɑVZs�Gا�,��]��3�z/i ������/|���n��Io�L]l�+V~��ۑMRX���Tn�J�@�r:٠��Z��*�����]�cP]ip:��Q-{�O�F�f��
�9a��l5ז�`oas=O�_!288(QP�.��1��1�0�F�i�.��l dP+�O�";���������\������b)�nZ_Y����@vo� �q��fO;�r�k8��!�ĺ�P%�E��͕w�kP����GL�;o�ľ�ߘF�Oa��.x-8�P0���8��YFR�_�y�AP��cha.p~�oKDP����4p�(��'H[F:W��.��F��/��1�mĊ�N�!̜�*|�$\%��d��D�1Ս�.'4��M|2�9O��^.��nws�hh���"¶j�6qţ-�k��!BiX�w&��`�a�H-kf� =6����Lֳ�T���|89��]�	V��Z�� G�������ص�0О�ĳ���3�<��{��K��aY�f#�a�CQ��l��2E	�Z���OB�!&e�rj&����y��	7�⠖�^����U&j�8���>}�-6�eOU��qs�������PD��n������?�%�@�i��G��'��j���D����J�^?��t*.��mg��>ا���T�D��v�<7�U� �Y���ϫ��J�����͕h��4O�O�������!�����l� |/��DͶ��O�:F��EO6�Nr�u�湀����q��)���l
?��
ݽS�Yu�7�^G�Mj�
�T��E��炖e�e�H�>)�w�{~�	v���p�sد^���n�n��Х���{n�i�)�3��|��e��fH�<�莽�h��c�b�j2�3��`�~7��So�Al6W�5�AWp�em,��@Lܴ��q��z�I㩬�RYXƀx�w�(��tޜ���q��#J2�!��.�Q�l��m�s�x����m��'�䡥/�ڥ����X���'�����d���LL[�����' �K3���IA���l�yk�s9�}����۱4��ձH�P��]]�9z�;˽w�Ra��g�3$��b:A�����'*��r�[xn��^�<����x�("es)��)�)��]��
cA����_Ox�م=e~Q�+��j�o�Zr���/�kca�F5x	;�ʱl��N����P+ �~�]\P�'MB �Υ(����CoU_���t�?O�h��̘S9�_Hb������p��]����[�Ė��a���"�?i��ʢ�2� ���f��u�z����EV��;�/�I#�n��Ԟ`�d�.66iS)ipǎc[|�"J�a�r��$� hF�qQ���U�-_��!	 �yW`fe�mU�:c��"����{^ m�,N���t��j�rK��j
�2��`W �˦]4���d7mZ>��
��9��vh��0C0Ї��?$�^Õa�����+�H�ǺbR{J��#�N�#��|T`c���:���ԁܕ#���g�L8N̲�B�����N�T1�O��S$�L��C/��T��-s�t��D��f-m�j��U��H�g��ܬ;b�НJrh�����d�4,����o�cW	T3J�X��oG���o�d�Ɨh�^a��B�����m���~)'i�E��N���~�����K��D=M��b������)�#ǸOP!Z������IU��X�vM�ɀ�
��W���u{*��ԝli�Z���%�����%f�#mT�����U�:�����-���2$���w"�W���a�$a���J�\%�+4b2/G�nvmm9�"����~A޳��� �8F3��M_��]���-dv��$��Dc�(洩��mm���:wi��X��b�@�*ȹ
y�m3�G� �	�u�|�����\����Z�^���'Q�LKt/�-�tю�Y���|eG4y�,�y[��J���z�U��������o�a�>�P�+x�km��g����
�0^�0�Ze��s���q�l����+�j���J�XP�~N"��E0�5����ꛟt|�b`��������ΰM� &�c�yH�:�.�V��lF�2���d���/�d�p,0�|�t˽9��ym�&X��?�E��1܄���5�vŝ댏S��Ny��t��60��g�Q�v� ��_���T��T]G�tܶ�b����J�^�Ɨ�e>}NUv��>�re��3eY�R�'Ewl��B����M ������/Woe���E*H��Q/D����B�{�F~��񋩿�����۸��r%xTL��OןyPM4�A�jRZ0S"�#E�9��aue��%~��'�O�;�SZ�ƽR��M4axd���6�����˙2�]w��u�˜`9G����R��ܟ̴O�o��z���jpl"�N�7h�{�W�o���>���ު��90�OG0ޱ����LS5v8V���.�5���7Ҡ�h�16B��Sah�w�ؽؽ����% ��(H��Q=���\��ih�02�ژsoUè�5RÕ������<��&#,U�*>28���HSd�i��̀?���[eT<������W�ޫ���\	����yi�d���:e�}-���&�~?+4j��5F9�	�(%
���3���ֿ�k1�ӎ��;�m�	7oƊ�b.Tb��������p��&u�U����d��ɢ=�8��r Ur<�0P��"o!���v�HM�JrLb)ۃԣx૵ Z�ͷ*��q��c"�F����t�4��FS�mi�S���X��f۽�f�خ5i�7��jm��Z��D�\O:�`�h� Щ*6��{5��Y�PX��0<�8+�n�RY����'>쯏��n���HD �q}y�����IzU�f޼�`�#,�W�eg3@++ޯ`��z��N�h�k��i���T�(���tLG��S�ئǋ�6<5/�c�*�_?��b�ݪ�#���@��0�e�8A�e���]�.S��yn�gS���-������<�ގ��`�f�w6^{���Gg���l.�j�yyg`g4�%�#���:ZR
��0M2��w��v����I�V�,R�O��j�5�2}%{��$��JhO73iA�F���x�䐛�Ums����5��~�,m�����.��� ��/�>�Lb3��qJ/��+
H۝<�E������e),K�!?���3C��jq�w��9����*U��w��4�1���4�����m
W�Ǆ=�t�97Z��4�9E�#�x3z��ɸ���IA�GJ�����Ⲿ�'[��]��% [Hz�O�AN���Y�S&�^v<%�J|�����*&RW�7m�Q,I�s�a��o9}���z&��q�+�A�c��?��՛���"�;����t�_jA�Wcs�zY*:w���8oe����ь�u؜�p��#	�fkc>uy�T�Z-|�=�J�RF"�B'	�XvG@%������؈+0`�{ D�'�l~R_�cn�0��}!U��
�vv!�w���ց�T�!�E�}�Í�(dfΛ�oP��:P4��C���0�8#�$wb*��y�񟣍�`�%�[��R%)����렠^�� �̘����Q@3Ӹ��&Se�:z%!!�i��l�
k�2@`�6��@0����$2�^ڀ�G���f}�PB�d(�-(�DQj���d��&�#-��K��!?���÷�T.?�wՏ����5�Z���CX-[TڂL� �� F���~Q�1���)�3n�5�o���kdf�n���<[�tR"��HdJ��5vT/(�Lɵ 3	^�$(?�G���=�c���3E�c	�x��$�>��X֕���&QX��J�������MH�MP�h����Ed��	�s��οI8o�ɗ�h+�1��
_1o��3��W���3�
e�	E�����اZ>�p���mz��YCG��-����_�j��!k�ߖ�L�"��T�&��tԉ�5����l��&U �,�aWT�^}�
���OQ���a���eB�X۱z�'�������p�h&g�w���{�a����I��q��8	n�~�p�[�1����A0₽M�g��6M�xL�m��y�T��}nEW���xk�J�&')��m�^��$ƪ�2�NCm�:�S
�1�ޛ�۔4�q��\]���_Ӕ�Iu`	�[�d���U
zoP�Ŏl*b���[��Y��41��G%�=�*�&Ʉ� p��8��sÏ������~��E�^[BmsK䗷�E�+���&����+�~B�0g�CviΞ��E�.N�H��P����do'�	�ւ�[$��g���V�I֣�o��4��%�a s2� ���D%��S$���Oc	f�W�[��U�^��n������DclPΏ��`�*�.�~�"lz�����*��F����@S��=k.k�'�l/;}��p�`����^le���P�-Mr(�[����W���-�yKc�g�A�x67�L��zk���9��c:ř3�"��ɀQ/�9��ku��L��Nl�ք��2V��]�5�tjeWPµG.�u�@K��Kwm��7z(��?$�f��P��^>�0b����V�5o��Y
��M��E�����v�R��p�QI�G~��;��oP��'$�a�9i|�_�QE���+�.���+�u����=R܈��<�}������c�#���X����Ly��~���d#�ˬx��%f2v��'�t`A{���b!;?���ւ��DA5Υ����.�ш�7~Ӿ��KI��|�P�$B+ja$�	������xS��KK�}��!.jIy	�{r4���]n�3����z�_V���<��+�&ܢU#�6�اO�؆�*��#����!�􄇬��'�b�7�2
_�>��^��tA�g8��=)�}G�`U�x�v<����#�%�xWЏ�X%�����-���T�����@)|I��Ԏ�t�9Wf��k/�h�p�N6TI�TY�@ o��Z3�n��Z�P�Q u����7��oZPF"j;r�7|������~���� �cVd��0��(^�����K����ΤC���5�.�LeSZדn)E@��D2�"�XS�2�����5�J��>���*]�l|�Zs��8jğ��QP�=`�7���g����a��L�.]��K�Β��.��Ts���Bנ�'ծ��j�����P�:*��f�y��	5�g��+ڜ�R?�sì䨞�w�"l����ha�1�p8�3yWEI*�O�����x�e7�>L^Ut�q��>�� $�}��%�A�=��_�Hch���ۙ�{� p��l��̯mS�_X�=v��N�=�g�+	/��Z�,,5e�n5jR$TD�z��H]uFX�t�o�ů߇�)��i�@���CҤ����\�:�eؔepۋ���?�Wxf�z4�p�x��;F�ܝW4�8��HκG��J�][��W�������9y(x�3�G�(���x2Vd�������i���c4�S�ɚ�F<���Q+ֆBvm�!����{����n@G��#j\JT�����=���E�	���ƥ>�Om�R�� D��],6�\��:~  �L2�n��d���q�RB}���V���F�֜��>ѫ��QA����}%��7��;�����i��=�ʘ�'ߓa5_QƼ�G"���`i_[l�k�L�Ȩ�-!��j����̳J%�P�u�hCQ�2�V*fyo���G���$�"��t��n�7���L����J\H����1�us��R�U�C�K����,�^Hl����$(����I��e_H:��RE�T�������u��O?�1�V��z��� �Ntg�-�������@x�N��S�0$�����|C���(6�ט�"+��c����3|���0Rá�����ɐ��Y��W��m=���5c�D�g�p>�kƝgx�XA�`���P{ �N���X�FJ!"�_��M��{��+��b�V� �G���>�ȏɘ����4'��g��ܼ�/����S6�7�H����P���v�#��5�&N�)�9rz��ڭ����*�����ɟsL���`����0Kԫ��M��+�0��W�;��7D.��*��M���V�������z��u�!ؖ�R�2i}��T�7�z�T[fU���j6ݠ�2�MC���Q�A���n���	ү��2�p>�xOЉ�{�Z��Af�+���|��$i�{Z?G�da�$y���?����/@/�cȀ�z�:�R������],po1$˾�zUT'���e+�hc��j�u2����%��09�{�����L�'	
�BR}�e�s����9�h�]�e�������q+�-����!�]T1#nc����oܔ_g��P��֒P��P۴�M�����(���<$v�5���,C�e2h��U�OG����?0E�=C�Ww�y�se��W���!T&��NT�+ .�\�31r�xQ��?!�*��� ��V�?&rj�/SM�.��?j���f�N�sa����JYژL�cy�����R�'����c-�6����Vp�n�c���x(�?�g�p
�dp��و{Q���4��pW�ŵ-@��Q�T����4}�� #D
����߳8�+a�(߅h�l2Xm!ɦ-���1�T��v�-ճ@$�=L�,�����>ˡ0���q��.�|`�c��*;�V'�n{�'n�'�{Bw��p5��߰m�\����Ͱzt�����7��=�%��wuxsf����
�P�[I�������"Ѕ(������B��d�v�n����Y,�2p��2���4�?l0WЛ����v��Py�D��tOŕ9�|��U��[�>u�>$�(�.3��j'�۬72:�S�}��>�nQ�?��K�H�Y4�I�j�@����Yej[!��!��
�Ò�{T�gu�t(��`H��Ƈ� T��������h�>����e��9��=G�z�W�`�f�d#�J�f4P˺�����7y��JX_FN(�(2L��]�6p�6'�.��?Rk��^�R(M怺u�z�& ����֢ҙ��}���M� �sBI��kM�n�������+|t��mp�D,�ˊ��� [|���UVspl^�b�.}��b�Ibow\1���p�Fç�)T])+7րC��<�������A�u��h1�	����%/�*��0��!�.�ib��	��pPb�h�ߤ�+`*:�f2�8V��w�:SX��B��v�n)~^H����FY�����l_�s}�`��v��Q�j�^\%9�ʤ�c�E�X�B���z�$36<~��&>q�L��JE��}am����n������̃]
��*f6M| �J�{��f�|�aͲ(��D1��#^�v�!w�,�K֘�"�v���63M'�<��h��H�?��η�T6<MS��K���� ����X�J I8�hјR����͝2��q>��Q�3�D]�e"��1��P-��P&��"�K_��e�����B��ܛL�a|i ��n�77�݇T���V��ǅ����EgHY4_;�)���)�p2������Q��dFΦK�\`����u�u�QM��v���4-�i��Ǧ���y���(�Ofw��_�A�Ê"��Q镛�&�R�B�$�K��Rʳ�D0�8�����h��Z�4�)���qи��k�J2q��イ���)MD*(�e|���F������ѽ7��n��n����&g�U�hB�����/�0�)�5?/)���C�����p{IQxQ��8���D]�À�X�a��z�By���õ��\;}^c�I�8�A��=Kz�� :�����s�AW_�'�1/��?-<x&x�i����(#�ԛ�tj����E�%�G�wo�E��m`�[��"���7`ߐ�?w�1���G=|����|~�7&nբO����2�Wao��R��������1��������4,ӱ����z����rjg?���Ͷ~q��JO���եY�(�qJJCX���M�%4�xz��S��*,��b�jP�{㔴m������UՑ%п�c*t��`{�l ����l	�����\X�кw`��4�z��)��.���Jg�Q��hxٳ�ܥ�Y�%��B5�su�zX���0�,b��-��׫{�ޠU� �H���[�|1dk����8o��|߉�-�_`�rn{�čE���Ԧ&L�g��K5����C�;k�o?�͂���,�`��?31�؝;)ܯO)b�/+�P��S1=��>6���y�J%4�M��>-�[��a�H���a��r*?g׀e��KUݴ��{�6�c�?mģjE+�S���+?Ρ;��M�c���mI�R�Xiv�GiQ�}*M�4�潤�f"�,��c�T�r�n��Ӫ�ü�� "m�8=��U��yȜ����t������ ���3	��º�.���ք���ҩ{�x�b���L�g����L㫌���ꪴTjɠ��kJ�*��T,f�U���|M�w���R�M=nÕ��J�xx�N�� �"�gT�S��Q�/�-L@&}$���u3�̀��T�0��AP`=��12c��bˍ��S}��� i�����%��7��{W��pR��B�Œj{P�I�O{=bvg �{����P��r��u$�--E%�4�0���L�o#�,�?��0�EIV�Ə�@��M�O�i�*C�1;+G�RE ΄YYr�#ǭ|���]��	&�O$��E���9���ڛ_�'��Cw��\½��*���Tn��+z$�itw���@p\C*Q�diz�[#�|Mx�>�Mf���������qOk�S2��å[��
����m׃K�=c0w�-�=d�Ȃ:�(x�A2���[QQ]6A��
-!��wv�v���ê����طZ���w ���{��X!$�vbfB(Q�Q)��x�t�
�8f`�_'�[�0�9��H��!�+@⸁� ߹|��nt���/�����gE��(�҆A^����(�����E�S��cuO="���`���U��|�'6�z.RD�"m
�a�u���r�hA�t�v;/�W:���&*P�ǝ�7)�[�����> ;�l�.���&�I�2�]!,��4��)̢�~��"��[&�E°�8^$1Zƾ��,����yU#��k'ǕЏ�&�F�W��b.�}A� s�w4ۥ/�3@O����>�e��rdKg@��ܛ�bO��dkPe��/�(�X�z�e����*��ä����V�5տ]�I�BB˂#��/��t+/�\��QKZ�۶�<�Į�J�BA�S��Y������}����
���Ȅ��b��+��Ť���^����^�ĺ��#0ɶ^��k��}!p?w��gwrp��f��gi��9�&R�5Dt��sF�E�"�X�:�+�AS��.U2dȹוu��>&DGZ�7uW��+V���Q,��8�����&?d�ZqE��q��<����G҂�<ޯ��?)�� l%P/�3�f�lXR�.Ǥ^ʼ��a�+m�{�<�\��S�9/��)��ѣV3�Rvpo?E�/ETU��	g�K�'��M���
Hb���VB�&ȏ��g�z���	�7�4�f>�yδ�$Y��u�ޞ���(�����H�5J.O�[����G���(u��$#B)��t�wmZ��o��%aܧ�x�r�������㐠�ec��Q��i���bJ�Q���V�����T��ǈj�0�)F���ӣ�`��Y���^�KJ/_�8P�;��[tlZ{��	��V�nX�moj���4�ev��qG�=.#-:9���Ub������Io�K������h�[�5���c��Q��8��\@�FP��a3N@�}$��o���k�w�P�}]�����c�`�UyBj��6���Y���|�vL3)� �{~�q6�^z0��O+�i9)�ӢyJ4�͙hɻ�y�F�x�J�)8�ڂ��l��L���|գ7�E���o��N���q�f�e(�^N �ј)� ϧc&�=s���6d
 �!Q�	��7ޖW���A�k8���7����> ���I� u����I��-f���@��H��Qk�^>x�o8&6��ZX(]΀,p�{�9��Ih�W���8��DU5	�c��	�����'�Y
b"])���PʒQcZ��"��%:˿,��2c!���H��!0@S\U:�I�w ���?��3%��lV��O�/d���1�VcdH/=��j��n?���u�v�Ւ
���S�4�z���_�"VVcf��4�6�7w�3t�=N���2���U1�R��F�?�ԣOK��FA2E����i!�c�Eܴ�Сs ��C"pA�5�� 1Hp�ThO�ܾ�^��\~]��&��g�BE�
�.lh�j�A�,����N9l�pqg�j/U���" �ʜ�)AN�Z��]����U`:��Սx_0�9~��u)z �D:�d�k|{LJ�UK���L��R���{&'}�+i9:s��������fc�[�m���/úН��_* �\ț�����}�ʘ
:����:���H��MvF�@�)�H����^uo�t7��&GP��q���c�8e5Q��훻�:���&;)_�y�r@Փ���1��z%m�)1��_/��u #Ơ4��:�N���X��^SL�qJ�O���`�+t��w/�>,FW�g��	R49Oe���]��:T�M`�����hʢ~�����Z�͒�.�%����k�
�'���,��Xz�`@������|F�8���gN����X�G���߮�e�8���S�V�����f0 N�ʋ�ԋ�t�fŨX��@�3T=PP��M��S�����u��ӝ��lg�*��zP	I�.�][��l��"0���T��Ȝ�h��#K�����^'-Kq����+�ιGeh�U�L��ʎ���V
�	4Ȫ���A�Rt�&�
x RY��c	�=��Qx��Xj,�W�G ֤����߉���,72�C�m�*i�n�N�M�]H�9�A�p}T���]P�"��d"�E�j�ܐH	P���N��k�3�f�*��=l�9?�]���B7J��fdd��]�������\+ak�l)��P�t�q����j��@�Q�� 0�f��r��1�(�̦^[r�t�0��w;�<�E�h���#�����2�����k{����Q�ƨL�gcݨ-��8��=��Ϫb D��z�]�	Y�-�Gh�����Йv�Chdt�9���ak
M��&���	���_v=t����*`�,��d�V٭~G����'8�5���7jw�Y��"#> *��[|��E@��(4����y[=�B���ܠ������E"��B����I��b����rꖐ7��k���i�P$�N����H�]O��xy�X���,$o�g�@�&YL�I��C��l��ߝa;�j�z���&`cw(.��#"��7R�	D�1���χj8~U4�c���Q���r)�:L�'5���)֣�n�|�&6NÇ�B<_X�o��!���ȼ!J�'tn�lt��_��2�����k����v�_�I��
���0��m��X�V�MIJ̊z��2ko8��>Dq�=1���Z��GsV������z�-d��ñ��eu*���0�f�f�7�D��W������u�n���.�>�F�TtN8W��U؉�θ��=�(���=�@�m�_�
w�#6�WfF~��'�|A����7������W�?`���w�ۘM>�d�Y���8w��/�;�[0���s/�-HI��5m�����!gm5ə� ��]>;'��˰�����+���?����T+$j��lN�dxh���2�v�,�`M�X�i>��?�<??C�<d���3'$|��3�p��啧�O�O���p��)y�����^L�d��)��:k��}�V��)�~S �u�D��ע��"�(�n�����c�WVT�'%W�{�7+����N^�#;U����:�>
Q��&�c��m5"����Ύk��0G�Ã�:�
��Cs��]��V��Ѐ!������7��r�l�c˨EߺD��m��m�t���ص��r`�g�뱧s�g�i^�@%�������й) c�F�K-���X��R#5�;t��S}���Qz���'@smF���|�s�_�#�ګ.+�BgHu{���C��O���a��Ք��Q/g�$+#���s��M�_��Qͬ�����$���*��vZدg΍�/q+��܅&6l �q^�w��'� �{'͹���=��P =��;͙f>q��>u����hq̖�7-e�˥ ��:	Dx9��$��ώ���$+���x�k%�ǂ<	f�k~֠R��s�Z='ڒ�zQ�,M(<7�[�8��̊�Y#=EM����B7��d���B� bG��XI�%!�<Q�mp�w�iI]O�h��^EK�Lp��<o*������iM��T����	I&�G������ �H?	��ôqh*+�=+���b6��'%�m�׏׮�x�^�Z���Σ�6m�z�z����؋0�O�$�����K!���!�0lʜ��)�ǈ��-�=ԑ5���>�h�����t'Xz��������%��߅3Cl�u��U2dw%�\V���o�=m��z>���-1�U�����>LG<��9�Qtc�6Ƕ�	h**�6Z$nF����L�g0����[X0��]��35>"7����� �1���Un��Y���hׅD��f9�����U��g6�6��,��d��rқ�g�i�:��[�a��D�T��$�E����%��[m�� ^�򢟲�F*��A��2m=�;q�F������#�I�Szp�Z#�D�n�~��P�v��5�o�m��1�*\��.l��M���jܦ�b�rX���֖�}��\��1'�	?Ͷ�EV�5���ݾ� g�1��U=�w�Yd�*�����+D4_}5=�>0��]&=�gl���.;�NԀ8^�NkM��
s�쓼X�3�j&;$���z扭<G�����b��~��4�+B�M��	n��l�mJ6�:v��o����L������+�1��n����Nɿ��`�Tp4Q����v\ot�n�7W`�ү������|�cy'9�!eP����1�_=�H{�b�N4��^�|v�c.�^tɔ�1��Ex CoO�pE�nD��nA;:de+a�'������+�� 3����c8��/<�vb���gw0���3�
�(��|��䑢�4��Cn�h,�Zc�܈�/Gi&"/@@[G��{Y�oJڀ%P�(�\��'<��9R��B����*�l-�^M�?�ugl��ٰ{���o�g�?!���Խ��ɷD`�??�#�_j�/僞�*r��O2YF�S�FMF/�������5*-?��zӂ��rI��w�cy�0�nI�����B��ڸ����Ѫ1ݝ�`���@�H2�c'���:��dCZ(�j�)�A�W(���B����\t�;,h95|o:��+i�� ��1����S�ҹM�/ܚk�
�w���6CPї�p]zS?T�]�#�x� ��k�R��t���;�{�{����g{� lJ��w-o�\n$EpM|`悢���b���v��J��� Ne!��a��(���y��.�ڀ��vsR�Ϳ)@N����,�3�Vg~0꜔Z�1#�v��M�Q���&�"�?zŦ�丆��@uG��{ؾ�k(�K�*|p�9�v!���v���R�I�\�@>0�@���(D��%��6h��2`��>�����P��O��%Y|�e���!�e�K����}봵zN[E�UK�0�Q��n�_pa�\B=6L��ǯ�[��R����.&x��C��$����9!wEe��b�"��WO��m6��A�F�E!g�XHQ3y�K�^j�9T.e�|}�U/�nT��;4���Î�ĳ�5��$���xr���;7\����tgr�ِ�9E�G���Q��:�Fs5]�K+�4n+�sjUQ9�!oK�ى'�� C]Q�+j����mR?h"ٲ�ϧ,f���mQ�=P2V@����������X�ǰhzL����C�>����7ߢ?�;*����ݹ�La�Q��������'��f@0Ť�6�h���h��K�KE�mbܬX;Rn����k'�09��18��ւ���z7�_�y��0�&L���g�ߵ�fd����i^�8L=$U5l0�EU�0o]�8H)�sS~�s���xU�,�C�α��!�L&�|'��&�T4��@��K�D����C��21WN�+
��h���}=>����|y�XT���� MiI�%�L��=;9g<�Hh�] XY5j,+����#��Q�y��8W�jcW�d��^;�]��+I�
�*�K1��X��?��;1�Zi��	�7�@s�|��p��5���8��� ����W�`r#^R!�xDap�-{$k��J+?jq��-��Yi�Ν�mŝ �w�k*���N�T���J,2��܆���}�/���j��Tb�����O�)��.��7[�o��ѧ*��i4�� n�u���S u�XM�nqrn��=���	[V��m��GF��O2;��9S����=BXQ>g(YY�'�6����Qx	��=��sSz�%����Ł�v��((�>�g�E)`��/�Q{�&a�N�� ���	x2\�II�6���4@S�ω0�rG8�y��)W9�3H�_➳C|�����F�ŪE���!5�j+po'Q7K���`��#\E{��U��}/_]<���-�����ٱò�`���p�,<<�2~�i78��)^��zvx�|��&6����7��b���-�(���z��� ��V�i���{�T��a��.��D�8�V��x	bS���ʱ	_�+L�Uu����p8���S,\���3�c�7h�q'
�� �z�t�U@�5����r	#��-��Tʳ
u1��1H���)JHd�4 �..,c��$��^�X_E(��f$���3
}9ds�W�؁P���"%Tv;o�)��
+�<q���c=�@�ߙ�Y��7�]<4	�w�U_����$C����������fv���$������V�e���d��=�S
��W�+$v/��T����M_���
�pi�*�B'����#]�A���|zo�,8C�|T���t���߱b���L9�9/Y�)����|1���l��F�<��;<g'QZR�~��ԫ�Xo��Tjt��z�J{a��
�$���?#]�>/���7O���D��z�43v��7մ����{�GƸS|R<+9(�m��b^�`3�3n�ΒB�M<9 ��
��㰡�V/�z�-݃���4�|�9��J�M+W�G�^=���R�� F�
����g����!z@�#������������zAF<���!֕is0z"��(��κI@҇U�v�YM"�C���Kz &os؊��������{/�,��2����K���M0��`��ߙ�1<ka��г���gcL�,f��ɢ1 ��)^�r4��*�;L	o%bޖ?!@��Ĕ��q�#�;� �D��&ʺ�W�w��H=�����Z���)?cd>��f�Z-�6�En6�N����V��h�[� �ݫIC"I/����c�,�4`��vH�Y�-BIt.�@�7�V�6�K�-�>����
:i���c>����jR�R��m7[�۾T��4=����+�MV& �����GÝc�T�޶]#���, �]���1~oꭳ�M>�C�OK�~jG*P�>B�$���G�/[
)���k����������Av��CX3�V�'��Ӭ� �Iw����߉�����&�w ��?#
 �HY����9������2�E�HP�gL�􊟭�v����!��B�/P�J��(��;7?8�Z�-��aNj��ȃ4�H��R3 �����s!E�g�����+P�z�J����^��UD���� �@}��4N���:h���yr%�-�Ii�c��U�.;��yJl�[w�$H�Ѓd�!��k�B��ڡ���1���� fhc�]��C��a(mNb�<ۋޤc�p3�)��b|<���?�965��F�d�[N����C7 �Qu��O ���l�������kzV�}n��ﰅ*��cb�kKȭ�C�"�|(^���G�x���;?+������s�����*����sf�%2,'c�#��P���I�G��E��v��6�Z�|,����7���%�+Y"I0.x���(#���)3�0�6�!j�>ט+�d����@{����Z���Dْ��{g&jCȡ���r����Pδ�������qk)�D*���f������,�e���~�;~��蘩�?p|B����Gm���~ـ��ı��r�'׏���"Mk���T�F��H��h��@�P1��˩�2
��-�G7i�]��7�K�`��#-r�u��e.�fk�	��UC�n,�x��p�D氺���bgp[��4��D�:��4���`MQ��<�%�ڂ��*`�kt#���3��I��)ۦ8�n��S�����?!~�B��]���Ͱ�Q����O}���1��E��ʝ؝��Į�d�b%�u�_Y�t�Ԉk�u�G$��=��
C� �t����
6��%����!��+��xJ��>���=��7��IM���<�p\|�g��p��4?}[|�n"�]8E�6���ݕz�1����_����CB���	�KRy`Lv������|N����%�4tA��ۑ>��K"@O���m�p-D^ew�p�o�Q1l
�&Ǜ�p�����&��E���|ִ�L�j�m9	��Z�'V�U!IQ�H�oZ�w,||/V4�罀K�W�(pG!&�	�����|�ng�i<�Y��<����m��wy.��� i��B��;a_���y���w^V�	�����.N�T���3A��L�Sz~�nԃ#:k�l0b��V�T.1wbܸ
��9��;A�z<�m8��79͍�%���%�����
V�����f��W���!Y#��������k���l���`/� U�53L����nʥfî&�t
�;;b���,9�QzW�ЏZw���f����s3�*�[��;g^5O����Y3�ʭB��W+�#(ބ�ݮ5�e'�3�]o#��ddL'+/���f�����GHY����4�o�8���(#L�ĩ�_c�@� �8����r��!5�Uu�ރ�n�	|��R�M�� ^���Ei�7H$��[<��ޱ���G�[Ahē�t�TOT���-�&[�X6�E����}q��1��7b��^�\^f87}(��!b.�+����م���~5��C䗥6�~x[�w=.G��ܓ�������� svMH܃�rx�`Gg h�4����<SZ<;|���3�^�W\�r[��o�b�ke`�'�('�@��������K��ʑG"Y��a��������d�qM+�p�h��'��&�i�EU��q��`�2���9 y%3j�ۑ���AF���=�0?}" q�(�8(�5E9h�?�ָgm����z�^�N��B9��)�.Ȣɧ����W.���kռ��!��H�[6�H.���Z��I�����D�c�$�'p��G�-%�͌��I�YK�w�����C��*0�̭�������8����3�op�D���|�GDi�n;3����I�Z�� F��JF~��hmI���L�*�n�ū��T}�@�{�P. -vJ0�>,W�j�%@Y0���䩮ĲXS%��`��Ki�f̊K�Ef���X��G��C����l�����#���^4p��z�v<�)ܓQ5TP��_pe����ND�/�f[��V)F�:I:�gQf@2k/��򄹈�j�%����dɏk
�`i&��M�h�p��ǔyP�첯�YREWT��m�Ƴ{�j��'�&�A+5�`�ɵy@>�}�����w �iX��.��vb��@�Z�=�6�ˑ����(���ҫ�m���2��������s�4a�p����Y8ERI�x� ߿ƲWÍ��;klu�iW;��p`��ӱ@F���2ֹ�ר^?Κ�bg5�U`�o|�i��2�� wm��t�N�śFDXf�]�ڍV��`A�f-`{�9=�Ye�]s&j?*Xm*@)$��Pe���>@�����¬=��P}w�V��ha�c;������W`��#�jb�~� ]�f�l�qui�W�H�H̸	�����Y#=A�Ŵ��2�M{RmWM�s�?�1P\�H�X�@R �)�bڙ;�B������f��P���֢
�`�zM4�bZ
�dN��W�'W-� �;���v���B�WbuN[b�z��`�%ʊ�=$�#��B��3ދvW�>��[��f!��J�Z��&I3�.�S�P��b����]�^�� V6�̹����b[�k�n5aO��ڈP~N|�e0�
,�̤�z��O\���4������jY{e7���xtd.%���H�sĪ�m���Wً¿f�Kˍ���{�i����dߔ":��Q����}crK7��vͩ�C8�c�4��7J�g�E��R4�W{��(�Mo��|W���L?�e㢣~��8�%�$�}/׸Ų}�\mV�
ԥGZ6+2t?O���7�{����60�D�a}G�*?�F�} �,�غ�6�����"GuB�좜sa*���Z�qG�Mb�������_��i<�3�|���ȹ�?^�;�a����(���Ye�ۑ�glj�[~	���\Z_ϥ�xd$pk*���?V^�����wE���S;�w}�ݿ��B�#�Dhћ��xq,�~3���8��s��b�\2�
��"*N}X�֑�����&[�u����@˙(Q�U���E�L]φ<M���.������sۇ��髄�U�Q��g-���Es�3�M�
z�'V��1�X��)��di�М��ߊ�?�t��S������S���]	r�Ŕ�����еb�*�p�"D����>L>E�g�Xhcg�\,� f�O-�CB��x�񳱛��C MK+����u��0j���/��p�2}�!xmq-8.�<���~��H�2[K��dTY5��emyU��6�a9����x|K���l��g6���!�g "��m�SM�$���0/�3�`3Xً�����+�d���<w=,���/ғ=�\������ª��x�~�",\����j�^�I���
������Ӌ;��[>%�.�C�����m����x/�@w���Fz0Eg߼/�
�2�J���አ/�3P��"黊��b�-��4i���X���
��cEtl@�a��N��x��G68���u"�{l��k�j�n�(h��KZ0�&��QgR�\�<�0Z��a���C7K:��\gz̍ Յ��W���k�{_x����eφ��O�(���=���S��"9�[�Ӳ�iez�^ �5�pin����,l���2�+�1����.�_z�t��g�5�a��g�OE�c쟚�E����_�*>ך:��n��.�C_}�/�ʴ����ep�	���@���bʂ��	H�a���-%�pF$!�BY'gT�w�c�#L�ѫ�⟐�DZ'�҆{[/�Y����K�R��@ �wcC���"\Ƿ�ӂd	��#��k�E^�iF��u�m�'߁�7Q/���Z�e��nz�(�g�wG�F6tO�C�o$~�LcT�u��6_�2�U2`�z:0D���4o��<%hV*�j��RX��d@p顲�eAbS@��F����5����2��ܓXC������ ��[Z<fK����AHRݺ���F��t�c�T�a���1���2��g�|N~�4�Jt���.�+Hh�
AA����X��(|Q@���~�=�3�W�C�=1�.0��77:�c��K��8
=|�ة��;��}�23��@�\E�0�]d�*y|L���}ir�bU�n�B�84�_�e2�̒^pY������MߡYAR�5{?i<�$�S0���DM����_.h���1=�og��m�M�7���zM����Q!I��1�^Y�˴�!�i����p���vxW�1�\�Y|��3�+;[���Z�	V�LK �_��;�I���8/eH��Kf�ҍrq���0�%I�⼉���t�l��	����E�3��M���$�`�<�gf:�_(�H��dI1FEv�sS����<!����哐0���w�6������(��^>�c�-a.��i�n �hw����m9���}�ʹx�1<B��'j�J�__w5s����)�o<�*�ܚjڑ̮�?0�������`������+��?�{d}�����bpq
�!j$��-_m'>�]!�g�k�R����T�bc�%�2��.ge�����LG�.ȏ�au�1]�OU�YN�N�%�"�6�o�(�F�jz�0�����ʅ�û�W,p��/�Xrh���){�aD����1Ndٙ{H0�4�/��]�@B��)P������sb5d�U���"��P�� �U.B^j����������ʰ�׍��&�p�j��!ٍ�L���7V��_E�&�J��c�_p�6����<�1�X5�l	�1�xm�(T��N!(.����?wgf.�g����� �����:��=l�d,LSz�:MX\�Y�U���5��E���`.#Ѷ�0	,���>τ�p��#l�>cKB!�o���E�3ޏ9��͓���W���P)�(wЗ�Lմ��Y�Su���g�<1;��䆇Ŷ�ćQ�@�i����@^߉*��@',"C�֤�#(d���(�ŧ���9w,�����ICL��G�*{�#��tp�"�O�,<�B��~��5�u���=8va��ҫ4�O-儒{��/��2F
�b��>�;�9
I62�Y`6q�
%h!�ێ���֬�6C�SQR�k��Jm��A��s�{OʜIz�g��[�x`��P�ܺ-�a?98FL�N��$=]�ϝ�Ն@Jq�gʏ�@
��'l�U��R����t�ʟ<�.�B�=�h���2�Ӷ,�9ߵ #�e���~�XB8����ђ�q�5a��&V>e�s�?�U�@h�r��,J`P�<��焺��[�����|t
%���r>�ʙ`���Kx9̫��Q-1�L8#���X,�����I��C�v�S�@$g�^�X����w��l��_��Or-gv����p������ Pw��Bo�	���[q�����P������i��Ә^x:b�O�ͱU�T8W�y,�%��;�
��H�
.���/���;#d�&���8E�g��� ��5�ط�S�ʓ���|�=&�/�����#PږC�����8M)~��������c ��+�(ZVC"���9~����_�]j�Δxj�1�u� �_�D��W��VP티7�y�,�(�7/.AӫF�hu9W׼;�̷���-�=W�"x¯�ȇ�ޥ�hG�$��f��ҫxp��O!F{;5'UJU��B>D����L�'��Ǧ��
��
JfC�<��s�}qXC�� pE���%����z��둰g�r �Q��c�%,y���������7�u2����L�޹&�AsTH�?�Y�Q�i���ck`���A%:�]�-=�L����l�jt�>[\"N��PQ<1�,d�>�� ��⍛����o_*N��_!��n��!>�yE݇��b�:s��"�@C�
~vgՕ;�a�EZXlY��| ] &��������Y�&�ǁ#�=y� C����@Q�=�v�*�S�S\(�>:�K��F�m�o��M�IQ�;[-ϡ�o��i���^�3���@B�\NjD�o�h�k,b	�T}w�b�մ˄;�yU�7\�+�t�sx�Ɣ۟(�4b�e���Zޮ�g���b�zΤ���Ĉ�J�Z����
dh_175�=![���m=]�������2��;Fw�^l��e$��B��b�� ��:!���2�"����m�f�ssv"��:�W�����;�l=�U�V݂��AF�#�aDY��.ߛd�q���2T��h�ۀ*��ƁCo�}}���)���C�:�Pm�4(���czqC$�w��gʪ�U#�r*��=����|�ScP �E�h�Wu�$����G���}�Bb�l�^����vጚ�TkZB��e"�Op|��um��?�UY�'�|U��7��pec�aX
�a��6�͎S��h�ˈ�T��e�y�h8U��^ɉs)�R��C?�9�?rJ���@|��X ��\|��f�)5Vkp��ix`�E�J�u�ޮ�]�A�C����n�!Дy�[�k���v���/�p4�mr�j&W�C��4�"��^I�ſ`K{�
\���]m��>��om[��w�����`�z�.�#P���U&��B&��<u��o��C�,ԣ����×�ו	%��@�`�(�fv`W�XaG a���o���J
����3�vI��3@ �.i�7�T���3��h��[��г'N-�:�� o*��h�B�����h�_�N�]��kh�^5[��"�>|IO���t���)]J,��k���w�M3�͉mn�486%d�>���4.�
���j�
B;�LO^�s�
X���N����tIHMN�}�{�#�����u�/_^���T��%fE��̻���d<U���oJ��' u_�ހ��Vѓ��kmW��u�(V2��I, alp)7��50�r�'j�j��π�,/Ӈ-[N2�s���,��)V���-2������O�TI�~��O���O��?��򭃱�)�=	z["�%���]���~��Z�7+Jx�y`�J���W�&�����˸Zqm+m�f�^9�a���ˠC����Y��x�1�\t\(<D�[�eߴ�B��Q�C)�?�����G�Ў�q�����|�Y$���ԩf�4�"��D��i�&QN��pV�c�q�c���:ns~��7�D�d�� �+5��\�&�N� ��%v�ӞY��^�br���Bv=��%��1*��	��ĳ�`�m[���k��k�����&=k�LmPC��ǝYk��R
�1��d�s|�z�~?Al�6�1�슐��#�L09Ir]9v׵�:�$�7�2G���}�0��/��'M;I��/ð8 /l��͏��',�^���$FYM/>Sj�@5P�����6��M�D7>���Y����C'q�(5���&��ʾp�t6�l�5`\F�)�p��������xJ�0pCt;,(�A_!��
T��?Z뫖�'n�u��.����[-�az�i#�@H��6�2���!h��:y�����qU�� fړ��+^���L�D�/�Da?Y[�x��R9�vߓ�p(�Պ��	fn�,���ˈh������eMD9~�����ȫ|!���V�pRI����8^.��Lj�=,"����fx���8Y*����r�)1��ly�Q�5�2������!&����TY��Rބ]OV��];���b��P��ʛx0�d<�Ib��,��-bd_d��%��Xs7�~o�j�6�]����fXps
dHҋ���ƹg�,s�jtd�&Ǧ�a�0ۍ�i�}�|G��bI�M|y��݃�i�"6�aw6Ab�f$Q�pӑD����)�N�+M�T{Ω$ �|ڽ��^8��uj��g��\-qL-6k�M�69<U�!O~昌�QX͢�
-�yLZ�8o���.Ɛ�(n.�By%3`��o��F��x���g�"����+���[�ҪU�H������B�4��*����,�����o[m|hŽ�H���S;����\~�C
l�pP�ր`�Pl�V/�5Y�|I ]V������Ι��h��1΍�S+>b{H{��_�V�9Ls�����
љU�� M���, ���m��f�B:��U9f��hO���K@���na�R7�7L�S8~�Q�1_$1Vٵm�o�8;����N��b˸\p[�<���/'�@��(V!="�ȑl'S3��Y��(�����IzxTt_��EO�)oݮq�a\1�F�M��#u��ujΐ��$C���>�J�~���u�%p4b� �]������"�v.�&�ވ�lM��G�H�ȌK�Q��υ�!7	p�^D�����nŁ��:4�H:5+�q�A6�.�������>�Eb'�l����n/A�s߇� �+p~��',��)--x��������.�N�y��?[��\�7JԕT��,Oz���r��'��^����'d�S�)�d�l�{�G,�Y+v�^����h]�Z*����o��s�����]42b�rn:U𭘶e�!�P���0}�Y�ҽ�@��ك�����?�ќ,�c�
PJ�!����fR�o�/0���\��M������Z����H��VU�v�][���<�%��[#6��<����o�u	�k�j`�o�&�!k�b
�HT��#ݬ��ôIA��+=��������_�ʚ�(�\TU� � ��&��S�c<�/��g6�G��g9r���>%��b^ʧ �(#��G��س.�H���"GQt�Q]kK��H���n�M�@Ł6䚸Bq�����X[vb��'�.� �d\�S��u� wRՉ��2�n��HN��0g�e�H���H>륽]g���n<��=���.����J�����h���"_u!�R�$��a����M��}-M��=�Τ���G�~�%^�b}4�M��o�sl�Z��2H��i‼J�+��ǥ6U�zYH�r����Y��$`����C���	%����NAd�Q��l���T�-�1��F���]��N������	NЂ.�G�G��Aǣ��+r�e**�;��&| ��@���ۊ�=�o�ȼO��t?+i3G%�STrdF���:����t]�0��S��ջ��b�����ڳ<�j�4�j�ef�+?���Td�=ܹ>�3.)�Ⱥ�Q��&�)�Kp���"Y-}�(��5�|*R�~�7~�:µ`�� ����� v�V>R�/�7p�7�0�0?
�v����}ޏ�ʌ�՜��s0�rY��}wO�������3+ ��>0	)j��sU���a�I���54�QL����-�M|Q�����~�O%B~�����4,PՔx{k���zw�p����v�'�]=�X��Ʋ$���(pA��ԌB���w!�ɴ�?�e"��~Z�Q>?�in����Q��j���
&����&"rP�n��|L���O]h����-�?aI8,)5S����9��#Ŀ�x�ru\�����������8��s�1WͩP�cs`?Wv��'B���y��gB��'�\�w.��6d������1/�n�[��ؑYbk5�cn��R�^M-��}D[�䂼 �ǿ��7MJ�����n��^�z���Ĥ����obosߝG.,�5�E�
"�R��~��|\�X@�OD����$b<�]	��R�<��n�j����Q"�5��K��62�A��Z�s:���C�f%�쯡@��z��!����_��E����W8��v%�v���
�v�0�qe.���OVT�W">�xo����x�Ue��tIV�\9�Bگ5ܭc�c`}�6Mɾe�����v９�bLX֘x����WмY\���)�<�L����
g��D=����!�a����$�♘���ƚ%�>y�aw�p�#ۛ�����Զ��u!�T�)��P�A���{@> �(�*A٘���g,���Ixl~<V@��.)�[�>�5QI�{@������`�'�%�j-` So���X�h�`�P�z�0�=�B����D�p�]R�]����?>�`�ɽ��Qy��L«�W	��.Pg+�A��N�OF��8͸c�r��+ä;���F��r��ߏ��j^蹉�%�.�5���dW�++�0��l�A���ym~�
F1+*�?��/sm,��(��������i��uǪ<C+�C�6U��x/^��C�51����\@9�~��9�����>,I�vz,$-sV�\(grI��ͼ���RɁ�2#S������;���N�2��ﺮ�C�E��
�(=s�uո�D�*�=��\:,�u��tx֓w����RV���<��T\�* `>^A}�lZ)�����Y�4V]\��iM��y��r*����"���,�{$�[���|��� Ea����a~�6�D_Ȧ���L.���A�GH1E*�V���/�mt��-q�:�K�}d8�lh�����%'q"ޣ!��NB�D-� ���^�Ҷ���RJ�x��~?���x���I�ߛX��C�?d!���os�S�9Z��ro�c��	7������J��&�f7!{'>���m�1����_�����cM�A�5� �D8ER,����a���uR K�3���4�tv�%:��v!7�5��B�2>���	^5�3����ݹc�k��zM�
�D���� 'U��g���1?��&q�c�h�ч]������\ó�V�y|=i�*�٭[��w$�줱Ʋ&Ϋ��@}Dsp�ߛ��C��z�k������0߀E�>�6*��_W�䑋����s�=ҝjO��B�I���'�?�f���ȉ��ˁv���Ȋ2s��PE�NG ����\k��8,r�����%0I$�\l�ܶ����0.���&7��>Z��Ai=����S��ȓN[
�y���݊ZH��ؚߥ4��}�gc<ހ���A��qsTX%�Z�r�O�yտ�t����Qw��A�H
<-��&jai`�eّ�V��UM��f��2A����c:R�X=d���̕㶆	޾<�l�;V���K"�u����x\;���C�2�c}�u�����K�0��8�z�k_-�d�]�R��}�4L���1����h�b�Pt�7��������%�B�՘-!\_0V5,C7�7�.H?��Q1#g��3�{N���gJٱIv]!jn�!��ͳ��a��O�����<wG�h�R�H|�Mf��o2�͂%�F��-�iQ����ʃ�a��u���
�{7�f�B��R]�8�I�*w�>�[Vt�,�iT��&�2&E�v��oM�3�7��m?'1A����ozVQ֦M�h�'��?�ZN�=�α�����6#�J�z�y�Pd��\����#3�-T���÷i�t|������]�D3O����gX���@�IUh��e;��z����W�q��%�1Ee�e~��u�o7ڟk�zM�e�;�`�W�f��C]z�[�qիO�$�9�M��9����֚����@�䒍���;6Q����i�7�߃䀟�=y ���X|��g�:z�b��ݿ�(��..Mf<X�J��Ǣ��������x�c+-37�}�;{:2+M
a@�_|[Ad$��_5Oa�)������G��|��2�b��+$ y�6c����5������w�q�Zј��:�������E���ָ�x֤�B!�{7qJ�����CX�A�pe�y)E'l���
o�Mܽ7<�����2����`�o����Q۴$EÐ��&�8����>9r', f����+�b'N��xOY`�9���\�����U4���k}��lvk�\og��1�~���3���RPI��VZ�Vs�È��-t�v�)&��H�[Y�6�2���Xv_�����v�jd���:@M�z���	���M$W#��L\k��\���L������W��?�
�f~�6e\;c�^��Lt��܀b��?e�F��/�U�bF=�;I���ɸFE����Qx*�G]z����N��U:q�b���p�{�а�ܩH�Y���F�{��(��`�{x7�8��8Z�ˠ�:�-�������q����"��YRՔH3�aAR��C�iw�,�;,k����X(l-�5�����R����&V2��%�=�ɩ���� �3tYn�g"��GI�TU�h�8����\��4g`vQ�_�$���j��Ļ�lg�πXh=T5���U�!�j��VJp&�f~\z�	_\�Y�|X��\����-���w�}XKzEQ@sK��o[v�e!
gFJkτf� m�{���5��_$q��:H+ih�-v�@�~@�2)�j/��C1 Z�MF	�)����	+"��Kk_�){�.�_�T�CW�;6
]YR]!���M#�\]��&nB=g�9׽伖�Q�S.�1��Дx�w"+#x��!�oe��Ow`ߖ5`��4����>�g�a7<%T��}��'"G{謗��g0��e�*8�o��Դ�I�Y�[2j��<�%c�]̐��&� Aݡѓ\#'8�O~�J���߂��}�D�u�ᨀ�l���֒��e�zF��,2E�yzF\��Vֹ�T�(ae
� {*�;4��(ᤣ��*LE�>Ͼ��.��4�)���A�+A�Or�D�쐗����/#�7^��ϜQ�@�/�Ş�� Yp�r�xB�F�|V�2=�]��H�_.= N�d�l��c��b��Ҙm��D��ق��番<a=�v�����e:*ǘr���<t6^�����g��/�6�� Ʊ������Ɇ�}��Z��ŵ`u`����C7^�OӉ�~a�i_�1��U^T���3�B]�G���B-���a�Α�q�'�)|J�����~߻��Tz��b��ǡ^���E�����9[�2v�s���%�����
V������H�.jv�L�C�Z#�a���ha���l	�k�1D� ��?��w�T���	��UZ?�����(�yP puVW ���t���|�L����4�x�yà�p�ރ��B0x��6wFkew�b�ѷ���ϰ�.~S||M��r׵W�햆V�)9QXs��U����*FH�HT�
ec<g!`'�s���1�m<(ZN��uD�MCI��m��ϫ�������9pd����'��P���E��K�r-b�����<K;�G�٭� ����u��J�:@>����~c��]��G���j�-�W�&!�Ӥ�8����3Ez"s��v|��3����}#����y&\��ejͭ���n���ɒ�@B�Dl�hC�:�}��z9@�y�U�v��ƪ%��\����zf�׈M�;j?��2@�ټ�:���7����	����,�.b���El��������1�%���Dd4>Q	9"�����D��Q�2����0��e�<%��x���3�����>�{;���N�~1̷��h�tƽ |�;��&���]ql�	���:@�q�]����'傳���j8YaU� �ɇ6��
G~X�{���=��T˧!�QZ�ݢ쇪f=�yռ�YE�]`^�]�=M�.�Ae	=�.A�4�t��'�á<P����ڒf��A�P��ia3g<�y��Ψ�E~�T�3y?�I]�&"��D?�7�i�CNoa��[ѽ��H��� �D��A@>1�v�=Sٛ�!�]��v,� =c��m�%����]���V�:��Ǝ�젒�߫�����X����,5T��?�)��؀��Xo��@�]!�x�&5g�*�~�'�3��+y��UB'�\�xk����I�w���;L�$��QPl ��ۻe%�>���4i�)���8E�]|�E��\�&�i	����̣)� ����u�a�N51	�aS�G������P�"i�%W"��{��ı�]A-�y���Y!�=���%?{�v�mj�{AH^}l����b�� �̃7?��'�u��_߅=�8�(VfI�H+���,}�@"Ka|���2�JDp�K����Q}eVe7S�I��j���2s���\�������ubxK9�D�M<H��|ҵT�fe�u�n�.i��h�J�����E��������8�b:�{d��>�m ^T�V9A'm���ު?KƩxb�@�l�*C�4�S�xVv-��o��2���3�/jT�e�w~�<��ݑ)s����&7N+fx�8f;ƞ�Pv���o{w������x B%�P���ݐs0-[�t�Ћ���<� �V�w�F'(*��P��ԩ�=�X��܏̿�����φ�H���3}�2~n���!{�@��J�)*�p��}��Ѻ�w0�}���̈́��հ��I�f<�)�}P)�#����6�r,y��̖����W|Y��+�E+�b
�XSݘ��:4�:-BF}�
 ZA1;WT��l! ���r(H�7�J1�J��f�NT�5�I��%W�|���vRK&e3�PE���st�iJz� �s�g� L��II�I�TSM#/��l��_i�~��*����!��Rm��'*�����PL��ӻg~�r�+�?T}��Z ��~�x�"t�c�#Z�	';IcAi�Ȥ[�����c`7�����/3�����s��ګ��"9��9E+��"����m�����ǧ^%u���%!�k�,�oQ� ,���Xn�2D�*�S<#��:�E3� \h�m&����s�@�p�!R"s�1ˣ	^-�'0�ز�t�{����c����H��q��a������~B�K�Y��^WV�S�Evʥ5vǓ!���=���Iq����|�������1J�F� B$/=ι�!�Yl�OEt�=`�s2�~���@�,�e���2�7��p��h�x���9z0���j��]��y������B�=�yp2�#�T�.gNB���#k8O�ˬ|ʵ�L�mNJ�����seeW
[�ωnì���"�H8�%vtyrS�L��|�֡���>:��U������A㘝ǥ'<9��R�>ڗ������c?v����oW�NeE�E5��gӛ��B��y �����'5��s�P�I)VT�*9����9}u��0�����w���n3,��#cx�g�L�IǢz�>J^�,�D���w����������_�=� {�H���҉�H��}���3����@杺�]5�%����=�d���$W�k���"HU�ML&*.�G�q1e���w�ɝ�z\�vj[�:�= ��;�L������ �%��g臯.��.�����VW�L �Y��l0�+Qt�;���iJ��`S�O��W�;O��B�)�;4��1pL{cH6�j��w2��=B(��D� ��&B'G��5B��?�-%q1F�O��\u-��V���j�bxtST�Ԋs/)�O2�N�'��M��2;3�TD�_��,�ѐ6��pM���u\�ĺZ�0���V��¦,:���j�	���?՞:�e%a������r%��*V�wܫ���?t;z�P� ���z:[��x5��$��f��'�:�awi���upt{���e�$���X����yP����_�R�pa���-���$(�&m4��OP���� �k��?i��^<��<1=o^�`@����\�5��өW��$�kGD�'F}?��E{��Y�y�����+;��m�'$���*��M��$��2O���V\V�F�n��G�/�ʧIi0���L!t�Q�,��K�qm�b�����w�۟م͑����zd�%5�+�P�$������]�[�JBN6��|�)����jG��;�����E8�".�Zph�K,#�/e��A��c��f��S����[k�9e�u��F�b lZ��?�:��B�0�����0J"&B��}�s�s�%8i ��p�wz�\���e�8ŗ����n���o�q���:�E�s�Q`�qׂ��iD��x����7S,�9d�� �(L�Sn�`ջ�:We��oP��ٺpf��zD4���PX
��Z�������R��	HE6O�EM� d"@Q�@J�;�� �&�MW����uK��7�$���5�����Ŷ��݄	|{��Y��A��:
��J�O= �Շr����/������7�:d�fMd��}3GR��������)�^�Y��灬~��s ��ݯ�ܡ�H8f���W/֬%��
lA ����T
��L�
�ˀzD�ؼ�E��~io�����,'�1���:�m���c�ʗ^
:S�u�S�	R�j(�Nk�AL�����z$�A��A�)
��nHmY||��{�b��{��x���oC��q�_��î't�谾�q�i���?���,?��_Մ�^F�^��V�
����&������D�b��e�lQ��F��~��J�!sO����j���=�B$Q�bVOjhJ�>��iF��˦h�Q#�����j 5��FIs&�c# ���C�Vf�z+��\�a2���"�|0�of2m����MF����KY[���U�S�6T�C;�����e�!�S��#�Z/�=m��9�p��
���5æ��&��؇����� �����8�*�s��,�L��L�p$"�+m���/��X9�B��!:c��9O�.J���~Y��Y4#Aҙ�ߡ*gѰrӊ�_d�>��������l�����ٰ��q�3=�2Yu=�*����tӲJ��[t�,��o��Ә��p[�f}�C\�=������d�Ddz�tj���KS�v7�*x�����!�_�����n"z����DC�k�ft����;�m�V�]Z5?�N(�N��ii�~��?���@M%5�C.���ߎ�_{/�Y��HB�����딟-��l�Q�ڶ091�b"�7ܓCk��H%X�#z�.)�Z��7gxΓO�2��� ��߾�����LS����E���7'W�f|�Ē�m��[���T���w�Y��pɺJ´
��w��`��N9v��ԓ�#��j�r�����:ώ���}����
��s�@����$jI�����0X/�fȸ��Ǽ	�ހ��*�.��LM��?�B���(���:V�8���3�'ldO���y6	g�����"!�5I��NqF�_���q��S�cd^_�&.��m��Յ׋�3�,�E1�-ڿhlO�>A�R@�4�YdB���21_^�Q1JڴQh*�`'G��7ϔLd_'��d+4�à��L�#�J�1#ݙ�*����`t�<��/�V���V�f"�x�82���̙�A�����	˴����"ɇRZ<�iAĻ�\�g�ұb��ŗ`z��� �v��>3�6�
N�7+'�����r�i��KH��BrAk����G�|f�[[h�K^�խ~Hl#��G��e��8%��'��Ka����������{��"���s%01�Дg�"9-:�D�ʖ#t~+��'���yk����*$� �l��E����p�`�
���m�5kV��R���V	\��}��u∘^�o�o�W[��?qQt0 j��� d��C�4�ˁɋ�7��g�d��?>���b�䕋�n�7���$V���Sj��w�>�z��~��s�a��a�:�N��w�.slC�,�$Ou)�J��\�X�МJҕ���,���q��8��c��/5͗�c�6:�Mc&Hd�)�MA���:Ν�l�LH��$t,+�^����t���]�;
�nh��6�a�m5���uN�\1��FL�?�Sv����O�V�8����@��U754���w6�F�}��<-��-BQf�ǮYd�N1��%�g��!x��y�#v]���yVάʹ�gB>��� ���Z�NӐ���I��g�Y{ɵt��u��?8�����r57�����u�	A}��%fn�ս_�Ǫ���D����]��nG��<����:)��l�ȏ��6��A���å�*�Pa�G6�S����a+�B4r��xPe�t��WV`��N���ؔ�Ę�80�޺t�>g;H:���܈e�'K��@�40�@�W5��"4�6�`���A�m�oi�Wl�A�]%n�1��@��ܨ��;���l��hQD��Op����?%: �0i�fY��
Y|�W�;��ϑ��}z��]��wB�y�zы�[L��6㿷�OzG�.�k(����R?�lb�0�4��EHk$}�&�Ypn�����ԡ�Kq�AXY�y��+7������a�nX��$8��0�z
�ļ�����dsZ?��6@���.*Vs���O�r�<|h��d�� {��<�6�BG�H(.�i���8)�����e��ɷ1sF�'��-})�v�Hg��G~x�i��?#�I��Ip�ڰ7�C��hW[k�6�1Qċ��p�ȣM3��s���`��_�JX54,�Ýp� ��R�BX�f!w�ˁ��7f�t��H4�b1�-s�Ӂ��҉�_���-7h*"�2͡s�~*��?^+�[�J��@$f>��k��.������p�e��1Ȑ���S���H$:�4�i����|�l{���s(��%�T��=W̒?'rtD!O�ۢb,ʉ�&�j�ʨ�������d>�#&`��Ilm�l69��y@W����v)�2P�n{��%�]s/�LG$�����ZP6��4�y�|^ǆ�}64٪=ظG��}l�/l�,�B�]G
\��k,|wř!i\��o��I]��g�^�T\/����-Vַ����d���u�;K������ԍg�s���27���@��%��^��C�5oHw�z#����Y��	�3 "o���҉���G˚qi1s�Ǚ�R> A<��+]�-���~�=�7���*��TO�J����R=i>�[EFl� �Z�8���t$���y��o�|^i�Ab�@��bnZ���d�$�r��N����Z�R.|�}����'�t6�|i��>�~�S����j�3�����"6O[�H���]�D݄��2y �e�#��ٮ��*]��U�'!Í.֙A�Ov��TB����.����̺�b)���PW�H���`�����3�5��X��I�l������55�ځ�+ԟ�zÞץ�����DL���L=[u~�=���7���S���,iW) GMu��m�֌�Џ�)r��H���Q@����᷀<���"���7�Z�ԁCʂ�U�r�S����ǻ�;��6-/)7΂1R�W���h�*/G����W�{�䫓���nvE��H�ƫm����R�Q��b�bZ[�aT��c��5�5�xi����P,V���<GG��t�z���D&�O�!QA�u���	�m�B�� �k;W����!y���(�m$kN� '���m�� ��H�
�����`!Fd]���7 #����9r��{j�qN�|}+�����yl�/a�T���?`V��X�5����d�T��5ȡ%�����F�p!!5�A�:�	��V������q��l�S��8:�Pe�]K<s�*�e��6p�+(���Ă��O�41�����ZC��[!1��ch�b��V��Ð����(��CaPJ��)�Z+?��R	�1Kj$�d,����>:�i
'���(V���9L����4=���B�ਦU��g�)��������AC�]�W> ���D�&�v�I����m0DW��@�����K��Ʃ��'��@ܨޣ����"�A@����CX����M����G��o�Z�/wˮn�?Od�5�ì�q�
��U���⍬@�"�
^�P]� ܶ��Nb�_ȞL�;9�,��h���t?���]�y���z����^T�x��F���0�s?T� f��& �\)����/��cG>� ���#:�
\�c�t{¯�H?:�~�����g�x4��6/�{��9�48�+;`��e>�����%/i��4�ǋ��� 7p�GC�Ȫb ��L�����1O���o�K%$�^������L�	2b-̳ƇQ���6���5N/���3r��!1�=jE�`�f�Y��'��s~��ރ�sF�W��(�^~$h��HIHaofz��=��]���ħ����]Ջ�9��F�ޒ��\��<��/}��0	\�u&��4,�4���I]�^\k���YQc��9;=�G/� ,�9����\�mHzI,���^7�r{�Ҧ�㚶��)7���C� h�|����,a}u�Ga�]]������n�r�o�tg�ikT��V�|��Eь�D��Uc���֨6F2���@�Q�A'ɰB���j��n���X����-�K���n7���1���_"�(��(o�����!�nq�2��pG�ϳ�J�l`]�c�����߀�<�"���V�γ���K����H��L\��"�����@g���۹@/��&�,�	��vk�Sy9��xZS{'���u�i��"F���9�Ϛp��ۆ���]Òy�Aj���6jE� ��� hm�K�(p�U�>Is1�7NV�l8��ɊYv�L34��0�d���G�(�\=�
er�
����b����dX�,����}���w�2v5M�7�k�?��&����p:70!OAi~xl�1z�X4��q�]�Ƴj���6	�=��pv��K�g�Ρ��Km�Yl���`E�GR�����_t�՗���Z����Q�mғ'V��%�u�r��Yћ(�!9�{�/V�����u1]��4�Bߞ+:g\Av�Ç{0;[y�/�z�d@����D^�v� �R9�Q�~D��l*hR�fw�px�{ɂ<�N�8,����2��ZÒ�ߤw��_$�w�
Sμ@�J~n�h���	?��K�a�&��XϿ�	�	ټA�;-�uA42��p���γ�Z/̛$+��k��Bl��usd\	��Zf'5g-�#������#�Y)v&��ӣ�B�[�M��XP�/w��(�&���zI5u�����WaN�>��k)x��t#~_�:/��~��͇�t�CO�*����@��3\pۜ�d��,,����O�P�w����
�I��3U�zl}O�bH��Ϯ2	.;���*2�B���S50����w�/�x�X���|0x}�E�*t�0�Me�:kH���G"擃d��QEvl�iF0�& ~�sdV)c�a��g���Ua���uG8�	3�z��bq( ����YZ���S�r{�$�!��yU����֏	�t1�p긧|�t����q�o�u�/��R{)���kl飣x�F1�Z$	���j�iQ֘��[u���l��M�]����^TJ<�@BW?�p�e,F�K�%H��z�P�s���:���&� w��N��+�����]']��E��)IƋ�\��~��$u�|S��z9�������e0�r������x|޺�p���QWUUoeS؂
�����m��5�n�u�����W�[2�S�0|{�����`-���S�=�2�$56ř�va��}UV�w)i�T#7��J��_ ���������ŲӸ�z���.��ys�a��F��.p����β��QS���f�2��rȰ�7��"�A0lc�teؠfT��y5�!*���.�˧'3g���B+�����P%�������~j��y������yW�C��iߎ=a����ڐ�s�F)�_�V�~x�M��?<L�FI�.�h�+ .h{-�����|��Q��2[���<�Og��dyd�qz�e)@0�N��Ll>���	�sx� o9[8t�5�������u�x�?{��V����!yK/W�E3�u�f�=]{�j�)���t����f�~R���})8+������An��C�����͔\�����^e@��s���rs+������a���
#Gz��[v��}Xo~[�*���m�����������(j�|h�i<~���3��B ��:
BD�I�	�Ȏh��p A��u��1�h��ᔉ��q�8���a�� cm��������'6�������?ؿ��-�	�.|�B���L�x�j�Q�u����S��>�@�����&�j+}�N�pS� �Ck�E�%_�&�#|�\�9b���o<v>E�@��ɕ�e�!�}��b t�������J<p�Th����!a�à)M�]�LN;ȫ��l��h���j�qQJ1(j;�2���˾&[*_�?��K�����ɽkD�;H�&���H��,[?�%on6�q3�HXx����. ��L��r�W)**�����K�����t���0E{��~zk�������g����
Gkhiʗ;���߃�BH_X�&l���)� _}w�6�.���ȱt�W�^�^���=����#�L=�[@���R�W'(�L�?⭁���^^��mv�k���ۈ&m�]�����w֐�y`�2�93�U��c�5�5&E^��L��H ��!m�:U�<�5 R6'��Pb����#������.���b;�궁6��TT}��H������p�ԷQp��"ڇ�Ʉt���,��D忸=/0I���:���T�T=BġM���J\
FU�I���k�<�,������1yَ�=<����m��Z�6Ⱥ��r*l�GI�k�9�D�I��������k>{��#U�6�:m�B�^��Z������y�2�S��[�7#Y<�k	_N�A���-�~>B�*v8��7k[G�O�������|n�r�>�o�/�Y�&A!�V�#��X)� ��k�5)}���i��0*)~N1��DvbE����d0]���u�~!����J��^I��L���tyѳp����"/O�9�P=�ʲ�)�cj�-Gp����w���&�M	��,�ἔ�q�	�|h�!%٧/Mb��D	�����=)l�Q.�~^z��g�M&�Uq�	E~�@�!z��td"��b6�ץ �C�cd3`�9��By������n�ӵ<)���X&7�������Sh�bX\�5�~ӣX�w�R�5J;������K���g��Y�f���ۢ�e%�
Z��EZ@ �@�9W �H���*g<>"�}��,
ߎȦFq�c�S'g�����<�}�p��Y���A���
Q�玉q���	q�Y��ֆ�
�����0�]U7����D���.�C�d�b�滘SK��Ba��"�G�t֝t�Hַ�r���L[�+L@����͔zp*K*�|�ѐ�"qN8��,
��Ŋ��>EZ���V�"Ƽ��v���8[Q�����cNAo���:�b���si��S������?��Hs��X� �ƚE�3����V��E>��?������zz�狖��oFr-��������ڀp���و�-s�o˚�3O�;��_�>V�W�m��V���ُ�Bp ��읤�ϋ�Z*�L���V��8���~��O-Z��I	�>R��M�2WQ�.YY2��҉�}%�8��t�3�8�c��X��A\�-+<CaAY����1#Q�{��
��B}q#.���JW��̞G]�O��ڗX���b�ԅ�u:8�S���ĵ�Vcŗ2~eR�$� ������
\�A^:����B�ݱ2�/�Ā5��LƐ�!Uk��@n�ZX�惠vU=I�����!t��/�����IR8s���>+�Qә:��I��^� #��p}Q�$�#�Mc����Q��|�ȲNK�3^�Wǌ�x��zϰ�u�I'͒��W�6�l�*��%i�|��LTO�h�\�W�N`X��l��c�B�T�/X9����||��Onl��Z;��3�������+�AJعP|2�b◝,�b�hm1����vӢ]�^�\���R��x�z�M����A<H���h�ω�+�`��A�d'-61�kڇ8��X}��8d)4���-�㒚�ѐ0���8�;��d0�cz�I{(�|6�<����!K00uE�'���NK�M�F�S���r:8��H�H���h��0�Ra��-�Kf�kԚ�uL�d�r�x�-�R�\K�k��;���(7��,Av� ���C��7{[�֍��)��@M� ��A+	�-�;�3�v#̥,�k����)��w��;��9�\��`~����J:y�\Pn����?�9~�)��f�(����QЧnnq5�AǍ0�������n0��B�%�,Ԩ�����E��x�3��Zm�\ ��^��mFo������(i/���
i�YKNj$�M�\%��4ҡ��#�޶�ש���s�bIN��Ms�ۮ�x:6fh���aᡙ��-G	W�m".��\5�����w�[��oe�*��YK*ZqF�y�Ju�	�Up�Lt_�r_!:���u�"��z�0V$��:h�U1E�\�c�D�]d-��	��.l<k��ڹ#1���뛠��9��/���~��Al����ή8��貺���A��M��7�/ے�s���,(�"���Z�׮4��T�P)wݵ�O�����7�"��[�ՔI�В�37H�C<p��n����CAȽ�٦.���H�6��u�)2��wg`�3�4��G�M��ϩQR����/_�/��¾k�nc[� rT�/X�%����#e��]����kT�V��6n,�F�V�7�>{���B5��cܳS\�8�O��w�1t�V~7c�ߕ�U`��H��uu�-�u{a ��=�E����M�Æ���:o�D��^�ʲ����H��­�����gsD�y�, ͋B1�3�"~Tadb�m9��-��&w�R0���uG�����0�JqԶ[	B�P�8n�r�K٨������]�'���>��ܭ����;J�E	�8��g*oeVB=%R�.y���4�XFn�_���L��x#p^y�7.�%I����_](��_�O����
5�R���!"�7�K��X�g��{�\��^D|�hX�j�-L�������U�t���M}}P��N�*A��Zis��x��7�7a���+�	ŖX��3�m�ʎ��X��?���nt+��ёH���hT�{��`K��о#�>�	c+�&P�zLTE���첕��|"��+q���Y�+���"�뷹!j��I�Z�#Pr��#dx��M��L�|��md c��e�rm��/X���+��Q�cp�%bǤH��X������pr�T��i�q�Q��H�9Ŀ�Jʏ.t�+��.�A���g��7��f+��7a>�.�È�{�� ?Ur=�WRM^���W���&�%)��ep1�M@"���&�R�i;�c0!����-�go���U]+��
t5���"/�s���K@�����1|�� �i��z�03ǠF�v����Q�|�����]XM����w���s>�E���'HPHh���ܛ���+
�
Y�>.��Q��]�iD�@�Q�t16�����	#;�*��2���;#,$2 �4������PO��
�<C�Sy������Hd�i,������� ���k�2��?޽�$ؒ�U,&$��Il��4�}�i��L�4��C���Wއ=�-�]|������OTA�>�~Ӽ4.�뉀S�=�T>Iv�3���2��ܡ�8�3�en3�A���f-���Ȫc6��*_�c+`D~���wL�y���ڏG��{q�e��ƫ�ۚh�W����c�b����"�q|�Hrk���f�L�;���4���,���$���(;�p����h��:�Gˈ!��0����S��J�����Lb� ܣ#�`��\�����S��]k���)���&g���}��D� v$�ϤN��0dv��ܠ�m��a���+�)$r�����a�`���s;�JG��n���W����(+(�;�ŧZ�M�L^A̝J�[?��H@.��(���˹>��݃��U������V^tmZ�(���̟����>6|
�I1*?��\n���ZɈm�n:\Kt��jh��#Y�(���ѱ�R�ƛ�����L!YU�.����v���s^��>a�N"G��n3Σ�A>��xhZ�D���U$RoM�#TG����@'��Y�:s�{T�<�O�������P<ӷ@<������u_�<��p�7�4��=��,R+m�����A�a����s�-�M-lw���@���ǽ��l�&\��Y��8�f�l [R�/���Rg�S�Vm�����fT���M� R��]��i� �Eb�!A��V>�����M�l	�p���͢;�<Wi��i�=�7-����k�v�?͵��V��1�
��M��׳����o�V�ȥhѨ�|)�;7��C�#�a��+Tp?'�<�lb���w�������%��Ř"�c����M�Y�(֔�l0�*�� P8b �Yv�{D��n�$m����*~3Xzu�F#9��E�ɳ ȗ8X�뮓²��eU  �����n�(h�>2�������""/v®�J��� Wl<�2��8|?��J��H�s��~~�C�S��^	T������yXm�!�ܵܲ���@�̑�Y���r�f4<)�����˜���Yx�@�G���i�Op2�� �.qi��p����"�]o[3�qV̗֚�(�>�i!Q���("�#ɇ?חv��r�Ŝ5����p2�G���6칣�x���}f&�W�n]��_(�_ �kB�)�M�-Z��#T���֗�/����w,ʾ��CpC����$X�gߤ�r�f(��?�ƻ��Q���8�(��4�M3,'�ӈ��p�|ܗ�(n��W��2e� �:�dc�B���5g�HƏ_Y�8
�X��Ҳ]�0�r�:�Wu����v=K[�q~a7'��+��{�/r�����ou�p�mΫ�,��n�p��^�u���j�:PaO���4�����<�d�0]���n�Pu�nM4a��xIĵ	�MAFcՐ7��CƔY(L/�ݽ�������k�*���Y= av'*���r*!�� �^�G:Q����89�^����D�1j��n-k�y�oUJ�e�|������ݗn�gHH�(����չ5�.�#L:���)O�bξ?�i�� "�,�P����ȇ>���!d�!]'�ZV9�i9�>kQ����T=�Eg��M��%TD]���[���y3�,��;�hE^���2x �	�p������)������:��m	Q>L0]��>�a�<#�XR b��yw�i�w�����c�0b�6O}�߮)��e�o�\���A!�'v���������^6���ٮ17qҠ��_}'�jD�Z�2cV�y7����64��I�,�T9U�������=�#��U��c�4�� ��:��2$E���* N��dI�� α�$�'�	1t���9Ĭuت���q&�S�4�vN\B{��Y�D�9�q�81tc��iKGem���t�v���hr�w��\>�W� 1�;��Qx��U�!�Jĵp9�ɂ����BIW��!��q�Z)�7����h5Ҕ)��n�=����[Dn�b���K��B��:|�к;��ω��,9�LXm�/��u��I��R�/6�ʛd��+Pb }w8��k�5.R�lS����.��W��sjM��*��bB�����b���xw�����k��ܙ��d�����3�]zL��a����쬈/���!*��l��9>�@���m{~���N��q���6�>X�M	����?7�|*�̟�Y	�`g�%�\
g?��Թ��8�^��zo��8S�		�iIw�rO�~xk,a����������{�G�����ł���#��H�5��2��K����NM�/�`�"�S�[̮۬]�������0Z�}�\O�Z%��>	h�Jj?M4��Msy9z��j�օ���gѰc�6x�#��W�ŮȾ��Ɣ��:�[:�@��縂���Ǎ��C�[�p�! ��!���p^IMM��lyR+o.�~�\i�ϪiX��y�����EѥU�ۼ29a���9����������bE��{��s`Vt���Ŭ�,��������C�-,�B.��r5�q�U�GN��z6�:��O��P��۸ٵ4�����OF������D�~���$3'�̰;Oi]dYh\��3_�j���C����2)���_��3��*�����#��K������N��(�s��� �w�!�i�E����p���E)p�͘�×���pt�-|��>�;����IrI1�t3𜹖�}+u����q����c��!���L-hSU�
����}�q~���g��h3�S�F�x!8`�đ"�%�5Eı�u5�����j؛%
��/1���t�Y2�88���=?ơ���6�7�1�tqN+UHYg�Ǝ�_b��'Rx|�7���AIc����Q��,�IƋ���-m`�įۥ.i]+Hp�rΩ��m�+~~�8�=2oJpu-�5J�e��?%��x��jW|�]��{���TOǍ�ݛ���v/�K������ �݅피:6�����k[yh9�#�

`?17H����ٌ�_�Jѫ���EI`���|��=��zU�Ի��1�\���Ɂi�/��\�
�h&�S�����f륄���z�°1�����a�o���ۑ�ִl�2��c�]*:��͟"#��U�>P�U\�<J���,�ӡ���K󍌧-VSk,%��HrA q�F��$��"�����ڏ�~����Wr0�iBzd<�(�vQc��N�k<��K�Z',��
�3�ӏ�`I�X�1o���n�'��O�� ��R|��r`���i)=��[30-	�i���7��C��ҟ���:�x˞��i-(�~���0�++���q�FO���G����8�����bEk�>��%��.=M߸6�C7��Y��^�daU/��Ye����
�+~�I�-V�J�����<�eF8k�	��1�`9OM��L�[��{=��~�������v�ǝ&����o�r*��T���mգ���:�;'m��U��x�8�E������2Z�J�.�����0�M1��wzw��䤫M�~`X�/Y�4&_��ޢ���4���$䌅���ŕ��g�������� 	Wh�S��^H�����#o�S���,�=P̈́�
k�̰'���~��ޡ��~f'rܗ��)�F�GԢ����*@
�k߇�h��;<
��%�(���Ǘ�� T��,L��w�btI�54rRB�E�y�ZY���H��[�t*$	#���_�?�T�����2�6��6��*Ip��w�.~�.�_�w�(�Ĉ����Yٵ�-Mp=KH���m?��-j;��f����73y��L��d��j��A�׋�j�,�c�i@��Ń/��6�H�lt2����Y+L������t�${�����e9)�n������yR� :��Sk������n8V+����M�w��,�{t���ڝ/��ѝ�����^7���ׁP�q�'a�X���@�/ZX�6@�M�	�|"�2�1�Z�X4Z�x�Lr^���Ш����U�O�QKo�&������'���K�Ds�|�w4L�LŃ�Eٗ�?�7�����r���9x^�� ��d���)r.z���۩��L�Z�~�`S���>w�L�"�Ԟ��z����l��e�z�m���	0J3��"O2å.Ix���a��[PҺu1�� k�ю�"�.��L���&���Ul]A��j/�Z�O���L�,����_�2�Y�}��B�[	��������6O���]B1��C�� ҂�ev{�����Α�"��N�4���s�km�Kj'Z�?\⌺y1�Mb���K15����GW���V4^m�R��y�O�a�ߞGin��A�%��p����_��У�}S��q��;���qy��>��<��/ϻS��X�[Mg��)g������@�vB��=��?sKϼ[����n6�J]���mۼ���"?fO��!YV~�Ib���ƀĝEKC�[xZ]u�FE&�lg2G����@}* t~&�;y�~��#&H�,��~�����
jBBj	P������Q��W�E P����4
Dq?��i��=�l���L䆲ǋ�
 ҽ���E�9�(	�R�E�4�����N"|�8����`���}uf����޺�7.����d�A�͘�R��eL�Ct����x�2�w���B��$`-���T!p��ϊ(��ъ1�iz�˚�4�cl�Y�`D���^��䲧Z&$�ݟ���}��!�\�N��ڝWT�m&6�^��R.�\b�0j�c��:��H�;_���@���9Fq7>с���e�Q8�)�/��=8q1�c��~H�:�a�-����3
��6J� f��{G^��x�&���O(T?A%K����`0�$X�9$|������e��ϭ�4zܵ�����6|n:	O���q�t���=�u� ��r���xj����7�%o-��������f E�E�v���k
�#1(�|�?�a�Y�;]�.�{�1Is��_ԮfZN���ũP�hy0��GZA�V�C�d�Ÿ�.��VO,4�3��-7_��-�f9�4	�W�%��y��҅���T��~n��<����O��i�:�*=�U�֠x&3��9�����t�j�� a����'�:褿42	���V��!r)���̗}���L��6L������~K�X�O�v�~����}^@
����+!�L�g�('��p��G��@w��ֱ�V��>>��m�L_��Xq����g���Ƣ����o�NU��,�+R�l��zh��"!V���)4�	���/Z�u���o����-��|ŷ�N[���	�5@�.Z��9��&3��ЎD
5�@k���0��Ͳ�=��kc���y�QJ��wD�1���8�i�_�h(�[��4h�%�t��(�|�;�(��ڸT٤͉��B!WC<���U!)��1���Vx��,`
=��28=�h{���ߧO���B<������@���}M:��G(�%2��48�p����s�%y6uu���?
����I)�Jx t?>K�jXR�l��8̳����}�0�e�wI}]*�	~7X��+N?��ך��TѰ�{����H���1�sZ>���ַ���P�+e�s�M�F�F�q�#���P��LB�w�E�<�hN�Ac�D(~��]^�V���AAu=���X}ZF�x�;Fv&�H�!`l�<c� ���u�&#+3�:#[k?��R������������s3��B��8��,,�
�m��z�"�����{Ū/�`�n(e�X���ن ���	?%����!K�m�%�䚯���~�ۧn��U�)$W�2\����#[we�`H:ڈ�Fc<�U)��K'ai���@q��k�I��2.'i�I#M-����|�X㾹k��1����K:\��n6^��hV�Qu%�g�J�.�RAE�!�ب���e��0�Tv��k��="+��&h�2Qt��;1���t'�f�x�}媭�6'�}(ͭ":�S�}L�B��-/=y�*@T֎3a̡�5d�:Rޥ+�-���/�6�����MsExהh��1
N;
QFn�(��@�K�{�e���~�Z2���`��V��I����0.�������JE�2����IT�V;�ց"b����V�>��6l>�Pmaױ�\W�N�H4���|�ֆ��4f��b�]�`Xg�W4���b\��Z�����*(�͕����wr�ws�	Yp�:9V�b��*��d�mya��L�j`2�A+��6��~yL�^���X�'�,���F��$�]YX��u,�@��`�v^'j!��װ�!�O�Pϱ�S��!折V*n�朹B�� ��Y�B��������-$@j��1*�q'W�=9� ��*m�Xi5��܄�g~���dv�����������-���͗'�y"BI�6��G�Qf�˪�J����P)�j��Y��P��\���U^}(E`�]t�W�2�Q���ga�l��*|����x��������zO���)H�Rf�4X"��R%.���h�K�?��Ώ��h��Uq�	�0�l�+���܉�K�r��DW}0�Ks��������ʰGr
������@�
���v���/!�`[L�9ө�����/m)�sm�ߧ�f��q���}����Gw-UX�j�X+�T
����Q���h��۵�A�"lZ"F݅�X\��qpj�J2煅Hm����*�3)��Fɖ�%$�"t�IajX��'D�~�l�nW�Ż��f���
������<���㓤��[�#Z��#��h.x^���T`'�p�ue�� ���|1K�L�(�&O�1D�.��N�P1�n� �V�| ��hcۙOu���:��sM�N/��HkJ�$�|�?{1��'+ ��� �5��<�9��j��K��H/iEE���q�)5��k�oh0�x�W͝4�(���Q�N0X�aж�Y��o�adj�^)#�;~��0���)�������Avx�9����=yE�!�@��?W<���`�/l�M���V�q鏞�@�(&��%ˌ��iBqYNk(H'����"�U߷�?ۣ���D��(hg�s�䏈z�cS�`:�G�H'*
��H+��#���Yˣ�"gc~�^EP,86-;���~B�wG9%���mģ�U�\<=:�����:��k����+�<�K`_�1����'�K-���ޕ�+�a��kIxZ�36N��ҷ��7sj^p�-���j���S�ר櫺lM��1p��B������* �3o�cLb�4|��v��l���0��+j9�
��mﴏ����7�G�'�o��B��_�bQ��S/ J��v-�$�Pأ���xd<j�����x����~��@����"D�������5�U�<�. �m�
ؤ�N\]M;0wL�_�0�07���c?]罌�	笅KLN��H8u����xT/�u�G���MK1�XS���Yе�I��V�������F1@�1�hj��B�<P��ڙ������5�����9��bŖ�B�)c�ٲ��#��*��e.d�O��B�B���/���6ح�q�K��_l�h�y'���z�W��>U��I�XF�ơ��A�ۊQf���u���(weKz�q,�\���);a�VW�{\��]���	E �}��s�X�]�>+pG����VL!��͊.��.����]B��XƝ�&ǛH�<Z�o�J�k;��?vq����*��J]�^r� �>(l������ݝYq%/8����yI�/K=���>��K�[+w Q�c��iڌ�e��F��Y�� ��E>n�f$�?��o)5a��=��|�!�?���>�gH�/����3�y��pmA�"����c`06�s*a�8�l�xh�ms�v2�lC���X����?t�,B�h��6ئ�qaZ�����U:��U�T�;����g�����4t�c�\s��ɍ����)ǅ��#̖�������l�Po����D�������@ԆA�B�]?���`-WH�t`%�qPk���e��٪; �Z�����#�Ӿ�k 4$9+[W!D�����m�f�+_��E>~GB�!��pf@�0��)Z=�,=Ƴ�h'i�8���7H���_��8�5MwS��J�&�w	cRH`����j~o��,��D���wKO�����w��(&:��K�v���R��a�uJ�%� s+�� �
-�����^J�O�6y�i�G/��ôn����!��⫚� �o�%��v_Ȃw�щ�>!�	8���)� ��4j1���2>fO;�p�KV������`��� ���T�IR:�b�}�\��쐤)�{�:��l�@��z���?�_���O���Y�s|j�����3�,�����U7(�׻X��|s<���D9)_���_�������o�Z��i�0�$��ҋ�/���,��ef�+'&�}�����#'M�}"�kQrW��uT��8,���F�X/�4�a�����s�{��'4��)lɛ;���Z` ��L�.��j'6�lA�PÀZ�3$�a���Q��#�d�~;1� _��[s#�f����O���_�T/�]�|����|Ru�5��4��r�vE��ݳN�{��?�<
� ��̾5�>�%Ia씊FM7)�&�HP�{䏿�Rśߏ6K�RM!��&�4Q�Tc���]U���)����-����N��	�@vU���m@踣D�>Z4�qۚF���'6����
�~x���Se|��v���7�t�`�u��Dd×����l	����O0N���p���e�V43�����)�����#��[0�tZ
�Ɓ����Y�5N�|9�e�D�e���:�P�a�n�������Ǝ.&���q6�۞�3���,\�ipNvJ~#�+��uiPK�x$M�wY���n�'��HDj}��X��*C�aW>X�(�ÀA�k+���I�L�m���=mj�N�g,onk�;\����������M�e�]��W��I�]��(X({��(1wf�E�赳V��{����'�zG�d/�:h�XT���ꈓ�����=K�'*���皋ǲ�&Iwl3Z_��Œ��:2M�.=qt����D�t���ħӏ�JQ
�g# 5���}��kKj<�@���ؑ�:�u29䕍lc�F�*�Χ�vvf+����N.!��ld���K�Y��W�~F�'���?,�8�3���G��<��%_�p�y���o�g�E�!��fX/+!���
d��Ι^���.��;��l�1����%Κ��0�;�P$��җƟ�{#�X�^��(���YT�n�f���7��q�u'TPe2Ŝ6�@����#�I ����?����Ց����Ll8Q�*�޷��v�A �N��ԜH� e��u�>n򻁠�;����o9_��'3�p�����i�Y�6  {��^̚����+XI�,0�G�;��A�g�xT����ˈ�o��}茯�`�bYh���>	#���u���+���8l���,���+�ђ���Z��� ��L�1�ǽ~Y��(��S��.��K��i&��RƁ��"���o���p�{��0= �T������K�+yyH�u���ז����-���1�~�j�<o�W�/��h�qs�#�k�f�)�7�^�7�5�t��+���;�ëF��:�~�U靃��y���ݥ��;rD�GƂt��>QNE+nEl�Š��� ��53(R�PmГ�n?!:ũ�GO��m������kkZ���6b��A>�F����@���0�(+����?���}�[^Z�^�?��+�1�b�{����o�E�ɤ�x勞pL�>�����|�5܏B���t��xÌ=F�!��bt�3���f39��5M�G���|5�\�y�]$����_xsb�}:�Ck�=�8��v6����D��U���|�:;��t�n��o(N:ˌ��[���Ԉ�T���Ո�����y��G(/$^��Tje������}�|��j/���44����ry������^�<�U�lΗ��'R��l�ׂ��Z�(�4��� a�Y�u�K���.4��]��>�����Մa����Y�%��6�u��j���H���8�~��bYT�o�m=r��r�&�C+9;,�`VQ�=Hq��
��6�-�۶�;U�E�Ǚ��Z��Zq�q�Z����>���:��Y/
�-n��ê�yݳ^��R���9�"�~�_��f=:wO	I)1�I���Ys?Zw}�D���Y��"b�TK��D��_K�k�-�i/_�r���M�N�՞c��Ii��K;7�f?NGَ>�Q�?oQ����T ��M%}N���rC;=ǀl0D	" o.���L���\&,Q��a�-����"&�O���Β�z=1�]GF}�1��5r����V�3Y���x+i�A�֧Q=4�*S�Im��=o�U9��n�R��`o�0<!?2�P��9���TN5tg6#6N��f4���>�_�9,�p�o$1*sǪF mX�i��'I�����"��� Ռ."�[�)�z���i�4��G�ٿ����	����l�a"�I5�~����=�巗N���K)�v@�6Pf����a��ڄ)U�_���č1���j����{g��GF�q.�{G!6�H��V�L- \��*��ct.m����I�S�~D�һ�s���	Q>��u'��aCu��O�������BEw�z-n��l�hr����G���B;�`�¼�
��Cߙ��ޱ�V��F����뉕�+���X8	Y�ۺ�Z�:x9~Y+�O�"zywhTҘ���L��/���cr�>e�<{��70Y9W������E���^���+(n���`dD���Lb|�0֨%b�[4�Q�h�n��p�.���d<7{'XV�h+�x;�jǕޝJ�<:& X)��>w��&�|hx��rs�h�3���?T�j�]1���Pw�j��񉥢x:	3�1*�Y���|	W^�3��)6� ^�Kf�Ƌ� 4��b�ܬ�7�}�?Zο�:ֶ��u0����VK��9J�g2�!ί�w࿈�J��,X�(ºs!�pa�G�-d�m�q�D����H�yȎ�0\2}���2�����'�`*��PE�.)��E�4�\�2p;VD�Fg��ng�ɴ��9�,�Ŝ|�ܤ9b?�۠�%f�j�T�9q?@���>R�B�Y�(3h\k@�9�f��uj�h�x��,O>x�
nR�a�����.���9o[ŷ ����4���]yi� 2�"��^���z$����/C_)I�(ڜ�Tg�0����l�|-R�M�W��,B�KZG#1G��m5�W���<�鏅�ݿ��i��'���Q���B��(�Ҫ�����R��S�^�F@�����r�|>5u���SӹjE�J��of������ /�i?��om�� ��Z ��۰C��w�ɯ�d�'��2e>3��j�+`X2E`�ʲ�3�Z�t�ք�L;-X����&��cu��5�;5^Z��8���Lp�!�/��'4^��T��r��E��x`�,�K�2f��15��koH���AP��HZ�5u5�%�<G����N�J����}�~vx.��,�ޛ5��qB�-roז�P�\ax����;G�\q���xd�=P�Z���+�,/�J��$M���d���4�{k+2c8<�l�7�L+֤�w�
F�R��3}	Ps1
5`����Qo���\��>�U�M�����Y�Q��`���]�ƻ��� hj���̂���}�L���j�$c)&^C��;���ȨjLZ��V ��)� �\B�6�Mw_�j�v}D�V�@M��a�$%�R��x��
�p�=�R�p�\Z`U��s�o`��a�k��+q�t&������@� �|���B�&���3A���+�h��>B�G�}R��F�>�g AQ�&Ae�k������vi�qpG"p�kT: �h��6���I�k,��ݰ��mG�_��Sm��!�U�ޚ(v�Kaz[�u����_0=7�;KnlzO�B�] �r(�����Sr����	ؘMTzV�:�&�Y.M�MĜ�&�'�Fi�5�1�Q���'��[�!�%!��Aeb ���b�����q��9�{	�g���� �'��;�ϩi�p�T�%G_�Fo�b�*!Ѓ� ̊���qͻ��>V,�-��I�K\^�(��\lS�Q����
Y�z���"�_TȜ����Q��$T��ĺ�ӵ� �>��+��Y$|QD^hsA�
�o�1!誗�ȟ���x���.�Ŝ�Aveg��K�J����QE�U[�Q���]8�:�<H[]�q�s��&��]��m*j/e���x��:f[c#�����}�4|,ö�+b����#����IQqu�;�*t�6��߾�i_�w�un��/)QL��xT��HL�J( �M�K�93��Çx,ͦ��Y̽¾�cI���MEG2ǥi��q����A�i�3�VP�j]3;S�~���V��=���� X�]1��}�Y��`��/��!ش��yr�*;�ǹ��N>lHn�
���^/p������J�Si�k�C�=v�%���V-��Kt�WH����tl����^����c7�J�-vFx���U��<{�'��	�~��$�w�d��-^M��>�{�}�P5���Im��0d��3��a�����,`�OMN�K��ʴ�؄sG3!rȨW��-�[�i21��G�Tv�a��g��AX*/Y��G+�#҇�:VB�J������6w3H���h>�{ ��E�9fM��uELDv�:��K@��26��Bٷ�"���Dkw6����n�AuT�l�����v:6�c���j]8aL��9煛����#�,u����[��|{�4]���$iK<��RPM�O�1�sœH�]])�g!���M^e�7����E�)���E��kt㴈����(6
,[�������'�c1j0>�h��vk�(ߎ��Ewu���i�5���C�4;�\0�/3�q�R8�+P�X�ޚ�~]ꇽ�rk�d-jq9��`'
���d�o-�&��E�	�1@7	����Y�u٩�lRF3�t��-��A�z~�_�B�FE�P H�M���\JYǔ7��A�B�1�C�q�z۸i��oUv�!5I&��au�#_e��yPCsIi��~3�������{��_�G���T�#�p����	�E[���B<.�3���j�y�A���*�PA}u��E�H���x=���J��ܶZ�����n�4�vk֛���EL$����[�b��h��(�!�r0_L{֘t�i�H��ͩ�x �˪����ч3L����ˁ����UgQ���Z��NL������S�>t�K��fo�������n���e�4Ν�8���p�W1<�Wz���+d���F�������T�jN�߁�I#Z��5�Td�|��yDaֵ�`��soG�r6�a[p
p�lȨ�"s1E��{j�L�
�֒���2�2`��>}#o\�:�84$��{��IVt��	�P͘�a�=s�CY�c�鮡�E���8#������Q�����;�x��I�^�ϣ0�kp��</N<[i���6�9̓sf�C�B�І��zVSy,��[�Ȕ�	Ӎy��Y-�".��@�'�r�����
�H�лU�Y�ۧ]�ȁ%^]Z@ި]��]�I���JP5 ��&5�Th�آ1�gu�����p�NC[_w]]]�����������M�i���{{]�zg� 5�v�����jj��;��|6>+���%�1MQ
�[ǧL7��]�����>|w쇈�@���X(N9zZ�OF�1	�p��W��l������zw��V%���Éʕ����z��]�]�~!n�O����f���B�C�:k]A�B����6s�!����Ĝ�~+���z��c^+�*���lwl�B�,<%�ґ�;�-�>�{�� ygy�?	֡f�LO�[&B�T��������g�vR���oK!�A%U������U���c�G�l,�eJ�t�vR	x4x�+R�Ӭ��6�����3Y�@�7؛VT��U���n��MwԨ�[֪/�g�@P�QVr��K�-0��������\qȉ��tٟ1�9i\��O3!����e�<�8�:9'��Cb?�<��h��ˢ�:I�Y����S�nS�b��Yk��C�d.�+�_���_�@:9ޚ�Ï�����}n��� �K(#�=�Bk1c�݁t�Ԗ�z�q�LgC��.��Wd����Z��u��pC2�v�$�D#���p���	y1�T���Jů_��X4��q/����(��t�m�(rB��\b��{a}K��s|��`f\�1�f,u��I���?}�����:��<L`��d �1$S~4��ͪ�N<a.��'ZaE�}}3�"��
�n`���'R�"Q��~c�(a`8��~H2�@��;���K9-WJA��EQ	��ja��"��V��-�2��tUޒV _�+G����+�O&��	��t�1���.�)G�~�0���F�6	�pj�o�?��d9Q�ȴ��S�~A��Ef��s�~��j/�!�>Ms׸��{��_!l�dF�񩵚 D�>�a+���<;�Rݦ9�8b9V`Z��W�Q%z�\��FC�
�:�L�Ҍ^�a��È�f����adq�V{�a�Ԓ�Cb��US�B@`Y��3K:�Z�M�Mh9�C�|]Z���a����;M���CsD�0<�ƚ��O�kVe�����"��*�a�h��L'.�%}��3X5sL94�6��
8h���P���F
�M0<#���D�`��-�ݼ0�%#rܖL dY(�q�mg��!G�0y���O��$H�Ǳ'��U%&��jn����V�7L��%��V���,���'�D�&e��`�DJ��d�*��<-(VY���7B� ��'�cθ��,���X�Rܑy�o�����<`c�D���>���`��EjG]2ۖtnL&蛂ݻd^u2���
ZX��4#�Š��:�\=@7�0 ��g�V�'��],X�b�'@op�b���Jz,T�'�5�C�Ī[�3GZ*�iQv��"�ˠi��$�H�G�m�]�|��F��7�X�ܭ�ݤnۈ?(�U8&zU� ���J��gFt9/Q!U*��S��Eb��$Us�m�G�u��Ta�w�W-��4����0�.�@O�SN��Ƙbu �K	�l���eU)�'P�[顼%ʲ�x�u+�#Fd��+��M�*;?��h�	�,��_e��l��7^��r9 ���ߴ����z�2�|驭R�h��]������DLi�:K%�*J ��yW�-=����4V�]G��	��]n�3�I����;�[�8HZx�q�kua�������ɖ
�����h��=�����Ȱ/e����݈B�`o�&�W[�7�~yb�;+IUp�̧o�İf�V�*��4�]�Z	���:<a�}6Atu;��qۗΧ#��d~���9ъ�|��Jxs��8�z���ԹEj��QY3��IB� LOi*�wZ��Ⱥ���FaI[�� 3zH��x�$�Ǝ�нv4����0�*׺�w��e��-�[M�wV�'CW�z��/��$�'�h�a~�L^��������Bj��yJ)���fn1j��6�5P��`"���S����cԂ#�loM���]��/ƮP�7cՓ����|����K���Kh��ACf�%w���4��3<:�%,g2�
�����w�w+a;�l�,�+�+oKD�'3��g`��A�D��Z@�1�:�4*ԕp�%�εx��A��3�����_�D��(��6^4��#�
�H[l!�5�k[웍��j��~����桢��ɴgMC���k�߿ Q�ԉP��N����A�N{q�:yͮ�r&�go=T�^ˈ����!�ߟ�_UX�:-&��i'�cUgt8�#>�Ŀ^�}��R�� '�i|������C�B�=�2ВBM�V
������/Z��������Wa����i�����b[�x��F�NW0>��2�Oֽ�Y�S�+��Ib��EgI0
n��n	{l&,U3�< :�ܺ6������<�e�C�h%��Ѹ4�h��B`�1,l�	��뜙��ݮ�v[��7�~P���Ɣv�R5�߱<�G�Qp(�"l d!�nS>�dX���#��M���<+mh��ь���.���w��?�q���&E��gR'W�%���)̃��XZ�5�j��>v��}
��	NzP��<�����C]�a}4�/O��~|��e"��h�Qk�_���/9���3����>O���:{��P?��������i��^�Vm'��6���	�?��)��4�MO]L]sM{��A��ͽ�#���ELw��0f�?6�<O��M՝�h�񶔢�R�g/yܩ��XV%����Pt!6�?�8	<��ƿ�Ĵ���&3��Lc��K�L���K�7��H��˕$��������Kc��ʣ�:_��y�g" y�=ۥ��ϴ/u�(x�pN�ˌܘ{m0�;]O�b��.��H�����E6���	��R�z��P�q�L����l4�s�FVs:���n���m��nE۽��T�8��ڀk�TLRi8
��N�r���@��/;8sP'�+ۉ<�%�[U�o� ���q��<�(�|��{tT~@sP��Ƚ3ؙx4;/-�	3k�޲}b �������@��
p@��KЭ8�,⢰�X]dV�R�븙�f��^9�	S��h�<~��O'�3�C
�xo�Gx;b&�u5st@jЂ\��H��o�y[��bqD���h� ���
�YM���:��P�"��H�jls��%���m�A�Z�}g�p�"p�<Vx݃�>&�_�?ހ/ft�����R4�cr2��q��M��/�, V2𲿴�^���G���pA����E\�hm�M�M�3�^kV��_�^RBlG��=�y����u\���/�b�]�$xR���^�����/��rI�m8uή9�N��=���j,/�,Z���t�
���2��j��R\!�o�8b�+�m�kHG����K������|m�)��TVhbb�訚 �X�������e�
l�)��tɊ�8�<]��V-�Xl�,R�iq�1����L�߮��~0��q
5^�������''�8��H�Ә@hbҏ!��sc�v祼�O���n�	n��A�z\u�F�7.�� \i�V�C��5��bS��e���C��Z��Y{G��!�7����?���ח�(��~q�:f(=��<$D}JL��`�����636tX[��x�5%�:9��4���΍z�k�	@��6�y=[E�-��>�]�3*��k����꽠�U�'���^��_$|XZTu�PrV���&]T��j\7ؙ8 am-ʫ�Wb�����,_�He�6"f�N�^�M�휚G��*e@�3��7�myG��̹�rX5�E�����|N�Ƹ�b�Hq\�ͷDk��6��q9�x�t�@*��`��z4ǼL��x�u�k&2�Xm��f�b�y>���{RFQ?�f��IY���i�s�EE��˥�(��g�鮡����a�{D��SL��)�K~��k�޻vP�L8�^�K]��|��]{������Qg6���̎�Ud͏/�֕2��&��V��|�*+�G	/8c'�����7߷�\���LE����[�ґOj� �s�~�l�a���m�{{�fA#���/ ��+t�՜JY�l�~|;���|8�`�ՋD!T�3	Xŵ���^b���&����W�6�#{�J��L�L:V��*�]Bߕ c�O�*���^���O�qj�uC>h�`��exQ���2;�zT��j��cd��@.��;;���/�<�P4b8��M���Ρ��ۂ���D�8Q�k�v�iU�(4`��a-�(�����`	���;7��IN;ڒe�u�7:P0�As}檅P;ܯH�Gt�^g���~xJ�h&C�6�J�
�:�,��yW���g�r����	Q2����/z¦����}���)�]�K�@��ܾx.ݞ�"�����A(V�J2��@���^���W�@���E�-ckA�sv.p2dr6�tf��I�@�7�n�+[`%��N��t1öX�:��?�{��j�T��8��ߒ��T���'l�����S1�,��)�׸�D>p����(H���X��Y�iH��E�4:��	�e�*x���=���H�k�eMhE�-�2���0����	�)��6�$m��b$�,�C���.�*���_�L9mV.j4{�\�Dq��<L�Ћ�l1���Ĝ���P.�.�@`і(���Ӟ {/��f0� ��@w�ǻ��N P���`��E��кi�$�8����GK��1vﰨ<��RMj8�?��T��������s�!�59��C�)n&ㅨ��YkȖG9cD�rO�-�����������'��l�6���P��=c��S��� 	<]H���t�ɘ�y�.��
0�޽�>�Y������G�\N��vd�:�kK����8M7'{��c>�_'�zǞ�s��d=$�k�U&h�M����i�u���kl�j8��8�+�gd#�g}���C���d��9�^8X��Iv�ɔ��������V&A�w��I�\�&�����N�f��#H�%�6������'F?�FV|O�I�W�m`�1ԅJ��������������B���T3M�]�M�Y�W��4� $�J��z�m���e�h�euN���"���Io�7��	{�j���R��r@Z��!Dw�����_�f�b=g��p�&d�>u2>ѩ���4�oc?}����#��e�`��18=�7�����HK�$IҶa��uku&��j9��d#zem~!�����kc�j�L��z�����,Om�U�q���e�45���7?�I!����&~3�
�n�}B�B��&��j� Šι�2^�>?���b��:�V�=�
�O9~��J3��1Fޝ�ߎZ�EOZ�6�-��N�7���d۶����@Y�t3q��O����I�0\�D�3�D�ɣ6� =���1p}�+%Q�a���/�����\%vtw����,e�\./~n��_�RȆ^&�~:�9��b:����r�]���
�s���M�=�pS+�Ԇ�8�1M[_']}�<������A�öXw���&g��~k[5zA��2��dqs_QG�Y�z�$F���ʐ���Ν|>-�f�!_)k�ۂ�C�.D�(-+��s��Š%�W�~ۃX�F%�z�]c������p������������|J��dHS8��
}�?�9pЁa���N�'x+�D�%���?>�z��u���<Z�l9���88A*+�f�s���ײp�1�y�Z��c^@r��[ɽNWm"����oi$��/�;��#4�ӕ�2e%]���[u#�T9���d�@����`��%T�cB�Z�=%�dYL�.����h���0��/Fg�7'@���ս������A�����I;���Y�b}N]Z���'��Gٲ%�w@-�����C\����-���l��M��'�6��~3oCV_*�KϦ�lC���K�3(3V�[��`�i�ZP���#��
:���CMD�F<(�QO�P4�@��pF�>W�m���v�o�\�(!lb�YJ&˜,Z��m�z� �1zKrp<�Rǐ[�#b��D��ʷi8=���Z'YP����a���v]�զ�.�5ԟ3�Ja�]�)��,����L��='N�k@F1pMC:��^Q�K�%$Zպ��WI9���8Ԑ�4�z�fpX����!%��^���QU�<���tJ��i�"��I�V���ֵ��26A8F ���`�qr��qx�L=�L�C��X	��d�W����I��i$�9�QH�ʒ�ĵ���ޜl6� 8��;<A$� ���N��I!��v����5<�]@�<���#I�(~J����)�-�}A�Gt謜	�����y������k$�%˹#.�yr*�>ϱƣUS�C홦`G�U�Pd�]9UΞ^y]	��o5��}ٟ�>����7�}?�b�[8���FG��?F���sXg�bH~>�|�P����D�Q�=@Cd[�|�Qs2�;����JU�1<QC�r��6?���	�Y5+e�c G; �-ǤW���&s&��Ԓ(��n�*�D���9iO%i�r������vB�JUVҁ���F?�N���g�/T�Pۓ�u�ʃ���۴��,1D�N@!��/ޖ<%�7׳� ��]�X�\���+ւ�|�Rxb<\�<o��r^њ�3&鿡i�{0Ha�Ig*�^�_|��:v�3Dv�&kK�/�r'�c�u���Hܩ8��˰T�Z�H�!�J��@�R�Ы
��[i_\5�mk���#e�6� JcS�T���ƞu��Е����s�L5�r��,�Bg�9�O����H{�"3Xr�f�2ah�[�@���2�btJ{�M�`TE������tDv�g"�R�V�Ô�ڽ�_�hm����QZ1�s�D	���]�f's\�����[��A瘽��eڝA�lZQtA�i��I��?��(]�B�,L_X,�tf�f�P��/@�Q]U��Ii�L� ]*�u�{d)�L�nNw�l�	������桶�}n�7�ؗBe�u+��
���q��5��n���Fu�ګ���s�rL��o�}���HB	o5S%*|��a~P�܋[�1ipwK��ȵ��
=g�d�S�٩�P7Þ��.I0���c����`g��X�gp��yL@���s���ğ�f�~\m�]i�:z1������H`���{�ǻe�]����^�$ �y�]~��੼ك�,G U�)B[P&�o�Pt(����zjW���m$V6P�V���1dF�L� ��\��4�ŪG�!�7�Vh�!Sv�?o���ނ��60UL�7ᓺď�t�k�LJ���(�-�:Y�,��f壜�pV�WpA-]����~/�iI¨��W(K!�}1�K��ZS~%T1(|���B��<�n<!�J�L5\[����Q���o�:��}�
ȿ�D�Q�3��r]#�ȁ����oHb,���V	A�g>&��������z_Z 	�0�54g�o� iޫ[k���&<3!!�ܝ�<�ͬ4w���b���_�����_��c2n,��/!'�Rd����I�H�O	x�)@1}�YP�V��Zpa���/�D'�,���T���b�r�r߈v�<�ZUzw���Y0����z����MU\W�A��wfY'+c���~��α5������G���l�A")A��N5�|�����Qfe89wD�nC��m�c?6�$K[��`����#�0�X�/b3�4F8�t�q޿��@��ogz�9�C��*�Hڰ�H�x�	����(��{���>҇FA�7k���޽J�1AyB��$L2�PO���c����9����]��!z�TN�O��scp`A�RX�b?Y$��_�s�&"��~�-��;<�ε:�a;�ap�U�����������#/-͟l���_�-���<����/EY��p#��J�!*��bSD&��!|r�;�����I� ��&����~m��f����*V�$�>�=w�|�}�i>���N���8��rw��ȱ*��ke7��8����Z��Iv��ɘ���wQ��k�S'Q�스3��X7����A�:0�r��a����5g��7x��n��UB������ZH����=,M�m�}�Þޡ_<ۢ4�>@�^d>X��Pkh��n�5p�oF͛�R��ϲ(�6�u��h�����$�7N��08-2Yv��O88�%gD~*M5;e�{|��KH�ԃ�=e�i�x�����Vn��긘�7L&�;ݲ]�`|^�3����r�(2�ϰ���_�l\��rq��[ �#a����@�.I�[C)�(P�W2��������V(��@�=�z �"�*��J�Q�q.�Ç�yQ�'��u�<���"Aa�C�{����u����V<�r~��ȕ��4��l�8v����3�{6	�������vg�P�a"��u���=t(�ˠ��︾'&�%K<��]ɜ��$(�6�[a��5�;"��<4�$pK��aή���s���c��s��Ђ�;�6����WgQvV����U��'�����*=zϝjC��sdc�]:���0H���f�����00*8v��.�lpS�@���Z�D�o`�3Μ���>�5�#���,� o|H��e ���W�5���?��⁴�1�U�����q�톸.�I�k�!Y-~��
\V�_��f�f?�댔�:1G�8��J�kؔBi�ъx�k�v"�~��e{����8J��t�]��ɂ<[[َ�a�Ip����' (Lf}ɯU.��h�J3�.�LN����$��l���/�[F	p'S"u����~���]t�e˟]��X��Z��9Bݩ��	����Q7ԑsw���Jյ�*����)��\��6c؄�H��v��k'�4��'��s��{Nd�wv_�r1���k-o��f|< �|�W�GӐ���S��[�K�=/ 3�Y��F����ŉ�X��=4�] ���<�v�=$��㬓ɘ��W�n���-B|b��A���%�=�x�������?2��M�ȳz �փ֠rr�#Fr��X��Y�nr��3{�2Ca5T�������tF�#/;�j���UF��ō�KOK�1�3�#7ٍ!u�Or���5�CːS�\�;HK�v\�H1��6E�Kڇ�HنA!�oԎ�d�Z+��8�i�1y4�.Ğ`א_�U��YȀm��!$�"y�<���Hs?��{)�|&v�|b�n�sR������ S��m�Gfka|]K�"|��w�Ӂ�%���ٌTc�>�~>�{J���yA�6me`H섷0�sN������a�hv�[L�]"6�o���7��ˮW�f�)a��g�I���7�L�K�9
�J���L, ؀�]�_K�����*&�bv�i�N��+����{�z����9/�m�DY[F��,�y�?���wDN��LP_�WI�6��ܰ>7�<�ޡ�uc�U�'�4�w�Ί"|zzUD9�����~dsg���2���c>Wcb�&2?�օg���⁚k/��j�[�Y�#�N3ϼ���g�F,�}�.z7J���u��\D�E!PKq���Ks6LU�\S���z�i��o�!`)!y��]�B���&�~���N8��� '�ې����(���/wK����vҋ�˥��K�Bv�h ����"�4ﳾJ�~�Ǆ#*e���[�j/A?'��]�fէ��ӭv3��"u�nX$���j��5�h��ξ�ژ:����СT�^k � ��Y.6�=X�O@J�r v�(��c��������t�� f��7��%y�y��-n���dH��COޥk�p�}�3{�Wn�~�����_N�3U�ؚ/��} ��{6��S������'� ��	�RMF�a�)�
6EHD��#�ۙ�d��8�W�����bʰiR�![�Ȇ���}���7�2��DJX��!ٚ�����d-�,h�w���	���;#�c�ۥ�J
�l�����?P	~��4�ۅ�+��҃�	o��^��|L��ڜ��ɠ���1Ќ,:]�Erx�G�粶����GI楃vF�vx�a�n�!|1�O	�b{3Ic�i�ϗ�G<�W��](���w���'5���d�4��d��!�Z�0�y�J��R���HL6�`#�QV]Rl��+>a���o���P]@Up���E�&&����C���Q���/?��p7��<��[��IVջ
U["M��z�]�_ߙ��}
�Y�BD��ѓ���\y[űr�E�a�Ӝ��b��m��uvs>�2!�V��H�&�~ϱv�o��G�/������c��u/��
G�k�Bd�����4����9�y#;kp4������c�;̞�/��[��1���1�QS�>�D:�;C��WU��s]���7�ч�2冥Ֆ/=�l��:v�<�ys_��m��l\�%[փ� ��Ý���y���>��s]MMD���\LT0@ѫ�W�gE�Ʋ���r�N��B2�9��P�5�jW�c��^A&2�H�����酊ʸK�^@T�v[A��_�ba��q=3b��l.�יr��'�&� ��IW�.�3@�} �q1��P�dyʙG����I�y�+��z������Z��L��(��� ^��ib�аU#Z��Vu�2-��gf�wC�@;���q�d�j'!±)�MNF_����{]D0�41�*iE�|���f�$m�P(L�=�?�F�z9:fu���� v=c��Qkg`RK@���2��f�3 ���n�t1e�����8l��+a�+�8AW1�H�;a�M����$!C���}[˱4���a/����4�a\�cZW1H0>ڽ�BM��Fz���]c�W�g��/�\��8��~��|V��)������W�wn��M����H�j%�1�B6���l��v�������B:` �"�oK?[B�>��'V���^ ς�D�V����hU��s�2[/7Aw1+�(8����,X����9����`��QH����<�).#9����^4�57���{�UD��LOCގ7��v����6�v9>�pҚ����:�B?C����ǫT���]�a�>\�/F�܇z	���@]= ���C�k:b-�6\�f4��_T�t��	���a�F䷛2��Êlb��n��Co�+/������Ӷ
�qFw�^]�κB���jr�4�<��������[V;
�u���K�I���Z��Tc�w}t���9&H=��#�0���5��9����͟bW��P�T	��F�B&�:۱%�W�����S�ݗ���N���{��X���ѭ�e�6Q�#^
�3^��ZG��m36]���w0�=g�HmV����5���u��#g�l�HN�:-����"+��ķ��v'�α�HЗ�{�Vϛ7��R���n�8ڼ����=� ��1z\Ts���@?Nx�;0�吶hV}��ش띏t~'��Mhx����:̂�XG�����/�o�Ŗ��b�3��"�Օ��c�� �8)�Qbt ����^�G�?2���J�_�ۇ���,h�t0�xɯ�LyS�d���>@Z��Q��.�ZO��df!��Q��{�s*s�O�����H�����X�6�~ê.{Da9F�w}�x�;�o���߰����r?�I˻�)�����-�XsV��?�8��U �� w�N�	�xΖ��N��)zX�@����;bn��D�,�y�G�;͟�M���F ��@H!*9�J̵n ���7��_����=)woL�!�r5�R�"���J'��J5� w-��_��tv�Pi����*� � �=J��l��a71��ӃA�^���|x�AR���g|�O(X�v2P5!��@xœ�!���'�h.wM�XLZbx_4K��T�v�����Cm|z�+�5,� k�#&3*ŵ�����ld�R�CH�|ưX��!^#\b�^bFd�v ����ܸӖR�u�x��2��7~H.!�w�bCA�_͋���J�����*�F�(��E~_�/��F�ủ%X��y�EZ|�����55͓��A��)�À��H�j}�4�4�7����x��b�AMD�ma<���iB�qD4��N�d���.�:�M����u� �i}�?���L�������H�ǚ������4����>��m�	�Am�b��2>|��q�o���k��
Zץ�4"�-���UoVr�Q[�#ZGZ�kre��:6&#/�o�gT(X�!�]���&�m�_��1L�x��������;HEA���c��N��yS��2ȟ6cC��y��O�wS��i�>��..mḲ^�r3�M"�����`M�`�ery�N;�4�x�}��5�<�Eb�"of����r���WR���Ld����(?��R��:'H�o���@9�n�b�o'W�&���epR�,l<P�E�+O��V�����X��������E��kQ��=�k��l>�.?��
�ψ�B�-h�緝��.��y�i��-N� �D������|ƴ0�D\XԹ�0ˉPAJ�G�}ߖ{5 ���(٘, i��	bE#4�WZl�c���p�N�2��p
���|�רI�G����}=���hK�g�Rm$⠙�8��.e�uT^ϥ-���5i�N�� �aQ�U)2%1p�;�Йx�8���:�%[�1�6�予M�@5��W$��)�ǣ(��=QN;��o!	|��	���Q��n�i�ͭ3�oM�����)~�$���>td(SX4w�/ ��$"V&M�^�K���nƺZ��%��jq+>��c�V�(���˶t��6N�>�긮+V�KEF��>� ~++b)hޕ��.
RSoU��{q������&ga�>�Ēi�ߜ ����Pd�NIx�s��,�kل�v��l��E�!��W4H�'_��G������V��o-�Wk�xg�����h���`�)af1�X	���1�>�tg�n'���`�i���_UuV�7�0cu�/ �����~������~����,�*C�q@%��%�����b�5F�9��� �5QKD���O �tA+P7�_{����lP]/������:�2�!�?��z��$���VM��/y�zީ��S�X
�JHh��%&z�t����-b#�`H����(�ze�!f�t���c,;��NPD��k<$_`Xh�I�ֆ�;55��%k6�D��������O���HU
��o���yKb~[
�b����S.�f]��4����+��H�J���b����?�����j� Z�Qn2�>�j'����X�xG��< g��=x16<�2`��x�5��GL�9�H>����r�KgX�"����*��_���=oj3�Ĭ�e3mU�e�4n�?��������2����{����(��,��f��������|З7=Z�V����m��G���B��6Ҧjs\�bmO8���l%�yjg�\7W"h�yͽ�^�v~���d0n�Ð68u��y�p�+?��Ȟ
]��P:gO��W2��i~Cod���AԷ�	M���,f!�)�xώ.�|]p�ìv�����+&�4Z�P�T�Pп`N��噒1���yV��������m]m�L�q�z)EO�@��F�(/����|h-�J��%q|_�`��r�G�	�=��XJr�*��K8�ȖF=��D[��3�C��1�?�*���w�gc�����>2����p�Z�K�.���i$��G�i�>;�\%����	~c��^|�f0�n	��ݏ����MK&o'��j���$(A�n*5�R�կ���L��aT^�mU>�Q�>����Z!HdK}�l]�oi~��!˿L�����R9+F:�31��F-�R�X}5�e
U�b�Z���?<��Y�����Y������
��Xo-�){ٞ�Ź������HH4e��'�8Dƛu!�v��'�v�W��{X�Z��orɟ��~���O�0dRp�Ir��>�N���s9�/��G�������]]��{�M�8^��K���JU#e�]Z�o��n��}b|�p���v�����c�n~���«ޠ�����r6�#�&a'�V'��3�(� V͒��`<�M�|m�dkϠy��V��Ͽ��U�o&;z՚!���f�1
/f�	���'ڌҏo���=:v�!�0Y4��;L�^.^~|O�-'_�n���S�����^O��Y�c4�A��H@8������	z�����%+Bb��u]`q�Ա�ța���L�p�B�P.M�9G�)�#Fq����m6��3��~�y���
��(�䳴��oP����g�b� ��68������x岤'�	��J�ѡT�bnX,�^�2�0�b(����nSW�f�U� ��2���Ҏ���U(��Q��O���A^�Q��c�j�;5	�G���~�<���"� a�G�b�"1�D�FɊ��	8?��R[�����UP����z��
��G}<��&;3_j��0¡�x�ށ�4U��㎟g�n�t�#�΂jB����\��^(��b��SG퇃>7o�N`� F.J[<��Sk�4e��g`ku�m֞A������X��Ɍ צ���ÅN�=��$pCׯ�P�`⻴(��^���g�5������ �����G��|��q�R��n F���&5N]�,�\hג��/E,��g�n�a�V0�;��t+|�}�H?���7Z�ȥ?��ݶ�j�f���럫"�:��n���ap�(+*-���&��
k�G a��uP�yY[�gJii�]o�H�+�"�'_ܓ9��U�8w,wP��}����oU�S!�H(?$KOP�D����&�w�fq�	�#1iG�^>��O}��M7L
eSc2 ��km�}`�Cx�@?jP���"�;����������ŏ���n����8�~�>�_'Z�M\��}���$�xULTW��8��Q�k����	��5��N��5���a7�j�vc��/0�-V Wmq��[�k��oU�Q_4�(��;(鑖a�o���M���V?lM/��e\ٱ�J^^b
��r��v����`��Nr)�*w�vY��8�P]?�I+��z ����5�����6p3iڌ�l)i��O���հ�;8���ˢ������hI�� ���.�iU��GW^{�����M��3���)��T%�%����= ^	��?k��@� �����q$qY�Ϲџd�6T�2LN%�ؚ7|7�\$7�i�#'�x[���1ݴN�Vp��N�����<ב�}��.r�n��G�KFgő�хDխ�9����Z��[V�[�M����v�
j}��v�SN�^`4/h�\z�������iK�Z�rO:��pX�h���C�J��H��Ү(�U�f�H�,V��,'�HV�n|�k� C�1A@�щdſ��}��fs���?Y%�Pu� �L�;XD�S���mХ%�����dJ�W�1M6E &$�q���\����"��BWn�m+�	ٜX��SP�����'_���8r�O�AAX�,�e1��v�׵�~V�Y��b5SN�I5Yg0a�C9e!�U�Ej1n�'j򯘒��p���ߏYu��V��Kz�?�L���+���,�m��m|��Kb��0b{���\e-��&�&�f�>�"�R�X_y����WH���z�K�e�*5�m�,�\��"Aٯf=[��C���Fb>5������kd|����ós�� �'���ik�\�-�O	tJ�g����~DlB�;-G�XU��V\Dq�T��ה��X�a��W��i&��@=�w�h`8���K�f��ӧȯj���,g�b��
(�Ϊmg��@����4g��6�(Ó+h��6�HT ��q���G��h!�,�Q��&v3�A����5��B�̖Z#11L�dU�Q�9�1��(���ځ"yj��j��W-��x�����W�^i�����˦�G!b�e;��j�̚�e�(_���V�ұ��y�X$E{��ɣRws�o%KЕ5N��+̕R�Y��m�������f��CB}�	#@�&�ְ�UG��4[@"v�*({�ʔ�$����B�l�k;D�{�{�]>�Ky�*��&�i+�3�&�{�'�PX���zǫADA?�ˈ1r�Y��.\6�J��ޡ��J��f3yBߍb�;#��I�VJ��=��_��B[+U卖+Tˈ3^H��v�,�S�i��-˥u�o;+�+���_r���4f����Lo���uU�c1g&|��=O����د|�?Et"��#pP{�g��X���r�w0��j4KًH���b�sV�@�б�I&Yޤ��s��H[%C�>�7T�8�jU|�uf�,�8�����eZ
�ZǊ`V�X�(�D-��;�4�F��G�){{Bb�\������L�K��ΪZEW��xrҋ�n԰�$���~#�����LK��02���E�����v�ы�����o���i�T���=�b�U|Ry��vb� |c�G}?��
m���y����j�����Z�=����iӺ��z��4���Qʹ�_�RL�3�{�S���}׫�Qaǁ�Q�̀���D,��7��=�ï��x9�Ď���=i�����+��ղJ�cV	������{�864=�!3�NϝMߠ*�ZT� $�� %ӎLddF'�i�)_�&]l!�'��������wϨt�ܝK05r��pޞ���d�)5���T�<��Sw�k��g
��*]��9��Q�)#���cB�
������4E���o�cf'Ŕ��!���I[9f�Z�B�'�[����P�`lM��$_`�>�!1�#}� ��/$�C�=�OZ'�	ځKD^�6�_>�"���?��&5CEF}޶^A���;���{_�q�3��,>H\�B�i�Q��-!%����X`j�w��e`�S��X�{Bݿ{��Q��^#����a��k����ԏS ��W���S�^P�ct�)��Q0�v����in��:8A���@�bQl��kz4�s:Q�_E�-ӫ\��SZ/���O��ؔv�����?�n/�UUʒ���<R ��b�� t���6���RO�5����"c:)2��l[���*��:e?�)�ࠟ�ݴ��/`A�����R��PeT�1���YO�:~Q	�a���5L���9}V�ɫ<�5�K�:���c�h��u+ӫ�}@
=a�_��˲�f��C@[QL{����s����w����H.dc���Y�5��­�R{Z?��� �˹��-�sO�k����[���Э�|�J]j�C��l�hG�E%'E��vC��cF\�m� 4gH�����8y�d?�D���K]��ʅ���!.�z!��o1��M,��޻�9�Z���f޳��}K�\���킝Gd���Gt%
t���\N�08�	�ĝv�8�� �Y�O�?�Q��J��A{W*�h�"�Qf�zڴ�l�UF%��F3W7e�bCA�kj��_D��uJ�Q����Kg���K%%�`�;@LH`^������Qy�	V�om7�<c�I&�P(��Hy~<����{d
;��;��<c]K��Z�Q�d�utl�Ɖv�`�d�IW{{Mv��_�~҅bƠaoh��-0c$��W��B�3f@"���B��=+A�4���m|G�Z0���,���Z8Xa���-gĀ�x:��:B���S(��]o��S�4ּj����ٵr̅],^�E�1&2�$�c���с����:5r� �9��������G�����M Y�t�s����|���|l.��+�:w�w���Y�s�K>ɔ����:K�n�����"[�m�~�6�Mk��W��?2��S�z�à0�jκ��DT��@T�]���틢w�)/	;P��}���{ahJ>��H��bX]�ï����p.v�bF��3E!/�;#3Cjk��Hv7.�I]j�,�������j�����_�>�4d����kn����a{:�ŪjG�{3C&W�4���x���*�0�)��0��T����s��u�B����@��NR�,`3�:!}��w���0&�m_����X#������0l�>z:�j�ꁉ8 o�a�Q����H?jWX�����Gr�����U���&���"��A�%���ՒI-ݪtj���7C��}���=�r�>t�V�Ҏ�3�6iN��!�o�&���!�̇�~��0~s`%C�������ME���V�"�3PX�,����#'�k�cN�2�O�&6�`�͞�������g�*{��Kg���}?�q�>|���������?.K��$$���0��s��I�Q@�m�������$����66( �u�O��&��+���i�����%����q(G���V��+O����g��66�Z�:�\q��o:���8���Ŕ&Kgl�]D��A�̬�ǏӂB`-�w�)��?G��	\q��r����p���]����c�{*�^�l��7�V�'�L0�|�f���m:꼴�Z�>Sl������wV��J	�}Ch ���7	�~�&
�?V��9�"�Q3~�5	�A����;����i���)���k`�KV�JY���B�������Cd��jk�v7��r��a�Q�7�[�=��K��h���j6lg��8>f\��
(Ƭހ.�.��%�]�m�z���Lb}N�a�ٛw�Άh$��"�������j�S� ���w�'
�mt�c��h�e1��~IL$pPrί*A���{{_���-�U�,�Z=�󮪭��y����e��W?^L""�$Z������7�ix��߶��ɗm?d��
�b��2�7δE�|#���	�Q�**����H��"�ڞ�X΃:�d�l�1k�����"�h/��!�z��Kz��G�7�����7�7@���"#us�RM�l��7L`��{	1hˋFUA$"B�nf���e!�.}���w�C�NP���T�h�P��γ���qq�Gv��o� �n�{ �� ����}dzV3��̣l�g]��m�Z�](M�+�/y a��p����>��8�:21H�7�;��{�
��y���Q�æ��]� ,�(X�i�
��"&�=x
*�:��8,�(;]Jб>@bc�W�.��ĶS�/����c�
N�����٦\N�H���픩FX���wMX�\����s�.Ɯ����9wvk2� %�S�X����Q��Q���W�gl#�'|��ys���Թo�[6<D�V�*:DH��C�����g��/���΄�*� �y�X*���H�t�����ݴ?^';c���s��B���4���ewц:�詼�Oǜ��2Nb���d�}�����%�)Zi�g��\K�����8e���-�a���Ο*�<4�Z�GB��Sؔ�`��9Ӽ$����BZ�ba.j���]����l�
���?���v:��u��d-��Y�jT6�o��m�	��'�Y�ST`�u���{%~6�^�Ҋ n@����_+k���h��#�}�T�ԑ�^���t�J�����z����޺�$p��\�Ǽ*h�1'Ϥ��B����L�$&$ϲ�*�����Orʂ�����}��y&��v���j�O�+�>Q���vLC�j!�_V!ro���2��]w��d2lC�����Q�̀�j�uu���U{�>|��/��%��g5:v�rY.�ٕE��� �~�G񑃷���\2Q0x:���Y���c�o͕8>=ڝ�-��J_�u�QuK��eb�֛���?�X��:Y�;EH˺���ՌB�XbJ�������	>a�s�S�^������������:��o���%&���ݡ_E$i<�����-\a8����}jT��LZI�I�$����ŭ�Жu`�#����4�3gMՆm	[�3r��f�����H��셛��~x=IFr����$���	�����-Lz�.-5�I�Mxs����TO���H���3D���8�P�\?���Q��{��ur]۶��8�1L4D�\�U����Z����s�U�>_��L0�L8j��*��ǣ_$�@=a!�L��=���iMR_$N6�t���)����)���9�/��0��aOa��ڝ]/��$�OVwd����x� �*-�����Qяp�p��@^L��W50��y�bƵ�p��44��9C�}H0��)�g�v�%�a?/�̭��}>Պ�T�� f��V�k�e�I������& �O�p�hn�Tm�	���i��ߊ`��4����2��t��K�6WQC+y���x�'�k�is��Xp(��>���&.����l�f;Zi>2�����?��o`S�'����e|n�FL��?ІwC�f�N���C8���&���jϗ;� ���S����/	��:i��Z"ȷ��� ����p�V���8�j9�s�K6���=��^��x��vjh�nbcB+g�m����\�v����8��jə�`�~bǼ�����ڷ��y�"z5G\�I�|)Z$P~!�"Թ�'}�p���=���8~`!ca���fAa'�7�q��ŗ��{������
i��"��x���3X~��aJ/������+�����sJ�f��4�W9Hm��5��oSG;8�q��D3Jq7�SS�}�!78L���R��*��U,�i���<��4�����Ʃ����%�⒥e����'���5sl1�Y��{CJ 7I��!����zT��&Ͳh2C	?YW3�#[�H�`Q�W�Yqh��\V�8�u�m�S���ϸ�d{A]��
I�4�����aO���M�X������o  ����a�?`Ȁ^��A��Q��r�u�L�v���4Y
��,�)?�P��#&1��f�T��w:Ë��
4ؠ[�e�;)�u�R�	{��=�V�.�D,�u$�|�X��w��e�*1�qP���2*�9caIh��g�P��[F�(7��J��hd�T�~��^iOb���dF��e��CN�8,99�1�>^�ߞ��"�����u;������כ��Fi܍Ĳ��"'e676�;=|�s��`�D�Y"��H������E�^$j��	�1"l*k�!�K�糐����0qU�?O�䊁?�}Y��$�DJTd�uAV���I2]<a�v��x^]��̈6M`��	;��g���TX����~*�"N�Y�[���w��^�2%�a�h5�լx$.6� ��).=�)Z��)�C�"��!��c�d��]�a@yxn����StZI�C���U��5^.y��G>�A@�wϚ���wYu(�+M�|�O�� =���%������M;�7C�a0��2�)�MinV�=,�m�{�0t��#�C���FH�bPh����s�l�*�1�4=|�Mn��������֎���Ll���/z;B�:����7b��s�%?�Çڄ�$�+�?������[� �s����qV�ԗ���4�mʹ"��,fBm?K��m�&O�U%���Śz܄-�ա�ӆ�ȸ֒dU�e�&�Y�&T��M'W)5�ce�H.�$� ��?U�b�����"�F���,�O��^x{�"�
I	M@!���?mF�?�$��V:�ff�BoD4������ -Uqj����%�=$E�Qu��+�x ���Θ����4#�����B'�b-��3�?�� ��<'|ۛWG4������,�����������0�i�
�fku+�ҕ��E�Y���>��'Rτ�7x0�IֲoU�Q�tQ���Y��Ef8���wN�2^p�L����e�3l�YC	#�j��h��:�C�{����'R�K�̈ϢŌ���Aѱ9�P���<,�Q�;6j�1!>b�`���9_(�e��K7@;)��k��)�#�3* ��$�x\N&�ۿ��sV_��i�������6��`_N��:'g;��J�hE�$�L0K(=t>���[�f�,��������Rl�:�]N;�Ҷ�f�w�U���uU��x	�����5��8�&�DF4���Tz���=�m1�2T21�?s�D�����R�A���@��ҹٙ�ac�v%�WL����}�aV�v�O[2���}�^f*u� ]M2�]�k��$�ᆌ�",�Le;�S��<wA�wnJ@��/����8��C!�j1����t��7��	(�,g(z�E�y$@`C�����2)�XxN-[�������1\HM� \8Ԏ$�B��ۋ��q�J�E�ύ�9��=���u]u���օ>|���9��x�ØWWD~?��c���E߇��h��)�&}K�F���=g�{��a�<��܏K�qF�5u��/�	8m��zs��dpb�FϋV"$Q�1���uԇ�M�
@��1�9��Ƙe�b�ǈ����q;fl{��k|���<Z j .�����%"���(tOД[�c�Y�*��R©��b<D���򩖝�$�'��S������e�Pzr��ҽ�[���Bܻ�O�2+��R�&�D� 8���-���5� r8��?���W�./�����v��'�pY�;{���@'e�nO�i�5�[r�b@e+�����<]�:��ɸ���۔]�acD�q+b�޼ ��O�}z��m��Q�E�V57s�
�$_TK!����k�����(�����K��0�#�|RtVc	C��^m�I��,.�&�m��H?i�0����[�(������Ke#8!0&.������@s�X�q��ߺ�i`4*� �(J#%尳M���Z�F�Vx
/�W�[���U#��̛�����+� ԙWi���	8/>Q��gxV�_L���=ʔ�&Ƶ�w��[�)]ݫ�㣗\�i��q�3�'X���m�%�험�������"A��^|�� 9����^��@m�0��M X�p�yW������,�A�B`W���@Ɋ�ZQ�h�[Yڐ�	l��jZ��Sv�|�죌�}��9og�c袴5�8�nQ��-�V^]�ε�ZT�O��1�Q�2<��k���,m������S��e�֠3�9Hz���C� ��l@�H����Vr���%���$[�E��Q���
����_�H����g���ĊH�zb�b���"���炏@ط���W��$���pL]=�������(p�pI�)O����jO��KF����-3E-��)j�{���+W��!���MA���.zʊ�����O%�L�@r3���8��y���)�ɟ������_��4�� ���
�����`�ƈ�)�vm?a�%Ɉ��" ��w�B7c�n愼1�-Od�ۑ��5�.��s?u���/������\��ԝ%��ڛ�R ����ʼ�R �ʜ;d����*TFp�{\'���E�pl�1������<�WV�i�6�H�X��^����m�N���W���Y�c_C�mMZ�N���BY��l-2��Qm��L��D(�N��7�bek�W5dy�޺���I�i�cc��6u`ӜvָR�(�A�E�va���_O9TQ�|���0vB}��
�a���ޜ�:K:w��[t��.�@�ds��jJ`Rr;i��R4P���h�7@�?�����=*�N@�*��?*�ӣs	�U�)�����@2k>�N%a#q�4ᾼ���U����,af# ۾#���O����˴�A���)(�!�2�(�(����1+����ծ$*q?�M�����N����b�?���1}+��`�A�_����� R��mh����RZ�-��|'�	%h�Ld��H�c8�]%(^�� �*�=ڻ"��&P|2q��QR5G���M|�|��y3
#M�f��I�Q�ad��;�i���XO�6=�}T�9��.4L�5�U�>�7E��䍝�^Z��>m��K
���/ec��I������Kc��@{X�*A�7��Kr\����8��|�m�<|�Y�s�¼�/gqKH�ֱf�=���я=���.����J	;ɐ�;,yf�!p`�+�,B]�0�jF�*�)z�X�q���D�UB�����j>|�Y1��!����+`���p|Y���@�f�3MI��#QRB�_�{�Q�JU��������fPc*F}�MͧP���3(Eb3�=� ��m�˳F��ŀ���AO P!,(���B���*�ơ�}�t�	�=[�L�c%�e�U���L�!�-�@8p|�V^�O��<����� P�-0!�*�����i������z��~��Z�I���{tL�4&~���T=��V�2�L�q_���e���P���Z<��M�sQ�RЀu^��W��!�]_ˢ��C0������8K�uW�],_�B�'�˱�7��C*:��z�U;Ɖ��(��9�h���&�W@�$�F�\�su����0��������e��/��O�Z��������'�ɩ��,�S�-k�!l�_�0����z���w.$]�JͤR'�_���s��*Z��ܙ/�G����(|��2�?{N���p.����Zl�TI��vFr�l"Tt�����#Ti$�R���-^��U��֣0�Ŵ	�Ҩ�+`F{"X}��.��������L �z@{)SQ����RF�Wq��f�m2Ѷ�^|5K]#''+��R�d�,�>`�.�E�\�8�}��t�Dnkh��q6�#@�˵&{[��WB()��_��$?��︳Q����;;Ӷ~"C����TM{b��B��W�+<#���i�Z8�~5�j�
?ğ�Yznql;��� ��} ����}�l��Yy�l���Z>P��<*�Š��V���t���K3�/f�1�T1ѷ���?4�l�-�w3jp��YN��!/c6ea�E�G��ۿe����f�W�;ӿf���`��ғR��܏�r�����Qr�:P8�
ٴ�HS�f�"�3���7���w�(A^͖���h����6�q�)N�~Jo���/�z�~�p0O�����l}�&ӑ���b�%%��>�����/l�{Z^��OWD��i���퐙#��L�2�&��^n0��1G�4їr��u eDX;�NA$��]I~�ɠ����I���0��U�� ����ix4p룰rp����b���-,�>�As9:y�o�����|s�3|�C�q�BK�k2�a �$�f��{g�9�"5��X��kO�PQ�����k���m�����-����Kq���ƈi���4���j�0N*���,\��g�]�HR�aIq��B�����tA��s��&^�c=��VAh�Õ��{F�����;�A[&�l�M@v[	�gaC��B��E��-�|�
徂"{1�\T�
�F�9�N�V)TA�h�M��������0�q�H�|�0���0z%��}�Ù
O�ެ��uG�����/D�t��Ԅ>�t�Lٻ� �'��&�.R#���[�_@\�^sDF�&5 D�,MPkgs���ʠ��a�]����Cb�b�^��O)m	]���-<�G�M�u�y��R"���zl���=�������_�q�[��� /yN�o��bU`�>�7Ǐ�-���� C�㔞��v�j�������l��	��w��l!>y�b�!�-7AvÅp.e��8J�Io�ܷ��~Vg4��]w>��o}��7���TNm�m�>�e}\A&�Gk�<�W?�KPaMR%;n��<��<��D(?/�ɐ2���.�Ɛ�3%ъ�f�o�a:���W��`��~����h���r��R�_JU4TS�Hf��J4?���U��*q޹Сj��gҳ.�Z��
��z�(DZ��V��UkBH�w�2���2��1�v/u�.bD�M�QZ�=S�*p>���/�yV؜���{��a��^\S�'~�?}+�c�Մ�/β��Xޙ����a҄��* ���5��i��z�	��}�0�<�4K���ّ���a����%.%�hڐ������.*���t��֠jUy+P�h�K�+�g�S�ٞ(4�x�����=S� ��_�Csޣ�3���́�
��o��'æA}3��m��jN�	W[�CD�}oeD��7��*����f�dt�a�#�/~�������X&W��W��0�f+���&��5�<�#�d�XfaH(P��1��Ň���C�l�`?���B�:!}�(�l�'jh�M�zQ��K�Gȵ8J�ZD�;_h^�&��Xa	�� ��n<e�<�}L��-J�Ƭ��/K��#HQ\ڴ�~x�'�Q+D�n����L��$+Y�{��1�/}!�B�+�}�=$��QU���z�s���CC�bf�B)К�_����z����y��B0h�u�_�G>pɃ���+`>O#	D�g������-Q��N~� 3��\�$�:#,i �����Fy���壜R�Y���tH!�*���ޏ)xKg�懿�R��5#���Tw�ce�>#wLM� �闄���*�0��;c�/���!XN��յ��n��� ��dM_����9Fz�\�Y� �S���) t���!m�����;z��4��:��|씮�VR�����_?����sk4E�i�L��v�i"R��%��V% ���lݲ[0���7��fzs:(�§�"��ǝP�E��%�:�`DF6}�IB�X^�([DG��i���4p_G °��l��c#��\p)`��+�)^����o EP-�������*X����</W�(r!p�����K����T|.P��=�>� r��MZt<!�T�[a�5��Wc']�z����k֓pKι�FU;��j�5���ޭ*Vt�
j�>�3�w�۴M�Qn:8���<#���Ic�bZ�C�C|A�#ee�����`��J�b���z!�P�Ԁ�L��2�
Q���-��j�#�p�Қ�>��/��ꍄ���;��Cw��9+��#�JTuP�W/l�u�
)7���ŧP�x��)�V�UѦK���~�%�� Ѓ�yǘ���ꂺ�t��s�ЛȘb��9zw4�
EzW��;�\ʄ������W4ٮ��MŴ����W`&�ڀ�W��\���e���ԃ��a���Ά����=�JӚ �HJD��@�����'�C��i֐l��1km��Oa�s@�hX箾$Ҙm�/�,��Gaj=<t���f��X�p�㖶��<i,�HX���Ȑ�4�v���%ŅvMMK��
���f2��Ȇ.%P&3����$�F]_�mcͲ��.H#z�"�8p�t�<�9b}2X�n�QѹN�LBóQ�2�B���~>�^�{��)gǉ�}O���N�;�~j`��e�����9����Y>�v��E�i��Q�I��A��{�����
��G��^
��˺h�LX�V3ޥպt�y4��G���'I����dRd{a�����آ?���4�������R�M����-A3�}�ҧ�]�ҍcZi�V�H�֦�５.��6O�P8��{J�[�-�US�!�I�U��v<�?�)D�3��=�HH�\`Ů
]��Q�Rw1�"w
�hL��i?��) �GU�Pן)@���,��s�>;E��Ri�"�dPi�H��<�ˋ�U;H��TH �b�8�r@�"�4��H�B���
T��
�RI_� ��*��:����~<��YY��3H�3JD�8]�B���z ٚ�m�D8�.SM�(�B⼍�(�-���D��^�R܎��#'zm�����˸�x.3�U[ZQą=������y��vԦ9�ӭ�v>��هI�������,�}�) �X�u���Ĭ�����"�pe	~6@`=��k3w���0b��t����N�����8T��nx.��
~��K\����b�=g�
���І!}��=����@����h���M\ZRd��@61J��[CZ����S�*��������V��p�%��5c^�Eė�Fr�F�8}]̹�F(k����>��\D�����$8.%�F�@�؉}M�oB�p�,Y��Ϛ�BAK��q�
���v��1/%l?�E�����v�;��X	�������n&���N�_B��ϹU�mt"�C���U-��_�ɑ�7�G�@�S��N���s�I���s
�{�&<���E�Ԇ� c� ޑ���Un�u�����ך�A*fQr���3/��ڪ�Y7� &��:5�(���G�q��g�t>q��D7���@��Sw����*.6'~>�h?�u�`WAJ��[ڤ���L�x��\���&7��.Y)[�d�H�zV����sjD�Il����#���d���v��#x���6��H��3�K=H��P(�ԅT<+��V�0��N�j}�ƶ6B�H$�ۊ�x�;7�z{�d��ZV�)T����
�oFy��`k��&F^'���8��� nG�<�d����~�E��ػ���3���j�{bn�;p��K��Q�n��Nmj��I���h���D��o��O㱳�r,��{ƧDB��8���cz�<XP�@���	����()��Y������4F;��P�fpO�A�f]�5�����Y� �i)�@��A���/5�_0�;�Ge�E-�2<��z3g�m%�x5�v�~L��7]N+4��$�raJ����U
b���U��U��H(j�^�[+��e�)����;�AP��CF��#���o2�q�A�����h���ʤ��wզ89�wR�G�
0����A����HH�����"!(�E�-�G��-֮5K���D�N�5�W{!z)��&ۑ�{�j�of~�r����,��f�U���4ɰ�#�+��c�9v��2fȚ?��#0a��p|���2������[E���b���c=j	�"�=�ʒE�v�̍R��������������;��j�N�T��i�ʈ͞�4��� �=I�-�X�q9�"ȶ
�a!��H�>n�m���q%x^2��זIw��	/)��xjrO�}!���9��O'��v1,b�w��X��k��sD��zI��k�����v��쮂�PL�8;=��x�!�#���A���Rk��T/Қ$���k��,K���� S�Pؗ{ m��[�u-�y�\�4Ld�w0J��t^B��v��S9��b3��H8=y,��{z��N��q��`-@)7��è4{_�� �:W���U}WCU#U���$)3�Z<x{�B�1j?O�2?��'q<��㍻�:vP�*�*���`��b�3"W6b����k>���#K���cQգ*F�̄�jk��s�r��(_����Y��Jδ�g��;�'R���{�C�
1���x�K��˧�R�r&�t��2�P���P����!EQ)1�������y�F(�o���s�TU���Fu�	8a�D���Ȩɮ�u���	�t��Sy�w8<&�8Z���9,eH1�	��G�O��� �'J��P�E�D�Y�Ԍ}�8"��=�*����P�x@���DX��(��6+(k�h��	��i�]�Dþ�,�6�Hp��.����=D�:;W��1��b�H���f����J�uS9�(��5�Px��J9��x>�:	��mǐ-	�bе��E�M�*O/�L�BZ��	���XOt[������v��T�Z�������Ϳ��KZuK�.�y/��Z=j�;�������oޢr�G����uN���OO}F��/�g��U�����C�i�+��� 8�o�Wݐ���:b���\*�e����>����%����k��*���u�L��fd�]�:�Z��2���Z��5�E�����N��:K÷`����ﰢ�nv�05(r��*,Gv�-���Y�z����7P���o\T;t�JL��W�:�|}�s�<�Zg�/X�{���*-�w���Ԕr�fpBŰ"�p0$#?4�w�%c$Ǻ�lKb��J>����0rj�c�*[c��X{���̤BQQѓ���A��X)���tN[���9�?�DP����9����H�oVP8! ���ª�*���nq"��A�a��� ��/�[�DP��ViUa��j��S5�D2}�q����a�f(]��;&'Y��\v��hs��ݩ_ �3P��Y'^�␖>'3�)�0��#p�T����;-���W�7�^?�@B��el��W7 �1%
t����'�����f4:��j)��lF�m۷���~zk�>1%V j�0�(~��9W݉�t�3��Zc���u��ijt���AŮ��'��|ek��\�sݖ��i#WnWP�A�P�;{�4ՓVq^�6��i����<�a`��P��P�w�$=��(�j���mCu\�_�S�	�������[{/f|��k^�:L��аƢjͱV��R���@悁R�\�-�0_�/���/0�#�R���x��Y�/����E��z��8��ylD���6U�D�X��+��«v1@��!����[�1L��r��郬�L��s��GBW���^������_l.U@އ��8�lI�NZae���]��E*�����F�����ʹ�?����!!Q:8��?����N���=�a?��
�W� �ە��T#Ζj�aX��W6e�K��bu������pv;�2:xu��497UѸ�b���twLp��v^�����yG�o�$�Ջkș.�Bں��	���03��4�$І&��U�6�Z�u �a^>�R����*ݒ�x.G��]~	�Ǭldt��ް���ƈ��"_F]ʄ����Af.�a!V��̌0=o�9�A�څ��p	����w���46�$or�.+$/L�ڬT�Ґm
\���v5<���2�V���|��A��=4�v�h��U�$'y�e���`�@� ��L���j/ಎgr�鯙�;� v�xD�LuqVc�Sj*�P�x����p���|�>5W���D�b������(�Vq��<_9�C�)i�3���z����Ɂ_gQ�;!w4s��/�h�&&�2�XZ6Z�f����s���.#�!�����Yi�ŧ�S9|�s��/���h����+�%x���۶j�>� �+���i���#;���C�|�&v;r]�|�'��Z�����_ԖN���]M��[���y��kU���<�=�!0��Xn�ȏd�5m��Y ����s����A�9�*J���]��L'�CYR����:I@zĦ����l�$�7(���J�j{��+�͚�������RދN�t؛�
H�+a�QY�ɹ�q�����+h"�0�zHS9[���A�v��_x�U��Fr�B��l�����+s�&]�.4�����M@|u�)�Y޸�~�hb�������M��a֧C�
^2� ��F���Iu�x��:l�7k�j挰���D��l���{U�%kN�N�g/�zw� o�ʩDڐRQQـ��Q4��EzΊ�Ψr@(-�Ģ�9�噥Mv��:��0w���E&��Q�u) ���Q�d��=��%�P��>�O 2�#�́9��$7�u�c71s�II��Q�btj���o}�ոM�%>GG�5��S{!/z�z�c�KJ@��]�[������u	|��_~e๬��Һ�Е��t&��_!6�\�g��H�A��o�dFD}@��GrvZ#^�d/�� ��sƯ�>BP=��B)A����!,BI@�|Ia}��x�$J�]b!v���m~.��(�_����.)�TΦ~�l�#%�W�ʞ�>�hQtT��-�p�i׈�g��Q���� ���01\{Ŀ�+�gj����ƤU~2�S��vu�_���!h>�����Y>j����ԝ?���.��O��,����(c@C]�F�u�;v�����2�m��p@M���F^<�ƴ��(;7��T�ˬ��������,,b}T��'�;Qg]�PO6w���^R��>�����|�$��Sk5��~Æ��硋��D+b����[ 4�IQ
������}]cf�o��<@!0���>×�7���A�w�aym�d�?��,�H��8]2�ݨ�'�Nu�Ŗp�D�_<�L/�?����.�d�g�_^���v���g�"�m������a����}��N��`)����=�(�dL�ȪM�p��ѥ0��\*+�gߍl�wn���p��wE�/�$���M=6�k�E�Kb@]x0��}#\<y>��Ł�i�x�-�)���{�0V0*��W|f=�ۂ07��L�H�(!��Z&��`g�TN��[����W�1�ug	8q�@�H/X%�S�	���C��u��Ȣ��+���A
�+����)ke����Xk�2��v��!��ý�E���a4|


Vk/ܙ��Bq�=���ڒ/*�r6J��S�_�`����.�����:�"?.P�QY@�vq�Dz3e���S6�'����<r.���V7�3 ����Kl^\�>�F����f����G�]�}d X;1~"��t�/�R8~�sa�&�����e�\n5���J���.a��?O27
j�D���_���g`adP�͖x�z,ǀ���RW��Ô�r�,��2a���k���6"����F�6�X�r�P����ɓ����+%��� 7�5��q_�'^��$�+���-��%���?z�1�Ky^rmHُ�=O7Lc����Ճtg�}½J4%��F��-ԋ@�ׂ�-F�.	���~�Z*Z[~)EYa���_}��)�.*��q����Y�n�0;�o;�%�����,PsZ���C�1:������X�8�$���:7.C_}��AHx-�>˺�
��,�
�}�����&�hB%�wi���p;	UOI��� ^�����?5Gc���&��]����n+z�����hL�ٻ�r.(.dޯ�n��0�Y�{�&]�l���q�윌\�?"�e��-�*�Z�9�BZ�'Z��xF��ݵ�r˙ʚ+�9)r�9�%kWC W��ǐ���[p����d��-�"�X�j��?pPW��C^y��B�x�����2�s4������~JzhB�ޙ��?�1�ݹP�*��*�`�yԚ��|�~l��5E#�֛hq�.y�e���$t�@����j �"@�9e��vk��#4�EX]Ͷ�6�Wį�#��!����j��x\��v�3�2d�N�qʜ(ѻ����n���}_ZMy��Ks�� �h�����BN����P+s�,t��JΟM�xb�u�д���i���3C�+so���Sğ+����LM�CG2+�e�����j3��j`1A5��$���v�iXSl�I�rmR�t�&6S3!�ilu�N�^�E���Y������,�멗�i��{NtW�f�1a^?0�%F�_�K�Q��j�$�6C�w�=���F g��m�>H�^�����Pcp!Խ�lV�0΢�yXv��ET;��댳�	�֖�#�1�wB2A���0�?'���m���ǥ	%B���)Z{D^�yo1�ϲp����	;� J��T��䓐ė�T֟�,ޯf����.}�;�S�49����_�\%�\����7,އ����W��08P���Ը����pms<qvO�����:F�| ��y��e?��敍��ǔ> �93��o��������;�=���o.'6ӽ���<�o����J�;9��)>���-B�\�JlY6�e�/8���ߐ�"O�\/�6SS��K����c���t�	��Ņ�ZLf�&"@�e6NA,ݰ�a�(qG2!?�P�O�"o'�r�~	1�R-of��u���⏜�0�ZX����\tM��-:*^H�A.�P 5��/Y`~[()^���4�s��m��#R;L�DX�;y��k.��M����f�D��L�yR:�GRJ�U���~��14|�wG�Ұ�㞫�^��Be��9�����H>FNl6��u��?T������8�V�+^�)iI�5��}Ͻ�UW���P���m�`�z*6'̉�v#�a�\�5cc٣�Z��mu_�p����1�t_��Ћ��r/Z��j���l�=,��teXC#�����5�k< �m�[ ���r�������}#���� =߾|2Z�P|Gp���Xsk�Oa5§�y��u��H��4�0�<�ܑ��5a�x[|,7nv�@�Irn��# ����z^��6�[A�dT�߀(�G�Z�$��~N ��O�L໻Myx]�H��U���k�
�/LP������jn�3I����0��`.�*U�	�A]5b���NKhQA��P��� 1l�EQ|$Ru���)h	���TF���*�(��~V!i�
-�%��l�%���>q�L�������³'����Ch�.`A�tl1����`���d_�_]Y`�XB�������� φ��:����W��{���#C�=���oㅕ�N'��_L�Ȁ�i�)j����ԇ��5Ia�"s@�������[��b0�S��\��bM�R"��:�[F��/���%��'�`x�5� �;T"�lrX5Q���9���*���\ԙ�0�T%D�<_��M���Qm]Ҧ��:m��!�^�қ�6�Es*��@��H��=5�th�I1�f�R�dZ�ܚ����$Ad.+f�������.*��.[�����S�������$��D2�[Z�� �`�����S�������X�^�������D%�1H,�클�|u����8�������n~&%��%F�sJ����Z@EB�"~�.�ꁙؘ�>�@���P�)�_�Y�:6��Hd��{�����i������E�sM&�����q��`��	��
��?�I�Kwѵ���3JZ�=.|1c��c�펇O'�A�+�*�G;��̻C����(1im'�8s��0��nh�{3{m���4���1�/i-A��|���I��@�k6HB�s�vj�S���S���L�r�^��� �TO���+��?��`|Ra���0sv�C����`�ʴ�ۉC��a���3���@���kj���ḌQ�vs��u��o����F��Wh�A�����;�l|���?{l龿�ph����7Q# �m���PS^�f��3�Ud�c=��ON`v%����8X|0��w�m�|C��Z�0Ԯt^�|�K>��?�ۯ��FK��VZd[s)��<%�4�h��yWV�}s�y�1=��̍^I:�#�i>���IlAj4?�43���	�n#2�`!1MgдT0�+'�+]�Z����:�����p�X��C��[Zi�oXj�W��VnW�}�ykk�ע9��zp_��Ԥ�,e�m�4+a�P������s7K�2ޕ����e�3 �x�=����E*��5T�i`��5�?�����QTm���t���Z��t��*�m�Z����aB"Ү�ם�b���hlp^��F��z]�%h�p�y�G>/]��;�U�:��
"�oX��#۲U��"�B�Qw�ւ�;�^k D�Wm|-�`�񮭣&n�Fx$xl]7�^�Ԕy�5��(=�&T��HZ+���M�4�3n��@���d�r��}`��ˡ�C�����@�'�àϻ?(ip��ҙb�"#�z>�%ЬuKB�H�c4�s{�0����� 8t���Y�QO��U.#��5+�
Hc2�� �V�7�K�ER@�;����v�u�=|�����-�\��ط��W�.2�dP�_�/�zO� ��L�w�a���g����f���&���L�
B��w�-u鶆s���Pxi�T9��
ڈ����
,Ћ�� 0R�Z�:�L�s�Du�`m3A�=�u����o�߇�p�F��צּk���)����� 4�k�?gc$THST[��	�����I��z��Gm�!+�����l��;�Xق[��@�#���.HZ˝��6�m�\�l�y��~ߚ�1���Py��"��-��.���C�͑&�Q�mW��'i�ѦmId�j�V�>��I�:�
J)�� [P��/�d���h�&���a1d~����r�hצ���^=
���ca@X�a�g�Y������.�"$�	��+I8�z̍�Y���NS8��Z�o��r�cA�;��
| �PV*�R%%�Y���T^2�K�����ùa�&u|�I!2��J��C�تc�ի~��L���=�x(Xюݢ5�eX���Υ�L�N�6��&�&h:���?�ɤ_Ƶ0:�yXD��R%f��9.��n��ޭ�_���U��T�+Wi�C/�._~y���z-�gm�X��g�y�p��E4�D���(Zw�����s˲u��BްgJ1�̬��;fVJN.�#�L�a����_<���t�����0��3'��(�=���e�`��M��M�Pv�̅ ��#JE��8� xc�q���#2�s-B��|�AsJu`\%?oe-����>Ӿ�[o���'o�HL�h��jO�/�g:Q�#�mp*��_�E��r&kx�+��7�^�T�����N���eKF�4�Z5�'�Z�05�e�J�]1sʃL���c$�s��.�Ҙu?�ܫ�a5���A 	{�D���G-e�(,(j��7�e,��"�A� *�J�y�"��d-��d���])5�i� �E&���%v�1��^�?ꕲ��Z�6�b���i8A��Y�C�_eփ�	�$3�{e���+&��'��y�$���̊:���>�@�e��#-�����e��36����f����&��0�UFlv�HN�� c>��m<8�ʚ���4]qĿ�@1;Kd+�~b�
�"���)B[jvQu�&,�������gJ�����kDp�б��Se�ѵd�x����}:�K/3_�]�B����)|���Y�A$���v�����m�qǁ$@^���	���d._FB(q&��"�,�#-�}pγim˯Yչ����+�2M���Gb��l��:�|��0���do����M�p�)B>�����(��	�����R�M��[������xC�`����\.{0�K�Ț�O����`�
6^`\?��\%����hW�8oxj�:خ!HB�ּ��ƍ���Kïs�z��L������/��"_q������ʍ
�@r�a�M�7��b׃�T��9��!���0b�~�іn�%s�*�q~����/F�\�b5���O�(h� ����^��XYu�p��T�\ؽ����L����rrV�(xF���J8py���Ƌ����w kr��g�\{�?�<�2��S�r���>9�
���@Z���(.�z��A�x���V���ly$�#�f���nSV�'�ҫ
�_�XHN�ElB�����	�������Lٿ+���I�FjL[�����7������ř���B�p��>*5�B�U�m@��c�}}�t{�'0�(�4���f��>��5IR�!:�+��"ĵk��qK�qq<*K�G�����A�BΣ%u�at�nJI<'���>��"��]�7q��"I�b> ">V9�}E=�\��n�>'X�Ż��Hs<��XXpT��*���cSk	;%����u�++��$�^��� ���R��G~�(��XTQ���Z�C����F�����3oM-�j��9uR.t(���LfĆ���ɦ�~�Nx��zZ����%�t\rj�}�3�ijvwC���mJY^��FiQ^q=��[T�~".���J�Y�LB_o�w �Z�G[�׶��k��+n��Y���]b��s7���?9=\C��:���D4(����ͤrUF�#$�
Y���2fU�.��ᴊ]�23���og�.In�W�a���μY�
�GQ��0.H����w��Uy<p����tW��^�PH�lꀩ�����+�E%��r�u��l����q_��p�q�]-~I��P��)�|ft�O,B�v-|�Sy���"�h��j0�֋$�)� 	F�=���Х��=��d��5\��]���K���H}P��l�;1��Y��˖��v�(���eJ'u�)A���C#*oSh�s�ȚJ��e���E<p6;���DIh�"D:AaˏWU4�.pl��a�8����Z|�Q~��Y�,�%s*'4+�|�K��x}�G��O�Z�U�)%�݂.�$ͩ����1�����𷛸s?���Oɩ@��NWŽNK!([��џT�J�G��ik�҃,��;Uz���崝�2=�dӯ��T2�����N�;����$��϶v�`�2)���^V��x�[2��m`W5�7����4S�c�� ~�*b�wJaX�D�t��#s�>d�A
����dQn�R��V�_�	�|Ϥ�B@� b� N�L^&�"�'>҉�7�s��!ߚu{�x(�&��+i�X�Xβ���*�o��	�0�S�;xfo ��%[�;�'��Iro9��JfȂ���%%*ܷ����r�*p�aπ��Z gc�"ep��<^���>�Y�o��t�؝�A2��ə�b�5xs�.����D�(�w��6����V�o��{P�zpq�\���'�@�YxT�����Af�Pv�1�u_�8H��џ�׮EZ%6cI��jV[j9ct'�U��`V1�
2W�J�M�Cv��]�,3@ʦhU����JyAU��q�A�y�@��X-S���
u��/)���$�[��n�۾W�)-�&��Q�hUeF\l;��I���]��D���yUxz�ʼ���I>���(�o�T�v��J�1{�f|�˅�\�BJj`_����?fA��-��Y4�Sپ��o�jF������	��DJSg�i���p@��W,1K�<�n�x,�;]�����a���xK�A���q�����o�I*�Ζ�K���ty�����I�d�cD~������MRVd�����'�OĂʵG9Tu��:���|?�i��,���t����D�	��8���/*4\J�DT���ya,A�����@H�fw�WB( �'#Ljnrt���ɓ60C=}Cc5�R�|Q����?�{� h���<�^���y-%VS��J��St��uqp�j��h��dE�:/��tB���*pC�,v#���3�g]��'��Y�%��P'�H��1L�V�ϴރ�³�=+
����`�N�m�k����4�p1go��<�Y�]�~�-\�>ؼ�z�����X���/%]Qմ�t:��<�[Q���a5VG��"S�+ѧ,�6��R���by��ø�����^�W4�r!���{ }����HxJ���m�E�V}"��?*$����=�I����۝_E�Ƭ�T��Ρ�ߍh.������m[n�q������KZ8"��#���"
�&�02�$��.�/Ъ�rk��R��� �(	s< %DCN��]q^97Z]�����x�?��ֶL����~�x�ؖ[���Wz��u�v�N�bw�W�(�݄Ǳ!֜���^��Qo�}��߼��ܿ����T���o�)�y�eU6����IǷe���N�Ƀk9"v�W��ЁK�7wг�n9Z'=q�͵�
��ef�i l���-������$���ٍ��8b �&����;�����b�
h��ǲ�h�m�P��ƃ]����"W2j{�X0��[w�D����5�W��>�jrbTVӤD���� �q�ekk_��u<���3o�4���k����'�� ��m�W�i�v��<��xȿ�:2\ؿRc� �=�^�^f�>ؗQ�V���J�3�>�4�U8�#eX�fK���^)nPDhB�o�) ���1���t7���1���-�L��w������}y�eu�~���z�ׅ� D�¡:4�p0�P���]��0���չ�P`��ig�r�U>��LV��䪷��nui��}3II��P$Q�w�.���z�*p}_���z�dg����-ӨТ�"C����'�/������A�&늉��1�AX���K.=�I�}��zb$7FQ}��ՌNܤ/��j]\��b��d��̷T�1�;]�WG�Г�z�a�-@��t��y�Ce���:���<s5qq|r2<o�!�ӟ�`��u����ju������>�}'gH�p�m�~-'Cm~��uLƗӪHb�o8\"%�X��N݇ ��Y�x���z��K�3�X����կ����B!����q��HR�m��{�`�\����U���[ܩ���.�P:k��iŃ������l�C���ԗ5�|���|��\�Cp������ʢ���03'�<�iu�g0gvZ�҆����l���N�Ұ��:sj��@��&�nY�'�����tqb�T:�&iAdh�u,��o��&u
_��D�A���XŞ��6e�+o�F~���&�.�O�[�j���n���-=����`�VE���e9g�o 414 �S�G%l�/rK��nP�4��z�7�"���ٱ���݉ÀϾ����w�)S��ף�9O�=��!ȫ@N�d�PЁ�҄�% K5�<>����v4�R��J��]���Y;�v�y<�*�}��.���R6�\"�#)���
c�Q}"��?��������'�@*XP.��k��Pp�J�3@ރ����T÷%���}�oa�.`���>*���h��xwf�m��������ꎋE�� ���I-YDq�.Y�~�h��ٞ�(yAEp��Ĺ@�bUIi\�aC�Q�F�%�>�_E번ji���<�0���$�E��F�wG�6WAg��oc��"��2٠��,3t*h"�� >����!��b˂�'J���?`H��..{A4/{�%>���ښɓ�Ty����(<,����+-��>ߔ�x�Jy�G��fɂ�0��4��=�G�2�n���d�js���MX�E>�����r�};��IA���z�$�,��@y���F�GVɢ��3�8�T�3��s����/�S�r�[�G=9@k[e�=��O0�P#(f`�*�P�T���،y@��(p�	�Y�{��������w��&h÷���Ԟ��7xIM�Y&�Dh7W�i��w C����e�-�<��:O�׃�Ͷ�4�n��"��ycpxJZG��q�8S�0�J���">���Aڟ�f��	K[Δ��.��ٰ�7��ǒJ�h�j��|�%ɕ�Pٌd��W����9:��(HWi���/�1��YB
�,Gɧ�w��Ϋ	��w2r�M;��9L�i/�dH�7Z�W_Gr�n���.LA�.cߠ�^���7�~GjuIʮ�Mzq���W4@Rp N� g���Y�fU?�P�1Rp����(o�����@q���<:�G���H�ղ�D����I�6絳���|�f�s2�{�Հ��yΚ�e��	��/��U�Ǻ�K�ˇ��E�ͱ�*zg��i����ռCA��q���R7#��K��} x����]l��em�Qń��ŝ�y���|�H4���&������F��8�M��^vg���
đ����$�Ao%@,�b<�Մ׬n���ӏ�� ?Wr�����4:�%<xgC��ֻ9�_b<b�:]��N�J��6wXQE��8����ե;�gV�n��MXX��|��;B`"�R�6ᮘ�Q�١�,��`B�ҶqT51�ݎ�9^�11͑���➳������la���f�-_4��Z�O�rb�l�v�'{����R�K�¯ʯ~�UCH��i��n%��u���-nz�]�x������S#3��p�[�d~���@�s�^���p��������=��}KVx՗��)�D���-X�7��.렡ƺ%�Lj�!� �c ����]e(
����j99��sJSQ	��3�T@[���]�5������=��)�c�XZ����R�V ȅ�C���Aw���z�n?�#�$�jf�dq?A7�j�+M{��K�3s�*��#__��D����u�dxӭd�t�`�62j����-{����C�U�Q�P88�ݏ��Xt_)-|�&ǖR��f�m�:([�k�,{��N�u����)ۘ����Kv���®)l,R�BZE��,�J��I�_]���Y��ߡ�����M��o=��_�5���ڮ3Z$L�� _�a}�?,�t��C�]8�c�h�,�MFŏ#%��[Y�P��3��<��K؏ӇWɓ��s�Y��VVA�3����+(ښ�-U�^��������A}�-�g�mړf����_��m���P�3vEu�;d���a��>1e7��#���Nz�59���3����{e���,����D����e����C�u�n�ҭ����~���W���`G�oS��.���+|�������eC�:���p�˷Ñ�>9�h�|KӅ�v}ts���oT��4k��`<�,"�nVT��0:e���k�O��.�هA�c|?��=�'���&L���g��1x_�*�����H���@^�Ꮽ����}�|���T�i7�un}][D�	����s�lb+C�8�~n����Jţ��Ο���e��~���>�6�ئ��C`��3s1"�=׀H��׷qj��lu
o�m�6p$ ���rx�K�.���S"'"�WW`'�q�P �}��u����qP#��;���3�	\�{ם��]�#t{j�sV�E���*C?$x��߀��Q~�,�IȺ���ڹ[�U��̥�>�!y<%}�MkT#�@$�=3�l^����=�n"]!ˆ=���-�C;s�6� ��"��?�A��X��-<kՒ��D%��{+�K�g��}4�D�v���VE�,�ki=������K�!����5�z_�T���)�L#�2�9�E�i)����EɁ<eX��"��=s����)	����ޙ�:@�G!s �pg\�!�O�.�rT���r��;�M����w_w�Ӣ�@���,b�$r�f��^5���6�ɒ����] wK��N������9P��ޒ�!�ع��R�V��V�G�8Hq�i�X������뺮k�IF�ʚ�d������>|�E[��uP-�_�Q-���)Lk~�5��;X���8�����pt��sXr"�.k^3�Nw�K�zyE���E���� nP�Nz��^��F��x�5��P�u�!�o
�D����cQ$,Q��ڐ8�鑨mR���P���;���v��Ź��-X��$��0�K�|�C��Y�EƁ77?Ȉԣ��ȱ�B'��8��4�@d��"RN#ݥ�ѓ��D�[�J�W�S������Fޑ"�44���jzOQ4�>
���g;�[��/���R훒#���̟��1�zmt<$)P�g��r��⍶:�7�f�Aɩ��>��A �êL�wNS���3Y�S����t�y=d�i�>w�X�M��6�>Z��Fn2R
�Rl����C�h�y��-�:�JrI�	��qIl$FE�#Z~�յSG ��-e���W
��84��`�u`>:�kZ������U�r��@���
qǕ|+��� y�V�w��G�$�����bY�*>4�Gt �Ú!�ދ�Қ� u!� �4g<Sܪ���3�#��RJ�L��,�ƻ��n���mi?��ٝM=}eS_i)��}iD��vkJJ�7N�aUY�4��f���Lx|@2�vˁo�pB�Z�P詥g�;,Q�mfd��o��E�F�A�G��#J'3��P��& ����$$=&�k�Y�)�gh�'�y�b:�2�X�LZ/���JHx���!/��2\䨹�7Û�ߣ���'js�ҳ��@m�_1���.�w���*:l?	jD��W�_�l�a$)�;�T��H�3.|��lh��I�����V�����*�����5rX2^�2���W��&sU�t��8�?��RHKA�V�H��c�u�fLX��0 �����j�&��-Կ��aE����/U�R�@��G�f>٨'���'�XP��HDwW�.��w��"�e��P~Dʿ���1Gw9%눉�����Y�,��Av��SU�C2I�7�h}��3Z��6������9���M8�����I%$��D~��`Ζ���-��a��6�;kD�[e�7��t��'�yQ8�����px��ҺY�-�>!#2dȀu T<Jx�?��|�c>�|�-������t�/6�T�v{�����^���C�/u[��P /4�^��+����<��Ȟ^��5B�����h��"�ӰEGt�A.�E��1�kҾ��I���#̕ ����� �e]�c
���$ji�!
G�}tZ��{����LxT���0��R�Ġ��C�07��5�SK�5!��Ǟ�=y3E�Zx��e`��G���/gaV:{�p���S�7�k�bA�.��5L��Xa�S_E��m��+bO
rp����3ܿ4��7���Ι��L�c�̽_c��PA�w�p{W1��*��K�3�Xƈ7@ V"�l�e�ɴ�����c�=�X~Z�7Jx)�uˁ8�5�j�Q��4J7l=�$���G��QVÞZU��]�<������T��y���wXPW��n}K^M���dl<4�����Ƀ�qK2��(N�d 8:���ge��"�4rF�9ɰ�����E/��h�q�y��`_���bcu����N<z!{4�� �yU���N �f���-�V�[���?��o��3��G��*x�Q�c��_kA���\?��vʏǇ;zW��ȿ��(�$X�����=��h
�b�c	 �[��o>Y�����y�zuT�q�����F�U�[�U�on+�̺�����j���Z⟰��7��wNI'��������P���L��įPR�7�%�,�az"zG�j�u��M(9BQ�s���ë;9�\ ��.��3X��2���Z=dN�]��-�I�!z��<�s�|�����T�ԖS_�#�p��� ��`��A�1
�OPSղdh��Sٸ���F��>��"L���x g3�es�� �����h��Y����>7b����mo5�-n��r��V��M&F�����^O��/:�l%yI9w��Zf��1L�]�*�-N�,	��P�v�Ъ{y���}+�3il�(��ιg?UhC��ٟ%&�m�����͸������+��񕜕��K�T� y%�g���9�	�U@�/)ͺ��	�
��^�%����t�"l�M,�`[������%�)�i�x���N	�z���?(����o|� 9��U;�x�W�������>�e���<Ǆ�f{�p�c,���������稹a$m�x�]���|��$��3��>���nRI�@N�Ta��}ʥ��s����Z��Bo�-��}w�S��d!D�� /林�B��~`h � ]C��d:���ʟD�W�ݷ��M0s���)Nڢz8}bBx�"1�\8�E��7����7��6x>/�^����Dt���!^~�qr�o�L����;I�)i�=�8��9	��Ĉ���D���L�تPMa�$���cj8��3������	���P�ߝ�k�v�˱E�t/��!�i�G�Z�ikO�{��CJ�~/e~���ɑ;/x���E����`*�u$W�3������n!7��B_q�13N�^��E�h)n�u���<C$4B�-x���'�����UJq�O=�º���픔X���'�j�1m�:�!� ؁�E�k�MRħx)�11��Ͷ2M"�p��Y<)��"S����ky�tjw���5��<f8�-X����<����NnJg
!O(=9އ�]��_�e�&��!ѕn�뺫��01A��e:;��j��b�?z֍���6hS�@b���\����:Z �ɘ�ldG1$S;���E	oCgLn���R�y�B�ƺ�q�>j�t�R(Lf�\�/� ub③�gж5W�|���@��~����0B7�M��u���	|��R%�h�f����Љ�!��c�d� �B
�<�Y������+ű�r	�������~uh�\ᇻ&�A2��1��"%����xZ������vC.}�d-;��M_b�j(�����Ε���"�Q���.��RRF�� $�h:��#�c-F}�>�6ף2��SG~VlD[���〞�}ʜ,E��~��p�Ѝ��_�n�/��C�|VY�9e��Ѩ�L��40�V6k�������n���^�O��%B/�������G��q^$�{Be�P�G�N�7�I2Nrd�
��y��m	^���d�T0�3潔����"���E6C��<���`��>�+����dZ��Z�����9�iz�,mY���ēn�EL��q�\B�b��I�WS<���S,�7�m��+Vu�o�-�y�}�v�����*S�T:f���>�خ=1ʨ.��:!o9�7/��X�y�T��1gĻk3ފ��0�T������tt��j����.\Y��£3g���x��@�̅RV�vP����.�ARI�˃�e�tr����#���\�!�
P6��E;ʋ�z�'�S!��/B��oZ�omI6]���-�	�|�t,vc�+�_4��,l6i��Q��]�wu�nr�p74�5����lf��3���qC�(���ͣ=�����Z$�9 ���5,��$2M�5�k_e$P��a������:k��WzFC�����6���2[��4a��c�� �P-f5��#�he ��j&)���ȟ��"$��ӈ��h@3E��v�� ;�ˁ�Z ��ᴾL5ѭ/���BB\�xo{����ܗ������>S|��4nA�e�u0�Id��mk��6=l_8�[$	�Q�Z`��Wj����u�?�I)�����Lx�O]��}�Z6�;�^d�O��"��{���Q��
1ZK�/�:kdFS�V���7Α#A/-���?�Nω����Np�Y�//eךLS�&G|�tR/�X���+孴J<Y�) V����R�]~H�$��|p�6<*8$e����ě���?����+�ՋǇh�)��G�WU�����{1%�* �/#ʑ������;n4$����B���*R�=B
�7e[$ED뺖A��M0�SM�y[�`Ŕv���������V�6CZ���B��^��ޝ=����}��-���������Da���W��%6��6�"=����|6+��ܢ!c����N���BHt��=���ti|��S�	����5F�_2��",��
�� ��;{����GK@r&�X�Lp�7[4|+�����/l��3
�Ba?��d����d�7���+�T���05���>�) ��h�W�w�iW[��x�����DeE���'�y����^��!|��g#�tk�I�$ ���(���"�� ���@�\��� ~�.+]�C<d�FQ/f��y��9�rm;��� |���6�̠��@�q�BV�0F;|�c�A̱@QE
��"A�~\��irh������QZ����?_o(����;���w0��w:��*U�jA�����~k��V}`�נ�G��Ŷ�����s$��M4���/�cX�b|��ZH"4pb������8�|�q�Ac�z� �į��}pg��w�=`'��]tu���%�A���lԹ�&��Ȍ���Ҏ�f����&g�8O�(#3���7�v������a�֋L�[O轠�"��@�3_�^�k���&�'��e�g����d����"��;�Qͮ9�GW#E��$.�7�����Ix�~_-�؞���#�UIg�`䥂CMͮ�)��ď��qq$]kXC=S�N�P����;_�4��,�wAv@Δ���4#���k��N�
<�AP���R*�HR���P��1MRINZ_Z5m�M[đ@bwu��O�?=5{���x��S�N���A�fXei�ܢ�$_����t��'�v���5k�V<i� Ʈ�e�����8Z�V)�t�%0���(FoE`y���$y�u�/���f�qj�?)G��fS'�,
��޺%�2{��mK�D�j����j���O��<��	Φ%�38W��o��ۇ���u�b�R���������Y'�X�L'B��~)s=ٻZ�m�;�[u�X8��P���~��d.�m����P�"�b�Ǫz�_ "|�  DM+ Qy��1���ۏ��R����Q�0�,���C���A�b|}_�#^�e�y�c�i�e��t�����߸���읂���>K��bǼ�Mzxt�(��l?�Y���_<Q�p�aP�Rp*�s�RLR粶�� ��b�����C�y�����C���\?�I���t�k/����vJ޳wF����L��+�ee���@���idt2ҟ��9G���ve{yB]ڮ�6�$����א+����b�C���OG������C�qv=��m=�_�8����~�/)��_%JS����y��I�D�T�]�Tv)���u�xsB������4��uP��_��d�&X�}�c���x:c�L�p�j�Lm�}?pixQ����;2��?f���p9T߸�4&G\/�vE\Ԡ ���Z1� ���~ɪ��ݦ�X�لSpAՉV��/B�r��L�����N�����5W�u��>��r�5w�(���&!׳��ќt�߂Fq�b~����Lʪ�v(���J ��لG*y���#�&TlӬ
�ĸ�d����Ѫ�X��g�Gl�Y^2���s���V�j�'�v�w�ꢦ�m�f�BN�(�D�Wyf����	�r�/8��&���5J�������g��pt���w,Jt�����d��#�m{!�[r/�����Zi$��i��R�`���{�j�O*E�A��>a���W�>�QT�*)ܴl"���kkP7�ǯv%�	Rp��2'��
����K͐%��ݤD�$�W���8���Q��Y
���N)@��M��U����ţ���$�pu�C�)F��|6j�*F ��A�S ��,���6�vX�w��	��+zP�W�����Q7�G�!Y�2�D��$V�g�=���As���Sa���L�H���ʽl����zFl����
'�¬����(�T�]r\(JCHN�M�V�Fו�c�	0E\�	�
��&�\��Ԝ�UQ*��-ư	 �.yCJȗ�\XX�K�]���@����K칣^�y�xA��Q�C�@�q��b�-u+��6�ٮ�����~�q�&�~r�e�ʓ֔	��	�j�,��T�29�߯[����'��o����I�z8K�}$����e��w�g�����d;�:%�bt��1��o�\���Ϗu!c��>�A&�OS���O�u�Lk�nড3P1˃��Z� ��h�٧q� r X���p{�5�wy���"������Y5iK���]�So���|@�SZ�ݩD��J���<l'�d5�;BϾ`.��O��קP�]��B�%I����l��j�9<R9� J0�|q�	�}#?�ĉ�Գ}�mY��J�(?ڙ#cP���7���2)�/�|;�̨�~�*��p��ʨ���o��'Ƣt���a�֍�x_���}�?��'Y�����"x8�q}X�W(L�5�a��:�ok߉P_�cHdx�n�.}�;	���b��ª��X�ӿ�$W��{�fk�C�����᪾#���-�HR f����x�_m�����:��1Y<*��"�������X��0��L I��3��~���C�mȼ�ƐJ�xp�]��� ��J@s�"��-��� U0x�yɤ,N���(��xl�1VՊԳ��O��@�O!a���H�����}�A��}��ѧa��Yu�{�מ���	���VA*��62#�m���2�#�^�0&8�ɵA@�8h���~�_6��}/xe�Z�d����ʷ�m:4�㧱�����"�S�:�R��;��
�
�o�%��!Q�GQ�h/����*;jB�v��v�F��+_]Ŷ�����Y�������o�'�6���=��h��F.O�|�`��^�υ,���h��
|�_��c�en���I�i���6o(X1P/����N����L�Wa0��J(�0����J��pھ��G��h�|CO?�ޡ�j��t��+�I�J�.n~ԷC�	�d���$�����R4Q�|�5_���="���J���昗��QX��ݫ_���4� ��0v�^b"��_�;�G��ˆ���Бu�d*6"<�ym��[F4�Yw i2]��ɸ8Mse�y3��h��7�D9���i�;�i�����t^8�P�e�:��w���-�1�Y���ɥہ8B�<?dݿ5�����?ށD��ci3�b&�1>��v~R5lҲ�K�4�{���w���P�^�l�R�����rșNc�PoVS�Z%G5RG5`_�s�,�:��F(R���*�������$Ӭ>��<� ��L`�ʈ��	Zp���}wϛ1Ǹ��ηy�p����y#�j��d���4{��m�y�����a��i��H�xˉdy(�kV��Ĝ��7{����~ ��}�S�{�*.�0���b����];> �A��NB�8��뻖C�(?��q����K��0#`��ϵG{d�:�����G��$��?�P8�iѺę��DrX(���3�SR�'�4S9u_I�!W�!���c^$Tc��W���������s_�t�g�J��jzb@*���	�'yࡻ~����#!jJ<95y���4�� �i�_�8�������$�xN���ZqfLk�����\No��j'�����ϼ~�W	��9OH���-�j\�Q|�+���r?�N)��|�����3�T#�Zu����c	��1�<I09*����:�gIơ髄�؏<�EQ����3T9���u�Kf6��[��n�joS}>\���y�ţP�H A�>�`��.�Qv�����YR��R��� {�b<W�����)��ig��E`�dO>iZ����D��i'η>#�j�"�,���ڨP�g��͘n=c�~�X�6�`rP�3	Er#t�4x>�1uS>���*�X����Ҥ��f$1��E��q��u��2^���K����cGbo߀T�u���RoO�*m�^��q{r�R�����1c���' �>#u�O����6�ەqQ�OA��.��:A-[ݕz6!��=k�t��W[���G\�N�^�l�,慞����޲��-�dL��ZI��\M���6����~;u&ͮ@�+�;V�f����I(�w[ N�RW���H��'+}� ̓1im3dHb�R��S���ڦY�E��CjC喴*��؊�p��nrm�X{�~�u.r��v�A�J���-�G[ܖoR�H�Uj'bLQ�)��|�O�X� ��醔	bt���:�߶Ƀ&3��Mm��M�j�v��v�C+v����R"�4ײ$��%{Q�.�;T�]��` ��/��^os�5Ý�+b�����9��QU�v��
⽫Me���>*�sz��t����Drmw�
�.��* �{����P+l�� 1��q���f^�x5��I��U5ۿ_�e���ͫ�k����r��x0�P��#���	e�eF]��:}z͘���+��Ùb�l�F>�]!�4 W��PK	Y3��u�eɍz��OI�,�x�.H�w�B�Vg�-n��3����U��+��GӸ��l��9����7[v��1�-�nSTKBy�,ib�$9;5��͕�82;z�^����v��o�|�[����~lm�S]3���ު"Ym��J����`�e}�w��Y����fڪ���+��>�c���&����x���@�h:o��Wc�'�tc6ȸ^��G˥�#{}�h70�mL7P�XQJ��"�pb�#��d�L^�Wx���N��k!��r����v����b���Hcݕ�ւ�����{�'�v*�u��^�$�okg4�!�YH�T�c����/�������|t�6C�P8F��ot��i��9ja��<��:��J�S�]����(�6�-��C�SV�8K��4�u!����c��B��T�R�Ħ����Nw����aV�P~P��d�#Ѩ�n����]ۣ��7���
i�H����P����t:�Z�q��Gx�(�ނ%-g�~��$�.܃��a��]��y6ꓳ���^�f����;��@G�H:��Z�Ѱ���Y<<��꽮�X��*f0é)�%3W�q��U���|pnrJ9.���\����$]�(e�s�hal����T�A|n��ޓ��g�~,5�tE+_��/FƋ��-��Ru��y麭�[W@A�F�Z�(OK��qre㉅6[gH�~70��o��u���X�e���:t����2u�Rv��ܑ$���d��3�	���N\	btE( *Q㶖�%W�m�s܎ٞ]`��(R���Iă�1��,h�,E�Ǧ���kRyˍKoC�-xPLܗ�,��  ������r^�}�iGB�*�@�'��:�f��[�7⋔��@7��۹E��0�>Þ�x�����9��ޮ�$32��L������eṉ�Iq,ank��LtQ���7y	�d��p�b�Di��x���N��m]!�N?���?�	��6�I�7���b�26OQSI����j�E`3A�Lkp��bn���+�1�E���3k�v��J��J+��U�:;l&�ݏ�'G��C�)��c�ԇ�G�5������ڳ�M ��<�v�����a�
������3�V�a6�s���������/"Z&JE��P(U�R罧Y	2B��2���}Kص�H�o�?q��`�5�@��Sƾ~˧�f�#�a��0������j�>�ez#u�Lm��E7��1A�Ь��=����:�I�+�.\��<���m
���\D�y(�\5��E�C��G	C�\jlkRv�q�`H�9ٲn�iY�I�w�"��^����ݲ)��&}(1����k����j���:���O��Gh����;��<͹�v�{؊pB��k�����ޠ��8�*zL�}n�2� �=�]�	E�M�SV���1Q��,@���&�Z���!�z��u��j.Du�_��%�	��<6�¶-m���u�����7|�ҨO'mNS�ƅ�{�*����F��������1J?9a.<�R5��I.� ��mE.!"k3BÐ�!ځ�vn�=x��_���a�M8�JW8�t�	�a�!0�� �Z�dd�lc�eQ'����(Y�s��J�j�-(R,��n��3m�+�]h?�K��ψ	�ٹ�l#^��E�M����1�a>zL�RE�X8)��Wߧ����#�C��L5�>�YV��x�.ܛTb���x�e����'� ��n�L�E����tO��T^[�+������4B�g���"���# ����~VO�����$��,�P��)�e]@�Y�h��n�g"��_���&=g�xE�^���'D�P��+r����ʙ����rȑe�(���_�aE���*��r
WN�Tx������*�8m��r{��{gVp����gj����"�&W�(IJ��p�C�½�ѻ��'tv�:R�q&�<���R˘ei�T��İ�4�.5�ˉ��Պ��b{��.��>|���\\�6ƌǥ^�ڣ�{D��L���1�%�������#a��cHi��ɼ/�Ų�&�{A;�E����G�y\W �aT �W�����eAQ�|��U�Y�jͫVقȏF��#�/�X1��Za�/:vei+��4�����
�99���+~^��$3?���"���מ����1��azȵ
ކY�W)!���:w�J����n�m:A�v�5֨;ң`���������_�\w�+�|�����|k�=[��Nj�"��%W�1�^�tӾ��4��'�׀"�����2��� P)����!�bpc�XE���rsܲ�0S���N�O\�$l(�Uf��X8�H� fx��H%C�"���6LKsq)�	A�@��BO�B�,��^�G�M���j�G��c���Ѥ�4Lh���"��늿.Pw��4��dΚg�&�\a��DPF��h�!l�R@kr��j��g^o� ��x��ib�����y����I�fU�?���_���\Kٸԣ�M���Ʃ<��T [�;FrI�k�fY�Q��,��PӣMK�n;@G�_�Ev�MhaX�uژ��JV�+����>�5����N|*#� �W0D��#v��t8�Zv~%��C,=���h�����`ʥ$�*�]����\L�'�سR��A2��Ŷ�k��f�n��'�2wO����w�Ni���J��v����/��!:�Ҹ;��	�pN�F��0`�{KXbO|̕�іJ�j�T,��.���������M+C�S8����,0�xrG�fl!��� R�6�{O?���ꧫ�����UH�z&~;�{!zL"u��P��`��)�b�-\��@*k�	9rw�-�;�a)܌O'� �*=k���+`�x���d���P i(�|�|������;�S(��QLg��� `��5��?�9���k����������%��j�f��3�7�����*\��:��T�V��έ���F��+�R��x	�b�󵑀������(p��(��&",f��>T����.�B�[�36k"4�v�~��Y�M)�ݠ��TT�䁪a:�2i�>�z��V	��\٢��v¼�.�}�#f�E�vJ�ݧ@�&_��,e�Y�._|5�8b �$-�7��n`�=���qNJ�`���#��!��@t�&(6��۰N��8�s�5��8�}��`\�{�Q��2�qJC���h��5�\�SO�Av�	���L�J��q�e�����/{�J��ˈ��K�)v~��UĴC �~��V��NKAE;�#�Mٝ��GIB`d1x�w[2�l"���4�by�= Z�|e�-�[�l$�J�ra�Um\e�K%�sOt0?�{��3+�k�a#�$a�j���@�3z�d���+�o�7�U���4�/Zd�^���Pst�"N?I����<�M]�}��-�� ��eD��pD��?����^� b��$��'\�xK }�����k�b+�>λ�z0�j�=3��-|��k�1��o�8����^�fq50q�B9c��˔��"��N��D%�)���8�rg �_Nۋ��4f�����m��7�X~h������O,dyO�x?G�<���Fm���3bS��b���'�De�lӭ�{��I�>�\�������$y��^O�cr)���ɈBZ2��K�	�?�-��pH�5r�<e�?�/�W�=��~d=|ǐ���\�s�t?��]z�]Y���h:,��JDnse.�\N�ߝ���W�Wp�N�uo�I���ֹrs�Aw.8���s��敭YFi����+��e�׬��2��aV院�8���m�1��X��E-���8תt������_�ix��a��bpQ��A�Ę\�ֲ����� }Dh�M��[����
&�<W�(���?���1ҿ='��#F�P�j������3wqM*�����֒X���ν��8�ﻉ�.�鹺 D���b����t�W�vsQʀ�� ��' "��sT�q-T9��;����~���J���},v�_J��޸ۓRt7����S����T��[t��� įo}���ܚm<S
���4�?����{q9Z��o	鴭]��9�D��Wz��v�p��Y�P'#-���sG�	m�C�.� ���r�-�H�[~����єS}�~	���M_�?(gm��;8�v�r�
T+�3,�m�IM�f��5��peYz�{��|��H�����^IB׋O���V_��>۶̨H�Qߺo�t�W�B�\6@�X��`�j�iUx�dw�G.)�}���ۏ�*�$1K�y��*�\5��� �3��[6썿�)
=?�7����g3��w��n��7ʹ�K �)x�L�D�J��6P��|���2�O�T�f���|�R��g�/6fW�4�Y�ζ0:t�x�B����㫺�m������ɵV�bh�^�&A��������ds,y��
(�������jI�:��Z�����B1�#��a��؅���H�긒W"L4�=�s�t1`��N�(�3Y�R9U��>���b ����x��3�}Ay��`��ƾ�nv`.�\'��$X�I4�b4Ȓ�2\ي�u#3.�~"����l���\���Զ���(K]	�i�����c�ڶn��!iK�>�����M'���Y����6Q�@����\�a1p�(��S�����Ⱦ{���ˬ@I���ٗ/��Q��M�%��	�%S?�<�F�m�z:�k���{�JnB�&;mY���� ሟOw/�����W���r~�P�,��`k0�h����3��'2�|�N�>F�ԍI	B9�u�5x�{�ŗ����ƚ�`�r#2�|2#��A��@USX�� M��@΃�h0�p����@��)ԙ��؉����xu&SkhKd�͏ڠ[�8P����+�0=#kÇ�1���mp��DzS%ۃd]O#>i�M��Me��$��O+֗@�r�¼&C�F<We�M֩;��櫍��u���Tf�D�ۏ��mV{X
��ٿu���!��$>M6�����fm��_A����~�&Ի�Y�j"ʷs�aq:�8�Ê27�YQ��{p|x��:i���Q���9G�o���8�����45"��9�Fx�8������e��V{T<��B*m�`�Ú��J�Й�6V�D��B37��Q�Z��'�b~�L���Jk�w<D͍z�!�,X���:� b�Yt�M��?[0�!�T8��T���ʼ�KF�vĢY�9�겗��z��/\��G��Gn#������a�Q-�#����;�� -��Ҩ }��mg��,�w�{O]^��p6^��+�q��{+۬7��#ѰZ�h��Ct|����=�L��}�+@g���rs�C߾
��T7:5����@��	�P��}&i�H�����f�?c�Db\*,�M�%�l癷>��b��M�+k���K`��M#�K"��W|�B�oDR<V��7~�j̺6i��[2OС��tK'r>��8���- �p��BDRJ=zhE�7�KQ�"+Z��c:����P�v�=:	q�q��8ep����zD��e9��E�&fS��1<��FI�;:g�.訌ӄi��&^צ����q
7����J#p�%�b��a��D0}��� �T\����K=Zw;����.:��H~���f0��%]3�DF�,��	1����3Be)�wݭ7���X���KJ�5�&i�_�U�C��*ץ�o�a�8ߖ\�WoϨ}����5$o9L��F��:>}
1��D��e���~��V�D�x�@O��	'̑b6eK��Q������j�,|�bN}��5
�`��<.��7P7�lc����+��z�����<Y��?h�5 ��{�q�h8��XZ��3���U��ñ�s������D�Tbm���v�A�v�*bo�i=��ⵂ�)rFO�@�/��{m�t9l&��������l.��3s�BA{�MbF�����! c�濽��+�L�����s�P%�r��#�5����`�!�)��,�����|�L0�f+��1��i^�!N�pA+�a��P��D��X��}�c��`B��)ݫ ��)�����"�dA�r�w��{ug���"�U�7�9	�Y�Ͷ�������.����^w��|բ��S�u���V)GF,]�Sզ�E(���$�~Ű~�g��Q[-I��f뉲ڙ�4�n�-J�� 2�y��P���c�w!�ަŮ-�  �#�x��=i�]vwP⧬�ڞ�:��W������k�#��#^�o����I�
`�q�6�ލbY�7�����B]_�����W�x|�a�n�/�8P]�K��:��1zT��2��~i�}\!�*���?��CG#�0O��G��Q3?����ԋ%m�DG���,��-y}�e���] .v���l�ekؔ�y�f	o���v���x�ߵR�m�d�K`����yh�C8QL���YT���a��gX|vݘ�$���[3���Z��Qb��5{V�Pn�p0�|H}|`�↲�����]h��X�i�f���F� s�5-�`��#	J=Z�O� ��.?3Z�0v��P>ëg���_*Ԇ
���7�����B򮍚?�H��\S�[���O:�;٣~G��rI�Tħ�RC���Y�r�ǵ�dy��`_��M�(�J�6�ՊHޯz�P0�x�x��=���4뷑� ��iC't�2`,0�u���>�]�EDp`]3?C�mL`��T)�\hOP�N&[���s����q�r#EG���ۣ�Mߐ�^��^-wSB��)����#�b�E�~#F��{N&��Xpøz[�*�\E6BJ\A)�Q�
�����iwS�N^�OiEkJjn�a�˝�����J�3�s{j��]��C������*Ǖ�b*܋ _�����43�컹+J��gd}G�����eY������[�'�Rb�5Tr ��zs.ul ?ڑ��!��@P�\�����������I����W3�4�A��G��/t �m��m��ҰG^�^o��O�
k9��LL�G~�3}q���zʖ{�JBh*\Ʊ)\+4u��" � I��;��&���U�.8C�P$��];�?���7�t(ݶr���ؠ4C�����˾��]���Y�*�f��H~�d���j�3����Wە�'�+M���y��p�I�I �
O�5���/=:(Am-@ �%	HGxo��XL�'�**��'N~�6����Ҫ��#2�!Ng���ꧢ6o�δ���3��MBZxu�G�f�E�G�Y���\�)ǽw`�\��K�*T���m슶��K'g2<w$��H+��X�`"���ÄM�/��p&34�-UӬ�f6�����h��� ������$����)��!�UoM!���g������B��9Y�H��$���Έ���6j7�U����{����ٵ����V�lf��Z��������i�D�}t#���r�_@�5�A�to5��)���>@K~��Xi/���?&��\iѼ2r������q�n�������Y�PJ�?ή��˾��]v��'�������$)V���G)05��k��T�����6������o`�KN�#$�)|Mk�2�EN�t:�N9��x-��*�e<N�ϸfy�|]Z��������)͈� �Y�qO#/���"����I6�D��׀p��r��wz��\b�5}��-����y�sz�"�t-UJ�?��R�ς6�p��r�k�xf�}�j�Z�5�m�*�2V��'΄O��Йr~0�&B�l�'�����blwRVvC����,�J��0����#������t���6u���ivV�N(�#V���|��=K�݌Ik��8s�4� �[��6po����M��V���Oy�xӴׂ���`$|�3o�|�z
���=�V�ݴ2��&s]��6�j�^�jf�#������T��l� �)���"�Q��)��Xɂ���[�q�Af���ᆡa�q�5(� >۹��������N`b�CPZ%�Mt���$�Qp�8�ӷz��h>'�����1V�Y���JO��s׀�\pa���X�^�]N����o�sOV�������@?��D꫈t���6�{�_����-�װ�x�9�i ⥮:U��cq�wh�D%� �Y�&�<u#�x��M�Bb	UY`�������Z����x}sB��U1�w�����ێ��u��g�Pc����=��Æ�O��I��>zیg��?[p����?p�χ�^G�"�D[��e������%P�����b�3�w���k����~QO�w��oV�۶�2v��x@�n�4��X�Ү����x��~I��������.�@�3bʿu��Ժ�������e��-��+��0��-?>�n �F���D���Oa@3�ߟ���U�����NH͖�olU0��,�Ip�������T6���\M�Z�$^�E��p����ün+j���M+�b
�1 *��l��)l����,�g��xZ�
-�3��.nƬS��� &�0�G,�@�P
\��[b�#�S1�й����VB��x\w>�-ϡ�ǐ�j\��1�.]#����w�#���)*�����b�{��ν�x�Y�r/}�UJjs�6.����5`m�% 1+$'��	���H�4ۺ/���or1�8�B>:� ~�g�UiT�ԤC�|��9��3'M���:_�)�?9�~��{��q�����̈���9�{����(�~�7�ɇ��Q:q:��z@=z��=��l$��@1 �-M�f����Eˤw�<�㌪7�F�{4l|c�{ȗՒz�풴�D7+�Á�Hw_�ޖ�Uڪ�C�?�Ø�Լ�B�Z6}W)d��\4���-��*���cTַq��ٶ� ����q�VS�HL#���a�k�c� R�-����Y���L�z�W>�yeUԂm���*�b~ESo!Ʀ{�[��p]B�ǀ�-|G�PTt�p��,��Z��͌7?U0~7���5�y+0�,wk�SN��ծ�^�o�
�$����=˪��4�Bw��Kx�<��[��k�V�߿u�;�%�$O�u��{TA�"r��N<g����2#
9�&������|ߤ��
?v�y~�:����|~QE��\f���o��Ox65�S�Km%�L'��M����t������ԫ�p�EG'�X�y0��3pRٳu �����5+( ���I���F�t/�}|s���`3��{;n�߬��By>�@�v7$�U�= g�.\�rv=�>uM9�e�����{N����Ğ��4F1���#�P����w�sO̥��-�*��	�eX� �}�zۡ�Tc�iG�;Gpg��7�q�����(#�����zި��v����+YM���6��fH�nw�n%o����e�����G���%F��G�GTb�T������~��k�l���f��"��@H������E�=����Q�X����d�	=y%�)�%3C�y������<��]�5����0]7y�L�wh+��ɝ�D��òs�E�r�W`�<W��2�}�ڂ�Oe���)P�~���b^ۋ��nPn��s���a�1�MW�O�]�`&+Jگ�BoBO{�$��J�4��3���G��@)�#��e#�.1VŇ�[�nc|�*+L4��1,&,��wH�; �%�[[Nh����}�JLUSI4�S^m~����<^�|��n�U#�Wgp���=��	I��+�-_�����1�s���P^�x�d<�)j�@P;4__�8�[Cp.��zP]4��,(���K��u6����bX|tcj�"�aa�{���֡&� H?d��YD���꿪��;'�o���ͯ�����3@�o5w5��[�Jn�jD�/��O��bt�s��'�)�P 	�����t���Wv�0.g� ɇpF��Օ�\�b�����c��	�uQ�k%~|ƙf��*���r��>��"����o!W�����0
�b,�"Y�鉢�6D����ŝ#�%u
�s'�|'�;��JYw���S_��ݨ�����lv��R_Y�yG�.�f���u�8��sh|s8��� ���;txuROe|d��ˏ]X�F7m��Ur��E�qmN�4b��Eb�<�A�&�RA��z���xv�j��sS�@��(������؛��X���p��w�%���W�?��JE�Gh�8��3�	ۇ��kڊ?%�w���J/#0̤jsl��8"D���A:��>��iݵc�(�SV���Lr���h��6�f��m^���}��V3�D�'�X�(=�6��m" ��S`7�Ƴ��dc͋�YT=����n�lH�:b����֣�#��l�Ƣ,3,�/2�ѿ9j���TF�S~&�3Y�󂭘�K�Z:Ͽ��>'�DS{�R4���l"~�J�GLJ#f-�J<�H9(���AHgi\�o���w�S�?����'5|��|�q�\����Hi���ӥE{��Ћ�[X�
�c��,'Je����AUz�f�#�j�cJ ~Y��*e[���W�U� �Kˏ�,FF���²-�������ys5j,��n"�$2��@`Q�˷r��yh�����3]��0�D�� ]0I�dᆉiI�_}�W���;k>au��J��\�����E�����q�S�,R�m�H�*<�FW�i��X����W��g���a7n�e�D,�w���z�4���<�ћ2��/�t]fݩ�,^��v����U�c�{�Mü�Ьe��$x����/.u�dqcH����I�_������^��"�l����:��r�ΰ���tT���f��rsXE�]x�q#/d��{�6��N���kC�pb���IzA�h���=������ѡ���iR�q�� ቇ���1.J.@xG�R�����6�2�W��cKVLf���Ch@�N��$u���6��ۉ4N��(5�7��E�a�ߣ�w˟Y��D�%
P4�{�+���ܿo��b�bJc*&�+���qi;���UտE���A��z��A�v�����qF^i+EM��<���X��aC  <z0h�ډ]�%�ڶ�'�ȟ��7��[�f�|��!/|(����V �����my/�C�����g@�D�S]>#����ZB�&��SG-�ѾAD���D5���z	��P�}������:m�K��=0���(Bs6	c��� MՑUɔ�Ԑ��#=�egp���x@��9_����$ԕ�4]���0CS�����v�AEl	�x\�f��	�0���	��;J�P����ƕ��!��L� �F��J���Տ�#�3J�3u��4dQ���@諫j���:ʴ�b~%̘w�%�Z�^�g��c�/
V��(G���:���s�����x�P�#���ޒ�.2`DDAP>$���������M[-Uwt����E��olk�s�3��PF�"�#9���3J�㽪m�t֬��#�nz���� �ldu�b���p��"6��"�S��l���G��Pt/Ctf�H�W�����v
�U��=�e��O��N���m/�\'��M���n�4Xm�q�W.�}-�(lo3��'f� �\8�]>+�����J�y�d�1�sW6�cr�Ě�,�(���?�4�=���ی�Ƭ9���sӾ�>�;S����v�`��>D�;;ל��׶��dV��E�K޺�۽��8&�<����"�����M��>�~n)_��F�'������įLІ���@�4v��E��&����|�Na��w=hq�M��[W0��;v"X�y����Lex�>RE�f�ޕ4 P���v���2k����}��(૰Z�&O*I^ɞ�����}$��j�Q���v{P�a�xwε������OgwJZZ�| Wi07@_�jH:pGL�9��� V��!h���|�C�����]�*��=kk�Yɚ����zht�|��
�obp������	�?O+����cژ}(cy��y����ɀ[�n�I�?�I`�?�E������zw���7�8]�Ʀ[��� 4�2�֤�O:<v�M�]'��er��w`,���n4��fH����OY�7���xOr�2�:-3gM#B�EvDM�|?D]��UK�=j�A԰�X�� �����6���FX!IѾ�����aۂf#�/�y]�sG�;P��Ś�����Zۜ�tI1��F˱d{�rG���I�<��X1N_�|�f��g��'#��	X(�߮H�=9�*Z.SFj�C���4vu�{��,��R������������s��I$`��~��2��XIG��nKu|^b�	A��u���=�u���&��h��i�iqI����z�i؃
�0Kv�k#"Y�|�X��އ���#����Շ�p�P�~�j�g�2�pM��O`�������^c<X�t8�����n+UT�uM�b�M�o��r,_�:���Q��tЪ��-�r-<~1r��	7m��� 3�Ikaj	�ҟˤ�\jO���9O��� V=���R�0���U����>�B7ǒ��'�O;0o^��n{�G�\�D�����!�#8��T�	��h��תawgX���ޛ��&/�S|�,��Q��G�<�>�<>�E:pl��~��{�T�wѩ�E�d�o�:&��e��A�h|��x�n��'Y
%4�R��or�
�aCr�t]�/�ߙ��!�z��9���Z'���t��_���I���'7^��l3�G�;q$�9 �BiE�qhS,������D&UE�px��;ͼ�W�u1g�u�'zm���%){1*��t�y���0�>�@�V\�4��fҙk���<�TJ��.��g"_+�~�Ǝ����Y$�[�b�bOEX�]������������ �J�D�&f�oF�S���M�g��|��P��;�ه�+�/��B�w��sB{1f�&�9G) ������w)@��Zm��J��E�R�x���" �y�"X�8�e/ǡ]�"�X��`�R�Q9�g�4���L9ۣR�r�/�rJP�O6n���g棂��m3�2^'�Ou.gpz��"#t�)�n�̠��fs����ʔ�E|�>��"|6�&r<QUz�t��|^�i�}U
5�����&�����������Xü�S�c��B��缊W3eG~'B=%�A}��7m74Jc��2�ef�ǸAk����s��E��]�t�'�G��ȸ�l��F�7�%Z���y	���߽�%�'��W��w1����; tN�N�W􏑁��^ e,F�����ø��i7:j}��	�;��[�����Z�9�7̊�F����'8K(���_PL7�MhI�u@⚉0��_֒�Tt�3��m$��R׮2���rU��:�;����#�І,D�V**U^�Mł�B�wȌ��CȢ᝽���JJ��w9�7!�8�y$·���04C8��5|���3��g�X��5�"T�B�$��be#T�<e4i���ȏ>|��KߊB:V$�T�O�<������r���<����:_�|D�sm��~�}�����Ñ�����>O�*'�ʸ*)��4X�P{��M��\xM�}����}��pI�V��56)_S%S�tEH3�5#��i��:8�v
�v��#Ԏ5����dZB�)��4��{bam�)FH�U@���.Ō<�#��kN���G�􏾐��W��ܺ. "}�<i��򤌶F���|.q�R�(�HV���=y>����������I�c�|�N�k�o��N	Hf���߈%�k��|��l©��	%nB�&�5��T�26��Kp�k�dc��>(z
���N�pb�b��(����=�wi9�^D���������K�(\��+QJ�0��*��LE�1x�>� �NG��QǈW��)v�d�>M�p���'���8O����MoJ�oa�Y.�DWG�֘P�~N9��\=�6��`���ERH����78/\�h��!8F5?-�+/Ӏ8��#^J��ж1<vɮ��2�RQ<�e�^��:�����QI�E&���0g�!�<�0���D�5\��a�L�5����ss�`�+"lA�D��=�"�sXT�K
��P2eL^J�{H!�ˣ�D�[�C<��Q~�3yg$�V3��b��6��6@��'���տ� ����B�m�@�0��e�z��Z~(ˣ�`,�fh4JU.)
�̂v0���VW�iX���*��I�w�3&?|0�x>���)}�xē�g �s\��
C���"�
�O&�S�e�c{���@C|��#��K"Ɯ��(f��NI�B�Ma3���z��Ղ�@Yy6�KpV��;h H1(����7�%�J#�ؑ!�`�30lz#�&�UE��Z��ąxmզ��/O0\%��9�T��z>����q���/�48�
�i�dze�hE4O�$�{[��hU~	@{����u$���;L���F�h<.�<<�uu�w�(8V�uV�5	ڬ�g�ަz+UD�� EN�
���D�uѷ���8&�)%�����]m��k̓	uL��'@k� H6��%�!�HѲ��'f6`5�l��5��e;ܵ��|�GwI��G榏������ɽ�X C2*Xϻ*�eR�vF�����E���vO_����櫊�l�^�_)sgbKkyc4�j��A�L�,=�����^:�>�L�Q�X	��폊x�XN��{#�ˇ_{'5tF	��c��~�y�C�Q+#�r+����Q*rp;�m�O���k��p|��u�J^,���)>�������o/�`��*�|�����v�RO�^����Hf��W��||:I,���bZMBU<�T\\���FQ�H:���Y p��@� H諍f��R[��Zݴ���'��Ν���
_�m����/#�"C�xP�O�,^���H�_8U�.pڠ�e1�6�N����z(�FoE�`]�@΍يp6ϊ�/w�{Z�%�}Y5�5;q:]�`a[gĕ������N������6R�k��~ �U��NU�,H��M>�憵���$Cl��G��'���u>��n�,�URݥ���I�*�\��ɫ�$(��!v�t�~:���$�d�9�+Mf�OfLy�u��.�~��.�J����~ؔھ��G��I��A,��m��0/|࢐㎏�A�7Z��c����Ħq��A�:3�,�saFNA�n��䱙�@�b���,��,����:�3.O	 )k�EUĆF�U�wOX(fÎ�	�|3G�s�xH'.�O�AE1׸zO���9?e��"!s��q����'YA�9*?�]�t�r��+.�%#��?;�/Wk��2�}y@���fX����щ����O�4&_����#�f�c�i��c��-&韦7���3����6�#P��nR����0��.�/�.���c�Yk� Ns���0G���n0�5G��4�t��yv�Wc�U����-'�8,T�@���:��RU�`�;DV��>��\C9߭��4Fn�B�w;f�aAr�س:z3���<t�D����淎��.���Q?xs7����]G��b��ֵu�-����W���DCL_�T��(*�����q��!��U��^�
��}�%�ʛ��^�Fޮ �ȸ�4 �q�Ǯ�`F:[��
�3����$�n���8С��X=��O���"�fґ`8� ��9Fv\�R��mGj�Ոaq���wg���Q�Wx�!���l@ǮR�/�-J�3���k����B/:2�죶J^_{={�,��Ӷ&��U�[.�Eż��/���uu����z������<	t�p$e�Њ-����v4aS7����]_"����ۮ]���T9�|�{��0(��M�tO8�j����c4��sc&S���?èUԾ'��~;qK J�� �%P Y/�(��%f�zr�Iy�����]>޿��t��u��a�#�j�E�Fan�����P�$��!�k���죴'W� ���,^�sl����S��}��
�v��dtItC��cW������7-ѥ�nu��9}�;�zy�œ�
CrJc �(/!-s���׵
��O�n���+^�_x"͇C� aTB:}J �޳�M�Cq�xs�@ӿ,�~�)EE��sN���P���l�J������l���ԗ8/���*�fg���=g�(n����.���ɋה	���xIJ�?��7I%���=�s�/}�txg�`����ht��1�~��k��yVrJ�J������P�~Ńa@󇑋��8�O��������d]�a|)���d�M�Az�<E'���5"l?`�r10 �H���4�M�?vL��A�����|I���d�Z�X�� 3���Y�7ʀ����e!<���-�>(J�_�<�s�L����p����W���ʤ�e���6��'_��$��]&wN!>
�̃��$�N��m�P����4�}��5@\��CY̰��ý�4��p�5'��ĴT5�>8)��uy���y�jF�NP�n,�*�Z�=9QG�a�Y���^��~�}"P�%f3[�Eg�'���G���f����æ�bĄ����W�waw���9$�:��xx�C�������o�n��!��j����k<r;�K��MD�9�bL������д��͍0#��/!��Q�Ĭ*{u".c�`�e�Y�cg�ȊK�P@U�=��R9x=��&��7ޱб�����w#!	A�}<0êP:ؗ��A{~Ir����������ӄ��f �Ire�7�CR.���څ�.U����u(���[a��Y@:�ѦZWm��d�ec��赶�4���X][����PGM��nP�heO�"���5r�V3��؍x-͒vޓ%s�Y
#��Ħ�O��S�oSb%W|e;�����������W+����Z��w�N����1� �u	 �!^�p����*+u���І�W�w'���n#O��b�W�T
E��6]�*8�vT�Ë�����>�@�P�&t7�RmV��(���>׽1��h������snfݚ�p����W1ǐ�:E��lF�|D�X4`c�P�����C!�?�@����d#�Q�#������S��b���OFb[,������Ň�vw�R6��7`�����f�ָE�v�vp��ŧR�I��FdT��eT��6��UCyY;��((�iȲ���L׬��䋟o��vW�حȘ��W8v��~�U�iN���%���)��z��.�r�]H�񾃽͎��e��ʣ�pS���������z��^y��V�N�uV�E�6�	y#��u���4�P��V6ϵ9��b��7+u;"��j%X�����6��>�6�.gR�����t2pˡ*L���|�������J$�$fG�=�h��w�r�߈<�*4�|il%m�lF���O�e7��]޳2`cU2	�ڢ�@�ή��6-B�+�cU���%�I��֪�GM�x�=��+Ye6�K��w���_���k�^�z<o4w�mY��&d������5����6I��PK��5���!��WK��y~�Jz�����&)��w�m:�`�"1�2��Isx�H�$�C��'�<�ц1zf%����Rt~�%���,��KKv���]�������51ͷ��i����<x�L��c�	SW��^6xΥ8xhI�Vot�+�9�1�iAr~>��aЭk��Q���.�Wg�����G�(9?6���}�̸�x�l��^��f�so�ȁӱ�2���#�ҋ->WT�v��U?-}���3�>A�b�	�C������̞�) �D1���{��*%m����Y��W�	��#ɁD���������d*��pg�"��f��de�TG�L��|*0U1q�&�&���J �}���y+�kԔ��Hp�٭�K��]�d��m�����k��,��+xh�l
���PGŊ����f�%U�/u��^�D�R��3�N4F�h��M��ˬx��=�y��a��E�x�|��:�xB%���Tv�j�^)_��i���9��!�]y�T@���@��_HFta��q���X��J���բ�s�<������d����oFҝ��8M���bA�g����l"E�H����飱��9����-=ތ i,���ye��O�Ҵ�gWc�ϳ$� �(z�p�A�wt�:Xf���`c}�z�R�!uq�Y�[������ K�S<�t�oK�HHHR˦��I��x�/H�M7�lpof��%��)�N�s�i�r�>u�6r:�� �7n�}��>�O�Ⱥ��V�{�9�<qڳi���I�J���s~�Vٺ=���v���e7̲�/�v�,g�H���b�oEi��A4����M�K�Zӯ��kf�W����Lu1��D]�\=���#���Y����S����OGZ<���T�[ɽc��a�M�5�`�2<��I��M��"�T汕`��{��E4k���Y6�^�B'00�z-!�4����(DQg��Y���Du��K�~�L&��|���$[��� tr���X�[�x>�M��CoK��`m�$b7[��C�#�ʓ�)HG�t
�v���~�ϭ���^ЬM`ĭ%O�նD;_׎K)�$z���FQ����!��/��R�*�U��%�l2Q�a��zidv�0��	}�D�
�������GmU����w]pY�'}1�p��ѾZ~����@�I���»�yA�![�R��x�<��gܷ�lp��(���m�Jlӝ�**�b��a� 1������S͋XF���w3B�*#�[^2��cv,�kd�j;i�|r�����Z}�Π���]��t�� %o��MD/h#��6ii�WL_� ��{�(&��ړ�����}}W� 85�Mo���ySg� pp�a. ���;������W�Y5F�-Ƞ��'J��E���9��n��-E����;r0�$ �YM���H*�e�7U�--��,��k����$SG���GG���)��Z�$ʙ��4)ݮ��|s��$�&E�\� �b�$�Z�ߙ����E��V����N�}	i���F��l�[��Ps�o#�n�y��
a7n��|�^҆�mZ1��1Z힠�����F����ͫ2�W~t
�m�*Şj��Զ�a��_����e��@g�_+�L�� mt�X��C��dec �#0_��|�(���K�����Q0�lI�Zy���]�(S��H]����FAuM� ��:
� "ix%��F�E�T�sOD�B �����l'�^Bur�
DE��<�Uj8��*�mҒ����5.�N@�(��X}�S��b��鐙���Rz�`����H�Ĕ�v8Q?L∺���;�/����_z��DO
��0Γ.�����j_�IA VQ��V��Z2�	^�MW��lX0Nn��A��D�8�s��b�5N���v���A�᪘�?`��?^R�o7�F0�c�@ަ��&�dvw�-�P�� &ԡ�i_���Y`_},����1A嘄���_���b˒�e4�_����#
uҖ��\��=�U������V��˰nRh�cb%By�'Aݨ1�tc�#26]���x�F8;��Z( �P��Uȷ��L&W9�y�1$XK;4 [/�Cz�6ʚn+��n#�1Ss(M��/^[ܴ�羉����	؉!�G�Y��P�R@N-!�KuD��h��P�4C��Z�����G��*�!��Tj��ր@7��ݦ.w+QT������߬I�����Fr�7ʳr�Z�sM�<�*�V#r~X���e���K�� l�ͤ�z
��W���N?��߆ 	ȀHwCO]M!�/��G�o�,$�
��Ð�ߙb�W�Rww��i��$ٰ
JQ�V�e�ӹ9p����4ކ%��Jn�nOS��Ndx�0%o�[�˳���9�
�ʹ��&��P2�{���T�6�h�/^8��O����
-�|��h��S�����# ��gUu��iN�W�!d'E0�:����ͻ��'aTXi�c�.ڢo��8���V"���aϕ[�2�D� ����L���p5�Ug'���������CFF�-a�?-����m%Sg����^�\�U�ߕ�e���N��Ϩ�K�Xw��6w���0�H��ama�H��2���t^������d�q�y�S��s$ouw��©/��w�?��"�Ô!��Gu�oϦ�F�Pɱ������Bؼ����>��C�&U����7��r!%���yM���?�]�xj��!�׮����}5�Ěr7�F	[/�v�H��{�.1��z����aT
��VK���:$��|Z`��C	��Xa���6� ��2�U��'���K�~7.��8����;x����R���u��J��\���C��ӄ��V`s��b�`����P�P�B��B?弃�Q��mS�A# ��߹\[W�L
����2���/�l0�-���	���)1o2��q�.�`�H{�o� Uk��6l���~tg���$S;������-��e-I�����E\��h��/�\v�:����^�=!7nt����vRɮ�n�����Ri M$��-T(�@�6塊�^���k�������%7�䍁"�2isP�df�(`f��Z�*H����|�L�����3L|�`��D��a�xN����^�nX�W�5?��S��+���pp��:+5`�B)���9Z"�D/ �� ŴS���5����3rH�ι�%~O�Y�=ڹ	��W���涨���w��>\�Ig�q4�����?(Q��I��W�s�^	�֕F����Xݠ4c���`6���T]����7c�N/����{�� P�J��U��u��fL��_�����{a�Lxj����,CNzG�h�%,B!� =F��k�����E'��2�� ^�L6z�4˻,��^z�����aE��>~��*o����ձI�p����;~���g�����xR�P'*�v�����?�O��we��b@h�;�8#�Z�Mơ�k;1�S9�0	�����x�E��Z�L�΂�ZB�0<�=�\|�n�v��.a�-����]�'��fqRf�Б����Ҕ7@G�^��]������	�Pw���И���pS�,x}9�\Yc��Y�/�v~���X��P}-�I�PF��Y5C%���nj<���c���	-��v�3�X�2�E�S>z
�.]��c�d��m-c&�6S ^�X��EE��[�Ms�u��F��Ց+���k>��媮l�u��
L]M�0yS1"����WE
�\�N&�xx]���->��#�K��-p��Y^�oF4�B�?��a���S��ѧ��+�X��i���l�c�-�P�ۨ����,�z���:U`�p�}��P���M�e�l�k�y#Nb��l���0���L>�34N�g��5�r��o�х��d��0�V�}��!\��db�JiU$�+@�tL�M|	��)��M),䝞hR;j������.�w.b0�yŜ�{�젞'�ې���/��~��!psL>=s))�s��C(�����3b<�T�D%��Q��nP��Q�7P�N���\b�I�V���.���.���>m(d"�;�Y�w�Ce���h��Z?�۪�iXz�k�ycj�g_�f*"������0=[G��!�~k��Y�.Lh������aI[�k�ΛO���Fo����aFs����o��'�LiK�״V�v��}_�^��#���*�̒�v�_=F���O����d�?��W�⾅���Q��.�%���Ǉ�'���H"�؍,s�O�����|��#�Y�*�Z�,���u�q��-d�<�Ռ�c��t%_d��Rm�&9�h�=�v�~��,^��U���Ү{��*x�e�+��0��)�Q�c�"S;v�_�#� ��o���;�*,,��q�o0P�Ӵ�x�1iՒ�*$B�GM@�Dq_�C�H��3�j�Йp�5�k���ȴZ
�H��\P��W&���a���
QL�*{֊�rѓk�@��,Zm>�B�]�>����HXOdn��7ݰ�9Czr0�Qר �i�VF���cO_�,9���hf"�84�F��]�����+*q�k����?��<|��=�\L�`���Q��st��7����/l��~�:�RmGk4�����Tи�U����.��.ߪX��$�6�Oހ�m1A�x JHr��3�-���B[�{E*|$�,�?rD�;3�e�u�Һ����Y5&�WdtzH�����ۉ���f���C	�s{�a�CEb/0���fJǫ$x5�IPkT���[���7��턧�$q�X<�iq}~(͉,��!��2)2�1ᓓa�D蘯U��̮7`�_G��]����ޘi��Y�Pb�	�� �>��$��S<kG	L5��e���l�|�`�ab3\2��������ӾcKX|Qj���>�,�Z�v�A�%�5 O�L�+����c6�����%�IJ��um/����}7:��:���̈́��#��_;�jM��r̘�amy��3�q�����}j��3ô�4��]@��3j�i${�iT�د����5X�=Ȣ��w��E��N�&��k������xӯ^Xܳ���~�ܕS�4�덿��Y���BL�լ��U���#���]�N ���n�ң���ز�`��X� x�oO	@�yNC�����`%E����;�q��˞��;u,\��Y��e:�DV
I���Pm�J�
��c�e���|��@�_.�?�IY�=�O}���{�?�o��7�)=���w��9pM�tS`kH}�c!h�N�zEb�aE91��bqv'�$V�RAC�Kc��C<{�8���H���4,���;(#��ǔK\�,BZ��	b�9��ɗ�o?�Bؕ���o�}���}�*��I���^�Nl��� T��b{��][9���MWH���W�ŵ8�tnl_�0++����c�X���
*���W�ʉ ں����_>��Vα,��ҙ�'�%����G��6�nvx�1ۚ�MD���He*yZ.�[��-������{W��N�D��E�U8y�� >uR�����|Ǡp�`5���UM ��k$9<��1B[�J|��s�qu���"sn�
����yz���;�O�mO�0/`^-�����j(^���ޛ#�����z���2Q7��j��Z�R�#��v[ǀYK^�=X�¾�B��?��s��%��\ƹo��)���'���m�ɪ�n�^���V-hl���Ղ�,
���Z���5p G���(/�F�D��$���~Y���y��"�b�9QX�S��7� nwx������[�]���iN�byFQҷ"K�z�>��		H*��/���XdB	HA�6�=y�ݙ���{Z���ڨ����A��Q�<\[R�V�+��&6�e{�`����:�d��*�N��J}�u[&�8�O��l|����»s��݌���Մ1�hf�4Tf���F�i(���������U:Fɯv�XvS���� ��ڣ�L��cB�ڛ;��
&�V�h듾��X\,t�v0t�5�;<�7�z�ja3���b�!=�|ӿ"^Omg��Q���.����XnE��A�ڳo�%1O
�?�]���8~�y�d�v�/��׌�a୻99T�����.w_�-<�
&�LN�Z@�6T#/S���n,��1����m� tV�1�6{�bJ�z��Y�/J �X�1�m����h��a;�,�̈́:x�����^U�������E��fV}r��Lt�{���M��gZ��1I�^+�������PQDP��s��V��Θ����\�U�gƦ�P\�K�g��J�g���yJt~�|�xR�ɔ����Z-���F���q�*�l��gĸ�^�Vp��AMpqej�݌��z�ϝ�]��q�Ԏ��+BH��O����m+б{E9ʦ��,���K�H�tF2���F�dJ�7H�r~dp�s������Dzav�����=�Ӱ�".	~�Z�
Y�J�:�	��X9M���sIc=���j$�t���ff�����p�Ric5>��?G�P�s����-��>�)�ߎGM[�5��2�n�#5H�t�awD !��C��+�C����'!+�&��KY�	V ����S���f�7��c�f��џd�7����}�-��#M���[ZOuqJEBy����4�9�]�6����p(&f��o�w�ˌ�|$f��ʜ|Fn]ѹ�W�B��6�IP�� I��� gK�gn�7�z�z%G���X^GHQ�׎��k�@ƀ��M��WB��^�[�ڝb����p�
` �A�H���<��$��[";!`� �=���Lh۰EiD#%�<����v��,�zm�͉9�4E�;[�u���n�'\��X�8���R# 1Z� ᰥ!�k�����h���[xU�̤}��_���I���7��c���ym��I��zl�b�iخ�ǹ�ufz��fT���2m�e2�s"0��	���Ǭ��:��$?y�9@��E�i܎%� ćI�iCY!�����(�A`���$KQ�*�I�r�Z�$�_3��AE_���ʪ)譓����?R9�A�;�ζ��~�^-��H>ǂji�.��fQ���>�`Ȑ�ǃS�t@����eda=�m���H��a���X
hc�U{�!���
�P! ��h�W�Y����s�U�5��9��#+�ܺ�]�)�w��.��ގ���4��>�����Fph�h��л#\��w��t����'�H�;7��ǔx���e-�$� ��]_i^�oX)���-:�C��jVGC�����匣��M �\�������4>C�nP.�/�oɨ��A+*�$���@���ۑg�)G5q �q��,��(�~R�� h��ڪ&�@ވ����{R�M��l��J�]󼼗�H2Q�Mt�V"����8٭ q����0�L
�3��xk�`g��(.��ۛ��g��b��İZ>����Ɉ��' ���a@Ƌ�t0_A�A�$b}2S�݃�r��5��?o���oD���������o0�Z�����0���?7��/�����!��fU�0K��U��薉^X����>:�W�}˶�5M~�E�����J#�}��<a��U��g�]��w1��0���dZ�yA=5�{���>��6y�i�F�/$��u�PϽ'���bm2��Y,�K�Jc�x��ǚM=8�1C�[����4�%'������{7���$�b�屣�)ծ�*x�� `���#�߁`��6��2�u��:�Ä��z��p�xq�c�fx���Lc�|Q(�_���nn�t V$�C�@�~�X���ׁ����r�ސΨ���0GS�`c8��Ss���r?�t�4����ѧ�]6���ĭ����tǣ�JzB��a����{�U��kӓ�����y�  |do��)�)��4��v	f�N�Ӿx-�gZ;o}��Ģ�"�Q(E͆�c{�w5z�`;�@vtَ�R�l��i�Cժt�
X�%�Z#�8�R��@��1�0i@=A�7�ۄZ�����k*B�@��Y�Ӧ����>�$I��&��**�E�
��18乞�+�nUY�F$�������8 УRp��Z�|����T����)w����\CL��Z����4߆�Æ��5���M��_���^�o��Կ+LU8�x�Q3����e���'z����s��6�
n�f?jx�H� �*8�(������L�Vʚ�Z�`v�W}%E�ԙ(=��{錈$RT)��4�H��&�"l?�
ڑ@���B�;	q��5�d�F.�:�b�'��ߣ4T2�� I�7޻=��~aA��[��)��PN���X!��b9��9l$�^�U���af|zr����D�xq��<���J7�e�o��C������d���z��x�/|`=����LU��fw)��ᜀ�"�q�W�� �[�7�7����g��3Τ�d��l/�m������E���aK��	GQr�(U���Y����!�����܃�qg�ڍ뛧]̓�v�D�L�#��_�52�=C���x�e�D����D9]r�)\���%��3��!A0�z~�>�k^����f`,g�l��@�������
�'��ˡ��H��$N缇�g�ݐ��礏ٍ빢�g(��*����6��0�(}���'љ����bDW�8Ͼ���;���hf�B_	+���U��S�gw��g�\<cZ�#����_YL���^���J9� �Y��:D�<=H�}����&
0C|��`�|ĀM�r��a���n����&�aI4�� g���D�n`�?�90�����>g猀r��ά�\;Rt��{��q�9c`�����yW��&5�[��f����L	�Y�&�u�:�eV�����C.w��T�%m�<ª�_�y+G�,�D�K9�lþ��jlקF������
q��n*G��KH�@��wK�ӹK��'�8F$�$$��z��@�r,=AY[q�|ߘ�M��i�z1��V8�23���3=-��|��`$%ͥ|lG0�3��ٳ�`�ٯc�-���H��1����x/�V֋ a1��n7�z�]�+�~������~�Lx�=¤�E�Ĉ��w6����<ʾ1�����i*K��a՛�Ր.jzI��+���1Q�y��Pq�{�N&e��!Dި�Г��0�O�T�2(IT�87-&~�b�E2t���L��,L"�|ఆ~� �`) �*�Bdm��V>-�2�����;9���O�?��g��"�FZ���:��s���[�=�C`L	aڜ(�,�!9����G|ʷ��@�1zF3b����T���>%�e5�nTbo�c4�-�~t�,YJ ��� �B��-�wVbX��=a�[�K��w��H��V��Nc�L.<l�MG�3x�����������F���a"W��<}y76_p\堚���r<�}Փf^�HϦ�ퟱ��Cυ3�5�<ծ�4Ul�;�T��v��o��J��{Dѐ�6 s�a`���<����Y�I\z����t3X*���y�����?׺�����T�s^�T@^���]�Iy
ǯ7Y[�ml�"�k�{����`Ӧ�U	�'��}ޒ�mԙ�3y�>B����]K޵�-�̑Uh����Wi+ѻ�j�#_��`J8
[�T1`�4�
����B�)ЮP;�����a�
JĻ0h^c9�y�>7��U�b	�w�v�VKo���>@R9)�V��!���̇��Tc s�<�8I�V�
@�
�����VK�ee�,�IV�yϖ�V�b�E�$s��lW���=��	�zَ4�kB��O[�󹪓�~`
��ZG<r@Й�[}~�C�mӉ��+�#������*�Τ�2M���܂�A&4Hs&P�� ��J�pG����V��BӖ��ؔ1���Lh���틮 ��2zF`�f_�Ńr0��!�/ց���|�V4b���'�{�m�F�:K/�Ch��.��(�
�k(Ŕ�y��N��5v���v3�:U��0+����{%��x���ލ�a��"���*z,�DbK���]V )���I�D-��Ɓ�I�dɟ�v���3� Ⰳ!�/��ԙV��Gv���O�u�.��{KgZ�ğN	C{վ�P*���ٓ��3=!ЦC�u�$[�Ʈ��u�7��9w���#>��2����#�<����&�I���[��MҺ�(�#�/[D�����0~�&�\W�@���@W|C{�ݢ{QV����{����z�S�0�UU-&��KJ�b|QxTWG�:�FG��~$�V
7 ̴h�y��#f}ˏ[��^�k�z�#=گ��|t��0m$w%*?,�&_�3�U��\o�
��]�-{��:}�9�������ޒ�%����xW7'ĥ,�դ�蔒�W�·6���Y�a��f��FiH���'2�����ã�Y��b�s�@qB Z�u�jP�q�n���te������a�� �w{���M��`�D��v�Ԥ��]�p��[@�c֋�cq��o�sH�!暤e(�o�L"�Y� ����	NY��y�K�L^vi��1ȟ<�-%��$�������ļG�x�'����[���g���E�l��àKN���8�����3]�w`^vL�8�pt�U%1�)��)�ϯ�m�_(#�k��[��ji^�D%�==��%~3�#I�0 ��VO~��J�YN.�l#�_q��|��dDl�hJ�@+�)(��;�kDqX���x�ۄ�K3r�J��ᣱG�N�Q����1�=hx�ߏ�ն?D[H)��gұd7���P��ʯZ�R��C�E;)�Q(�z0J���I3��-�>V�W)/~�z3Na:h�ij�T0Ed~�_�2�1��v�\��wϦk��_ϢX��E���mcK0Q�8��4i��h�B����l�l�w�O\%`�1�(k;d�:�@L��|鎹O��uG5wϲ)n,1?Bnwze�~�������[�ZW�i"��30�@HX�9
��ȥ�:���p�Y3T�F�E�ڞ�-��u(ǩ���x1�bS�SVΧ)r���+c^OQD��YDRl�h��䄭�U����u��Ȁ����S%���}��o��l��h��+�׏�4���N�Xv�ch����UdN���)�Q���
�ZJ�yD�ݸS/y�������H��c@�+nƄ�h��2Q��Vt��c��Ce]��U*H�>/G�-�����u�����`©u�r�/\3�Q�*�K͆N��u�K�-�����q��G�e,7���s���G�glg�xv~��t� �W�=dAhu��S���M�f������N��l��E����@�Z�O^�Of�q�ar��]�>�R)s.*1�*BS	W�m5��f����L�̰#���o>��'�
,<H�z���%�/i~E�A\'���WK[���ɋ4�.o;�˕W|z���ap��TZ$���K�*���ک!T*���Jl�%Ik����P�,���2C��UUS]��;���A���ͽ����j��L�}�J�I�-�~��I��glS�4M�o�c�5���P�3>sA=6�;xZT�P
1:Q�3(���c�0�&��z%�I�QgzAY�{W�s��\�V�m|�_�{��8�C�vi��{W��2<0}�/0u��� %f�"��v-N��%IIQ�s̵Ŕ��LT��lחHw�VqR��:������D�J��^���7��\�����r$Y����Z���R��pdM���(�,@�*x�-��>s|I2��V�\/���|?�g9�.(�NK�-�V+�h��>6e�C� ��qk���I1�9Ͱ��ɩ��wb��:��(0���F����o`�;�ף��b�E;|��@m~�6�̾��K�JC�Dv�h�9�eich���g��|]JqN�N.�Xl��.7��Y�����ƕTWnXfP�e����C�l�lķ�j��3�碘(M�&QU���U�i�?y��,�����N�0�2���^��F� �D�>�v�zS�c������VA��kO�J�����RТ5%���y����W����[F�:��t-T��H+��}��A���ڦ�s��ԅ��@ɐ��f`����ר9%��U����bT�k��V��]��d_-�U%_X�>j)�+l�6:���5+]4�C;� W��8A�n_v�  ��!�)�������`�]T�X�c~�-����@����V^/!��r�n�-FJH�m��ȃ�,Y�p���(=p�ub�m>ר�q5��m��`~���Բ�s�g2C�r S1����
���l�b�.�&��Q�QκKM;��	�ej)�����T�p�@k�r>�Pq�7����c�jO����NH%�ƻb&���Qx��F�,�����ёBt�7#�k0�:�������	�������X}���
��r�u���7�e���.g;_�-W m��++`U�H^�"����Qy���3(+&���x�m��%�[	��%�9.��:�\��.�!� +�Tm[�[(ȫ��u:_���Ǉe~��X��(JR��2�}�٨��]-��I[_o�� ڹ�U�r��8�3*��C�\�&���B����N�����Wm��:�EĐb5��#�⇟���#~�(�_:�2�OOv��bK�9�4�F�&LQZ����a �C}�a5)���i�j�r��4��OB�i6��D��YSBu��D�O̹ܜ���+���Y&��2�˷7
Kh'C�+�I�KP��� �=<��T:�ѱչ���٢�5-�!޶��D�+��Y�d���C���D/z���OF�0d�k�dE��R����]�u�V��=-b*���Jv'#6��(%Xť�g�fr�Y�Ǚ��+k����w��K5n��	ۼ^��	lk5qȞ�����k��^8�8����t ��6��j�܄����_�q����,a�lL(���Sh������?�k{Dk�+J��緱w8�'�W��U<4.�Y��+���D[6��N�cbIL�]�''�����i�1j��Y��b�I"������W��R�e��(3��R�1�L��f�M�:AqL#�rD'3\��ؘ��b�}@�4���	����B;H*$+G�qK��왃i�8����E��dV�B6����i��X*�E�F�9���4ӱ],!nCL�z�ef�	S�I��̈5�T�"��Vǹ�t�P�]��3K/Q�.s�� #���x{`<��^��u��_�BB���{���|�����	�I�_�m� )m)ҧU�=��@kC�=�R����%m�K���({������y�hn�nՇ}:�ʟ�(��~�r`���^z���Z��ĩ�sp��㯍823����1�Jc�)2�ܸ#2;X��tSG�e�sKJ�q+u�<��&W� ��b慓)��%Dkﰑ�Z1`',琻^�Z!�/��o��}M�sbH�����Z��7 KXC��Iո��q�mboj#.��*AuU���Ny��� U ���e��:7y�p��M���|.LS̔�c8��M�ڇP\�í�n���+)T���,��$�^9G��\�͸b^6��>��R�,�0�8C�1"ࠔG={qGL�oIkRJ�\&Dos?&� I�Z�}Z�ީ�xj��y�
�v�f�~T�r	�q�����K�&d��o���<�S{�D��S9��|@�؅�uP�nn�GdD{��^���+!&ɡ�2�LEI��� c��>1R�
�s�;�!��������%��ɳK{-�F�Ms��*$8XW��D��H��{�3�B����$����~�c��c�d�.IX���m�^&�`4�O���*�czΠ��ٔ&�ύ�Gk��������I�D#R浕���m7��_/Z�-�^9P�W+�ؕ��P�0����@*�Uk
k+�AT�X�,�em��9b[Or�澴_5�4���P�j����̼�=�Bx��a��[�`�tp��n�\��/<�K�ɚ��)���+`��Zxb��V$޸5F�:�/���";���,҂��|/}��ҫG�[��}������l���U���`�������}�1t��w�.�oǈ�#��@�5׸x�u�? #;��a}Im7 ��uN@���i�W����q����u�i��d�]v�6;p�w~��;7��9Zپ���D�G6�0V�PcSJr��*�ʈ"���q���m��g�2_T��+�{���g8D�vf�����3o���@⥪�\NUZ|]7���g���<���Tռ�3�s���˒n�����&.
Db�%$+U�AW{��	���@�}]������F5ci�W�߈U��S��DX�����R��٣[�I�:탂���^I��=���]R���y�	NkF���u(p\�Lw����b8nˡ;�I�]��"$���.�"�2Oy_>���S]�E�z���v&�,v��@�Q���i(Sj���UP�&1@t�������ޙ,���NO��lelVLs�sh��t[|cv[�46��Q����C���2'�$��_>�V����'>� ��������ۢ��������@Uϒ����y*j�!%�������y��Y=e��WH�+Ud +�3_�����L8>�(ș[5[�F��Y� g�(������1���GO���7��X�q�֊�����|{�<�B@���������ãϰ_o8���5�C��%���?��7cV&JV�+��#��ۑ�	�ðVK��/�}6�[)p�1!�������^�[$Q�=�m���|kq�F�]6�Mk̏ O�3�S��P����wid�cY7������{���/+�J��~�v�Y�}�ր�Qb�8S�*� ɇ� UqsG�=�Xvy��O�'�q�����&n0Z	�\1GPZ���t�6;���*���`�E��������=j�}�g2ɛ�:>��� ��ebޅ
���Vvr��g YϹ��½j�6�UHNpG�C�ű>\b_��U��.
�0�g�q�B4Rn��`Ц33��M3���$C�i�O�(k�����k�,��ڷ��}(��M�n�d|K���3��Y�Q=�%�w/���WP�8R�7��-w�DT:�em�j�;��l���}�o����i�O��7oG��̬>�َJ���i�Q�T�:W#��a�tm�,�$R��弄ςG���?<�b�"�B ��,�;��Ś�tY<3��OS� �\�G9g��Ӻ&Ca���n�3�M6<?�H�Q+S�<����y[�,��,W����~���I�s�h+��_�}E�JzR�U�H�/��g�	�&h>���k#v�IU�lx�g�@K�H7��S�o_���t�^�,���=�Y!=E��/���!�~V���r苉2��Ƃ[�[�$)Ϻ��Hh@_��C��hP�����Ztn����ͦ��Q��ȕH^��R_��%}��a�g(�ܩ��S�����Z�l�@�w����#z��(�!�Wō?�� {k��HϘ���o�|�W���W�	ܙ.�Pވ7�?�����#h��ۑ�1%!N[�<�)��5��U��<��u�Ĥ{7-8Is�/�°~YGDHrR>��5�ǋ|�I��%Q:�X`:�_Lt���y�������ze����ᘃ6��ߗ{45%����>|�8�A�Rڝ�����di���;<�h�Z�¾����
�Y��p��+�z���#�^uE�D�4Z���T����x�����;�tG���S�<�W��K��F*Tl��cF+�P�u�l9x	�8S�c���y	9z" ��N���fw'Zy�!��tNn+��B����H?��I`����IMm��<B���^�ۀ��z\��_�i����\a=,�W7���������6O��J:&�?�hba�� ��f�ϳe+�Ib�Am���S�/�r{��3e��I\�˨�.R�>��:*!gyȞ��a���D��sU�[e~NXZ)A��y���=r9��K���<� ���v��-a����a�c3�UĥZ�79ڌa�w'���>�A���p��T���+���<¤σ5JxU����3���h�Wk-�/�,�'�H�-�Y�N�������$i�?���/�+�y�j�7M��8��4//LԠ�p����!ӻѯ�V�;B��R�ȱ�L��m�S?r໳k�\'���k9b�y}i.��*�U~�M�u�x�% N�6����Vf�keS��Ͽ�)grax�Q�������QM��u�֞ȅ6���?�J�cf��{�0��!��J��	�I/dP�'�FkcԪn�cV΍����9�R�^��N§��Y��, ����u����a^��=�a�F5k��[ �kf�27�;�j�'j�q��k	f�b��]��	?�6hB�&�<������[~��)4���]�n�f�h6�>�R,@��V�Ѹ��>��ټe��$�0���Sf����ɼ�EJ���qJ� и�uѬT��Eo'�[�ICYC0�Ζ�3\�u0o�E��4����['�M�D
�M�lEy��n7�Hi����}?��\�b�|H�jc�����`K'��?�Or��X���>�a�p���	5��c@��Z�G!}��쬟��B0?���Ao��Xl��ű(�8�V�ޤ�m�:�����@���K�e3��
���u�?MʷC ۝O~w�8�AG�7׽�V	��Cg(T8�!�~��4]w(G�!�i���
�����X{��a?vuQC3�
�PDs� J057�yL�����N��}�n@����j��0C��.Y$w�!�NikpF����=��z��UO����(�Y��D���n�u{�n�����쯻�\p�T
v:#.�fԌ癏���&5�c��)}���������ɳ=�E�DH�����<肨����=v�*�B��֛��F'��~��'H\�K��g�	���� $QXR��u�3�C'�I�>y��N��&) �pn���(2웄Sܓ�An|Xf��}�9��@*�ȰQ�i*ď k�>�������Li�^f4�f�WA��9a=u�lo��ǅ�ѹ�	�;K��,�8�Wь���w[�3<�ۑ'��ί[U�`ďo�h��U����h!6z�o��0>��*V��*�(���U ݗ��'��Xnx���j,�Dq��g�t�&����Ԁ�Ǜ%^�w+�/������yp�9f߃�1k���J�^9����!	b���\c��-~৮\�D֚���(6Sƒzc�ʚ�J��	؅��4�z���e�K�E����2�$x���������H��O@=L;S�+H ��Z��6�+�D���+�� �M��<��� ������g5�=��dX6y��dv�R~e�Q�ld"�YGS��/N�P!	�!"�#E㋣p<jw��1R��xW��嬰�v����
,E)�ik�T�A˻�)�e��ҹ�g)�[��?Ͷx=]�W���O�f	�̤B>�~�I8S��i~��ZM�FY�آSR�I�:��q���A}k��Ѵ�C1/w��|�W;n��@Qh�9��X���3�.�U��ݚ|��6�a�=�㟮+H���D�o��}%��}�
K:�Y+(\���*���4ws"��)H��DI�w�
d BQ�
=\���d D�[�nK�� lh�w����Z�Z������J�[e���e�xӒ���[�3{�ڃ�?,�.�'�]�9c��iZTɑU�RS">3��O��U,���ʪ�=���3�当�d.���T�ʢƻf��G�P�c	 e�m��z��M�/m�d�H4���R�g�h��%,�t��66����Yb�pQ���é')w��}=��Q�?q捙f`:����@>�Ϟ�8��D7ɴ�΁q�=��g����e\v�$�y�w�<�:�n4�ㇾ�~jf���j�h���\�ԏ��ߦ�,�3�Ǵ��˾>��J��K@��})'�B��!�E̴��!�i��/�����y�wN��0B �}o���B�0W����?X]�l���axf~8�����+��ˏ#�v,��75%R��\��g�TZ`�I=��j	*����Y��VA,I�-^�GK��K���:2��Un��Y���jT=(T�d�"�;�S��P���G�_J���=44MxO�c�Wp �&�%�S��'�Ͼ($!�^�ڪL��g����"O��> �G��ч�/�<("�8�z S@D)��V���4[['�^/���;�i[������"��f�HD[�L{r|`5�'6�����Q�����j��i��* ��\3]�}TPw�2��R��{��(w� ������>��]����	�a񆾩WA�۲�l��$�A�Ԏ�yF5����t�wy�N(�_b�v����B{�`&&�X]��Z���r9oW�)ƽ��(RY�^iu�4����@s�=�_�ix}c��No;�8���^��R�oܾ�p*�̹0tq�=)���	Ͳ��N!/�6���I5`]��):���� �9��8���#��D9q�4=3�?��,���G2�@����EV&r�	n���5�a���t:ZR�/�J��'��I-�O����2��
3�A����h
�mk���/U6(�������#�\�.��4�e��N����ƛ�f�:������E�7��R΁j��G�~�ƽ��3b3D��vM ��xi���6BnΦ�+���^��F)}6Q��œe�[���dY{g�6˂4s#>C�&��F�;+�q�,�_~�9��$�⧡���~�oԬ�(ky����9�oE�=��G{���Ǭ�����~���N<6U���Y�3 ��=[��Bg�%��¬s$��:��^�gj�*9z�qX��jGܘ�4��+g��d�F����*+���~6N���}'���Z���7�(� ��J��-O����p��	�prq"˴[:��Иݒ��!�k7�������m�XK�S������c @�毦�H���r���]eZGZP��2����W��04�.��e|�4W6^QB��6o��bn�����4��4ح@}�%����Q~���Mi�N�(�g~C��@a�X��S���AE���5x˕���9�������Ɖ_��b���Q/
� ,`�*���������]��%�o�I�\�:�iϻt1�B�GqC����w>.�
V����-�H������^������Vb���-F����KW�S�+~��)y$#5�,����ss�͍!��v7��L���"W/Y��3������x^Dtφ��TT�\�akb��[��B8�LVƠ|��)��v~�e��C�T����l'`����Ί��`��r	�C}�����늱����T�j��|^Md`�V���h��c�Ĭ�Q���B��0�T�Մ)��|P����y�$�� k��&(�"�.o����V��KSG�fM/�[�WB M��V`=�h?@�{�L�_���9[�aƍ+��i��
����}�
�c;�s.}O���.�P��'������`EѰ?��*��d��n����>Pn냗�n.{��,�ɍ9u��K�3�� ѷ߯��T��Ie�2_s�����/�q��ڎd�R_��g�>�3�����Ը�A�aqe���1�N��"����Ȗ��0������l�Z	����&t��}|/*EIr�k;)���(�G���r��	�l�>�:T�%�S�>�N19�c�/r#K3��v��쮦H�˟H�*�'�������ܹP��G-ֲC# ��t[�Ƀ���rP�'��h(Kϙ9�7!S]��^��E溆C^���t|R'�;>J��A]F���P�X�>[1�8��=�o��p-�v�,�%@ql��S0�z�x��px�ﷆ��h �K,��R������(���*8���z�6'��Jx��JBt�tj1ߞ�Jw;K�����m\j�7�D4l	V�:�-�ȪXH��F�]���V�!3�a7I6K- :%�R��u�#��:\���Hc'��I�l%�e�$���0���i4t�y�Pq��+�\*o�a�[EW�	}����@�Zj��up�S2C5K_[eP {�N<Qc 6��
b�r�!o)�t&N���:�����Yqx�l�5�Q
V����w�|����7�`�����T��q���7RהΫ�E��X����w��C�w�NzGv鍒���o5��K�+�>2' �r1��H����"��lD5��{�f�s�n+�)�B;϶Y(�=�����B��h�l9�ྀ��}8T̠���-g�d���駆�a��X�i�<�M��E�U$�)]��T��h��q��{����I���a�V����@�B��~o��#y��f �r�5\f�c	��쁩��R,��]�g��������!j-?�{�XY��A!{K��.Q11&�D�����b<��j�ì�N�8�H�O���8��p��Q�p¼o|�X��ZW|��d �-�O�%bBP.��V����wS�7��
���F;����!��L<=N�_G�� 3�����L��7c+_���p�}}�*7^N�p�����	^젝�/�k�
��u���!͌ds��ܖs�T@b�f�nz�u�Yy�j*>j*V��rao��'Ȏuk��+6�m;Re�q�p����$rT�aӴ�Џp�,��0,�ɼ�� 7^�4,s�R=�Sns�� �kw[Ԗ��Ƴm]C�%�>~z����Vh׆���Ȏ�9,m�B<W0��M�/�����̢�rw�+��z(�sQ#hX�-m��yX�FZ�����jD�Wz�L�*^VWw�D���fH"�Y�c(��}���w�:x�M.�C)P6B3�%,�ԍ��CC#!	N� �����~�J�C�aj!����Zx��"��7���Åǡ!	gJ�Z�I���7�-��$��
O|'�����y����e����w���ƃ�>@���#x�ї�L9��=�J�+@gA���*�kÀJ�a\�P�pwҳ���Y��8�5�E�@�b��g��쫹�ω�8���./�F��� �Y��t�2�m�������~��y.<��p�I����χQ�_��TSxZ�tm.1{J��M���O]
���қ��A��C��s��4�i}������@��Ol�=�D��ߥMYS���[3%��C`�*7�v��xY�~pA_%���|Ӳ���[h2�V�uW�&��(=[�yhXؽ�,26� �<���Ƴn����
��m��*ښH2?�'>
�o�w����Ff�߫b1�d����Lt.��F����e���b���Y�7]$���8�N"`�_����ݒ��yU}H�]q�.��?FIe*��/A�f�uִ�F�9���hh�\c�K�,��AJz�:��������ί�;P��a����s��\�䧜屽��G(��`����RhF��w�C��>n��Z�X�`�Z,��s�b��cvM?H�g_m�>�>w�n;tֻ��ӱ�ʒm��H=ҫ`���Ddb��<�h�����!����h�&�!y��-�	��q�>|���˳���U�R��t ���}[G�{_k#�f�@����Q`ȈxD��֪&{4Pe�p��ͨ��m!��R�5@`$�1Zq�$��=�Np�y5�Ea�v�@�5m`����W��]���j���X�VY\#r�b�78Ha�m�,�v��B� �0I�������Ʈ���ӊ�E�d�"0�q���!�e �O��4C!��\K��U���[��~���I��h�0���!�u����e:Ds}�L:��~7�P�f�(M������.[p�^a��[��p S�[(Ƶ2���Ӭ���6I���I�w���1q �%Jaj%�8[��}�
����]}�dx@a�U`�����$n�P��+U-~��G3d��%�X}����$fPm{ik��E�9âB�r��.�4Bġ��E��#9�~ U��?�YW�1�C�U��w�鋲�,��Dհ�<yI��⸟!�xؿk��b�RtR��%E���:V��vV AO�׀�caM�"p�w��`�3qjY�+(sXڸ��me��zl�]J���N����>V�,�>��K��D���V�ph��p�����-���Kj�J�K-�	)�uU�tJ/�\mWj~��c�~������Ժ*��9E�&H�x]�4�N��Ur�n4�G���c�(�G'���W�f�+{�=0'�F��$�ҾXl�Ȱ�#���u�н�,�tsxb�������<f,�}x�E���F6R�k��0�ٳjz��=�����e�D@L�Kq��4E�1��3b�����y1-�ʏq�OA$lH�s|�Y��DE�O���v�Ӏ�����x��Gm�XZ�UOA |�$2�7�r�z��2��:MC����JN�Z��پ�� ǀǰ���^�o2�L�k+Sa�~8�w��/�&���:���l���y����)�<�ժ��~�\H����A
9�X)��ώ�v�W]�̯q�)��1 ���!�m����W��A�&إ��V�˖��8��Z�9��a��Ъ9�_i�?m����� �HFkX�!���ST�--���0�[4��L�6NR憩2#q\o@�5�����P0�P��̖��c,Q���H��J�[m�M�����w-����0C��62��q�T��X��e6G�l����%
�O�	���qҖ�X��cʶ��˦ �q��6sS6�b��s���Ns���,�����j�'��j
�ko.MV9�n� �V��C� �ڈS��?Ӻa��)@��5�kކ��j��ϛ*�:53��sy���~�9�S�EꖽQ�*%��
g�P\׉4Ky���4�L�	��P���UJJ���� �BP������r]�:V�=&zא�$�B�F�+�T	w���`���HW��)n>",���FSR�O}�<6��uL� Ŧ<�7J�]�t�7,YXs�hb�+T�-t�O����k�Wko�4�`���K^.�W�g{���.[����|mpK�܉�3��Q�xq�nĂ�7A�C��H�i��M�ee'�:���J_��ɯ~B$��d45$q�Q8��3p�R~�D2I�If�,�9�b&�[����q����Gө�sc��@}��SYƾ����n�I���Oz�(G�|E";��ϯ۲��%�U^����7Hf�l�|6�f�2�ڦ��?�^z6G�i�H��_H�m�	��$�~&�����aMm���< q�ٜo�}O���19Z2kc�u �x͢g���m֏�<�>����`��EH� ���u�쎺]{i�x<�������=��/��Zb�Br����r��V4HN��U������2۷0����*�!�\u�&���RF�o ��+xy��$�'o_��Ǘ3�U
k'��W�~�;��&j�����#�r8����J�݅���!jX1t�W��>��Riir������m
�����[WD���LM�����r�C>��ݙa\(�Tg'Io4�3]#a�3���6}���?�is_��ӵ�&5�Q��gZ=O����������Ŝg���k�o<����X�-yṰ�R�%�ƈ�e냻gl>��N�/#������m�8�LK�G���z��^��E�~�YA4��?A�E"���\�.�������s��̔3-Wz�A�3��@�#1������*�E���	�"��vI���X~��:����Z�}�����^6V��c���o�*�WL��.d��Y_��G{D��jS�� l%�^V(;�ŷR�Ǡ��aXӀ��R�-Α�1G� 4��F���*1O�"�Z�����F��p�+f߱�H�F�7m��Ѵ����U�?�+New��|NJB��?üئ)4�ӽ��򲺼�*����o�S8ռ�Gl����[��08��si��Ӂ����ʥ�ˣb�.�ܹ�{�[�y3�j���!G=�ü1�i{��X�16��9��L���S8���"��N�/#G� �H#h���9����O��P4u}.89Ie s>&�	H��I��bCΘ?F��.	)��l��FT��G��"��5�E�_yVwsUOg����9�R�}������g�����Ix�v'���0d-d�4��g̜����)�Ĕ&ud2K$q9m6�*q��OOOM܇#���)�)�gȲ�<#�ݝkxE��Z�NL��w�T�f�?��rw!����4�ۘ���c{8G׵v�8T����Г�۴l�� ����6B0��X�-�j]"vg��N�jOe'�O�Bg��@�څ�yX7�<$eoJV[>~/��xJ{2o5=�F��u��:�K�_�^�����ɀAN�ņȒ��9�n�­�j��'&B)�l�T��Th�;)r\x(��5�V|�����CV
A,�o�m��g�
H����׶�[K�)�`�r�t������y��0Hw7�v��_JV�)�t�j:#��-��QC`��Ok[J�~,��,���u;�V(\��� f�r�k<��� Qz���i�gX�ۃ��ѝ�j�l�iR@F+?q�?������$���G}�G��`�Gw�q�<�G=�gɣ��8$�K���
�V�P����
p�T��O`�@�4�o��Ԇ��L�\�*le���C��j��R���$�2F$���='gv�f �'~�r]����@i��[-Ͼ<�cs#Z�ʁdm+P_f�U�l���3����e��~s�1�{!�y��l�ӟ@k&O5����(�s&>�"�W��Q�U_0 ���V�RA�����%�/��31�^+0ԉ{��\�?�iҋC(�J�����AUJ�Ұ���~2����$�A��ȑ7�}�x��l��/)��Sn_}�X��3ɩ�\�v����(��T�k�W�1+d��S��Pd�ݙ�2�J��zu�JSj���\�5w�n)�E�`Տ?�Ui�*_�0�5k��U�	���i��KƝ�}�-��*,�ֺ���������K���%F�H�ɪ.`R B��X��	f����`���s3�H� 'l2���x~B�}�����ʔ~W�cLT��~��)Ta�ZV�Vfϱ^�E�A��V�Q�L̓*^:�HL���p�#RHY������+��=�'Q&N��$E^�Q�Ovz��R*N+�d������xό�	4�2������4k�����m�����9�-xz�"@io7�Z��>�>wG{��v�ͳ��N5?Ѓ:��q3�Z�h�azB�Z�C5O�Bn����������5�����:/!D��L�P���L/7*�/��x����}]1H�Ǩ�[�i��8ChNMCW}�'[F#O`YL1M��B�2W/�]%��C P�]���j�c�y��^_�EX6}�2�u�PP�:	`d���!:��L<Mֹ�v�*�g�c�(4>�����9�O��5(�S�D�:�5;.��DY�t&(NTV�08��qQ�jK&_�9s�>O��»hW�ƾQ�K_et����(���!��=�JeP"x-"�/|��#���q�� ��b.#�y@����X_`ݐ�8����js�鷞�'��x�]l�\ޜ"M�	��a�T5bX�����T_��Y���}�� V��iT�s�i�|㔏i����^n'KB��x]bÜ����=T��܎7�V����Q�Mցn2���ԟ�㇌�{�x�e+c��v�qu�W�}�����om����+9��J��Cg+�y�D�b��󓬄�"Xa0]8_�\Bv�"6J�E
�M^�Ɓ�8�G<g�t�}�2,�2)�����~�~�X@N��VG�2��r6�ܾW�; ޝ��MEk��Y_2o]���JŤ�3\�(=f��8`�a��ƘRU�����Øp���䀰[�<�M��������o+���[�nCj��H�;�/�b%�׭Y�qP�o�潍�8��(��y��q'c��3��kf9�.��t���>.��$5t�n���!�8$�΄f3e� ��X\����n����B��iK'0}��ry���y��N۴cE��H}�ޕJ�
��&9M�Y�j5��8�p��9R� �o�f���͢\)��e0�ӅL ���˽�y?�`o�d�Ҳt�2'��-���i�jPǰ�����2P:1�$�{%�p�9�y�&{�;�DF��q?0a�;J�Sdi.fT���i�8r�:��U��� ��֥�YUg���ӍX�����w�׿7��=l��kOp����hU:�~H ��~�>tR�{�f(8J���h�	�@p�l�w�b=�͘�K�&}P�#�p�#_�̬�X���e�[�&ؾKA���{������,z�̼�榐.9Ʉ���Y�[�q���,p���3�	YF�U3�풦#��d#�B˟��unJY1,z�O`�pg�"����i��<�k8�����% �����.��
����i�o�ã�*\g5���F���������Pyi0�5�:��d_}^�259;o�f��1��e݆ɠ^�X1�fY�o_E1VVG�Q��6��0uS����Nk7^s#2*=<�끞S�Ac��o�?��hDu���uF�
��C�B������ĔK�ŧ�dS�R|���[������S��Ⱍ�/0�3w��-X�ܢP�L��,ɼY�jBF��6���NΝ7!µA��+�LS�D�X#�ǎ�[c��*��gz�&�E��n�
�Z���й9|�7�}(�(���k�S2Cf�O��6����"�T�N�X���Q���#;t������q}�-�x���T�Y��:���P�ۊ�F�|
�RĆy��`E{�t4���B�-Ռ>$�E�B�����࡛�!W܉oJ᧕̓�c;�h,�\��r��lB<�rKL��\���ߨL5�C��Hݖ��.����F�?\��܇�ݨ�%�{���0����� ���Ѣ�Y	&Z��g��������S��6i{�/���|9�xl餤C&s%#߳o�z�aQ΋�b:�؞�f�mށ=��b<7f9�HK���R[/u�l�LZ����
P��Ss��JC �h3�Ҏ�H��F�b�p-�K��Ju(e�a�S`�`h�%/b"�t-+H8v>�Z�-ae7e0Na�q��w�O�k4趒�\��q9lT�8r���:�c��ȁ��'���	�i˳iZ�c���ޯ�-0,܈� o�d�pNR�	?�EZ���\�+�7t(D�Jܝ-k4�ۡ9w}̉i�7�z�M��+#�m.���ee����ds�e��6B��۴����ӗV�K��<�Ó����ܺ�~�V�	�j	���i���"Zb]���\x[O�`vS����aٻp�a0��=� Ȍ����ߵ��'��K'��ea���?r�m E�
Op��5!Ztp8	��_��̚&��@o,*�=)љ�	���E�T�����V�넷��%@�d&R̓�I��Z�3:����)q}�����{�q���d]�y����jn�R�0\��*��	��մ���Y�A��%뢱���,����Տ㙪eE��e@�ĝ�����������6��-��Qm�����y�W�GAi�#�|nZ�S�������>��k�S��|���V�ȸ9�H�:��m��4Hm�[���+�k�+��RQ�h���x�.� >&�;?�)ˁp�]�L^$�O<�w��Al����4[�e?���֭��H_ƿ'����<�j�&�9�Շ�ԛ�V!/��<\ڋ��=��>�������Ջ��C�䕳�0��0���jj�e]�Rf"#���R�xݬ�+����vi6�
S�������V���9�]
(������?�fDk��7a�;BQ��d@q���i<]�=����1�5�8x��Cs0�0$�B����������ga�7_�EaP���;E������:����@7�U��������1�{7i�U�.Љ��?�)��׫h=W	���yǑF��=�w���(ܲco�vԽ8 ���nP!��s-9�aǀ=#�Qm�������3w�pL���q��s8��<:o�Ó�7䚂>�����[�7��l���BH��_B����:t����1�g{7���JDv�4�����pЍ�|����0���[W��5;�+�zwB�� �.�����7�D�8RK=7�%��QE�W��lN�5}	/�-у[���>��$�D�F�W���뜡���<��+��%҄��~]��cb��>J�!������[d����w�k1���t��3���FE?�thoS:������-���E��r�>�i0�����;�L0�3L�{�ðe2i�޻�8���Qj�轾5�B�məMd�֋9�9W.s;�>n�3P��C�)nQa�XY�+�!��P? �3�%A�ޯ2��l�9��q�������ݻ\Z9=K��2?����_Y0b�̲RgIB�&�2�}O��ȗ{��%�㞣u7!TS}�$����ne�
[�`��Dn|���AF�>�1��qȴ��S���v��=᯻/�'�hf�]���}J�"�vj\�����2g�p\ց����S[�k9�����ҷ'9��	#�n�>�Q�����weٰ4�s��AT�)�� ��>#��SuIٿ�
���)����}�@7�Y���Q�/����%�H�H$�}����å!(�6�6�����S0��<��ؖ\X=F���øJ���8K�M����9�Yr��,9�9̗f����(�+�`��4O&"ݹօκ�����N��>�C����S�,c��C��3���+}��t�C5��g�6פ:����=��D�e�h��o#��a� �s����1n�)�l򓽗 [����>�����J�M�W�l1�ѭ�o��n�#�K5j\1YH���!^����YM��n��70�Ԫ����FW�s���)���G��#��.<����+�E�+	}�4NG�R��jmV�T4~�r��:N2W�ӏn��i}ؒ�*z�����`�'�����L�%���T�8��7S�B�@r���wN�0�(5b�?����i�Z�Ӹ�^-��sPA,���~�C"A2��Kj�8��H��A����hm�B���{�+�?��.����n�K�|T"��V����2�� �7�(x�QQ�lD 2br�(P�a�i��+�d�h�IG���I� ]�u�O�c�-�c���ݴ��G���\j��X;�ʏ�����E���1&��b�WW�l�~����]��
��ZE��]sX���A�~4���g�Rks듧�`�_в{yv~��\`ʑ�c��.C=�t�D?.�~��6�2���\�Fa�_�6�u�l#��oq-�����nn_H>����@��Y�~�����������3�Ґ�U�t��A��h ��p�rB�D�SD�ZP���/PV:t8F�d�,��~��q�<�EW����*��]P.�Ym��1��i����G�S���#�	v��vi�R�jm�ʫuw��)w�Z)Ȼ+T�����,�J�v��KQu3�Z�K��|�d~q��X	
7����Db����� � YF��4�<:2�x�X�+�(�����|� �)�I��` #�W�,X=	����R����44"k��'gS���h�o�/D�{V�	��n:�l���If�/[���o3�{ea#�,�u�`��u��'����'��S�5g\ChX����T&�}9�,�;����%�P�髥ԟ���r���t���+�^T����KX)nOx��M��{�ϘI,����	��A� ����h��]	���Qz�(xE0�e��V�@0�`R|D��^���g���p�V��K�[��j��5�4�!8��X�TMx�Q9��)c,7+\ϬU��H����.Q�H)��K�U��c-{���J�{��H��иe'g�fi�n5SI�����9wذ�qxr��B�}�z۸��m�N)f�����B�ހ�)�ew���5�����/�ܗ�a���%�$�1fa��mf-�Uh������I��9�SЩ2+J���&�)/��!���j<�Z�uꏈ�f���YL�pƻ��VL�ډ��zǳ2?�E�2��Q�^�E�d�f�/+�(��3�<Kө���m�8����n �����8����iӋg��6X1�DM�+eW:n��̲uJ��]�Ca`�_n$W:~��8�K	�H(��FO��?l8�d��o��O���'�cڅ��]��+��碇����ƥ3��kBv��
 �bޑ�,寠f�u�6�(Oکw��k��Y�^��2��p����/*#�g��dz��%��Å3�|��[A&�[�K�G̵;:]ct@"��fLdHM��[ͫ�W֟8��v#&#WD��YJ����EYl�W����ҧ��������i%	��)�H�ɣ���6�+��W�V;�O��؟@\Fp�R��g����YV�LK.紿�ZeQ���{gIWW�T���X���g�syj�eX?��z���D��@7s����zeJq�&��)��:i%���p�ǫ��C�IV�2���O`�Vj��`��J�mR.%0o�j1�O^f��C7� �?�/�C�ni\Mg���~Ew��܈��;'|�t���K:J@kj?w��Zk�H`&ߚ�
�B$���;�g_\�X�FaA2���l���*f��:f�g�A;ͅ}4�x��(�����	������i���E�ā�z��$�N�6+!�!u(S�������q�'�99=?%Qf	�:���D�f�cZO��.F|N\����i�AX��ZC� �u���"�����tv�+?���q�c˚��繅g����
!t՞��F�>�?�$ �����#�RR}���fyToH�
�:+��,�-A��U,yw�V�Ȣ������'�|g���AA��_Q�ɘ�)&{�^D���ޫCmGa��@��e�C�ܟ�1%L(��@���b<DjO�Ɛ>ܻ�US�n���<��5 �T�\ ��_z��	�`JK�h˯S�W��N�0<xK�J�&e��t����Q��p�*
e�+u`���#f��ne��f*�N<���7qx8�Ib|zd�'�=�es��R}��o]���U��\1G�2oQ���p>HOo,��Cojx�Hx�b���H�Ī�D0�� � �8�1)�&��l?-'����rW6YѴ����R�UP�}��N��Si�࣌C�z��Zk���i�?��<����|6�n���'�5�����ά��VXB�q��/��0�Q&E��z���·!�m��(��UdHp�b�zX�t��pE-����1�gJ�W�0[�J,9Z.��i��H�P8t���Ƃ�[W�~1���F�/3�Jj���\c��=.Bk&�?���/�i�5�,W��?����_|���`���Y��&?�2�z4qT���|.��
�9!EF�@��-ذ�Pl?�q�1�Q��D� ��x)_{�������N�o�KD��=��6�@��ky�ʪ�@l��(n�����2N��awC�� ��w�f�A��ȿ��xo%/��{����{Z`��[���!���SE/����8x�>�;,�pv�J�咖�����dC�{"�`�
��0�v�L���E�d�[Դ��}�F�nZ�s3v,�U�S"q>�}��6�Dݾqw3I)����S|(�bP��y��*g}+x����$��A�2]��!�d�p3§����R#���1d8�׋�]�����?��0���""� t�ӓH��D�,��n��r��a�?�M��d#�^=pTt���u���+�� �h��yC	����,�T>�
Y�o:�)��-V�3|���;��B!~�E�%�ؔG`pf%@��{�fx>��L?�h��4EQ�$K��Ozߩ�~1wS��� P������P����('Lφ �r�k��c]9l�%Z���MK�Dړl���e�ly���׋'��Mc\&�Iw��h�r��R�����s����^p!ˡ:�����߄��L��lj����ip��*k#��3� $�LA�C�������Y����uз"<�pE��tc��ں��Q��U�k�=��P�RY�U�}p��4�������1ռ��~w�OO֦�}��ڿ��T���|<��D�qb���Y�ĉ�+Ҹs��\�z#� Z�����|P���S���J��.A�5�q�MѮtN�&�&_��ONPk��F۬Z�Ҍ /���BPA�L��hPM:3�H/�lj�XRd9F����t�V�"���A��Ish<^�i�t�]��$���ǟ	_�V�9N1��_?�B�@�ְ�5���{Y"�R���^�M8��O�Ν:�x����*�XL-�5D5sG��ص��JI	\�bY1��u!��qV��9��=�2?/>P�HB�vBա���9��V�J ��b�i{���D.
��6S�������RY�ߎ��ZxW5�j�d�=�@���Gb\�)�b�	9���3�oY�$�TG��M ƣqӿl_oS���s���x�����g9(�B��L��u��D�b1���8���9B"Z�|ؘ�Z ����Ao��3�D�D��S��Y@�A�θ��T>#  �/K"�%��������j�xy�_sɟ�6K��D|��N��3:Z@�}��s&�nE���b�Da��
1 *�� �-��a\V�7��:�=>T>�*B��%$�(�sx��)j�����i_��^�2������J�Ʈ���L�R�n]��7Dc㑠�n!����p�<�z41�!�j/�tÅZs����:E� ��U |�3胶_��� ��C�&{�v׵0v͢O2z\@0w� ̴�' ��ܗ~�6
���E�\���N�[aAS�%�x��L������je�H���W�m0?%��=�"�
�I&
H0�KřG�ܹ�g*�+H�4���+��pfe�Jc�8h��O����s}�~V��\�pi@��9�%�K�ц����TP�nw�w9t�<��Ӂ�,�[U����0�j�x�ar�:*@C�5hn=�j4��F2�#����Y�����ءMZ��%5��1oo	n��Q��˲x}����DBX�B|��\��[���ITU�3�:�sY5��/�$���{Kl�.�-�9�*���g���Ct�l�O�C	��PY���^�z-�D�ne���LQ\	jGZ���i����
�h|=&�3����;=�{���l�O��x�(��`F]��f��X���؏�Dy�E��YFC�i �7xC�8&���cY)E�XJ���d��>���[zV��W"��`'Ŧ)�E������}�4�֪5;�؊P�vp#Xbd��R�+����G�.��<�G����0�^M��>"ulH��(͟u�D�\
[o���D���$�����T�>��{�4E�/I��3�4��Oǡ��G��"PG�7H��t[u��.��
V�s[��T�e?��L�y�gb����gS?0b��'T�}�-��H���A�6��w�[�l>�P���ȧ�@=��6�n,UK������5��\��ed�M�w0G���nQ�r��~���`�-/ٽ�6��>5H�U`0�%q�I*��(Nb_28�t�l-�9Gm퐤:��1qi�x�E;W����"�ɿ� k2�z��[q�'q|�u���{��\D��%e�y�M�Li�.�9��F�[�ݪ�FR)�W��v��}��g�IJk��Z�,�{���IoV�s|k���1��А�L(Ӝ:��"|���F.Ҫ
�8��d�v�Oѱ��@��~n8ܚ5�N���J5�_��_s|��g+0����R�~s*��-���?��B�����'L��?\ ���g�3/kX�F*� ӎ졆��*(O?m��F�I��;�TK����(�`	up(,��>bDm���CMr	�q��Ҵ�8����i|�Fvx#����� �u�#؞���l"cD����(���b�3�B.��#d����,35�N�ee/�H܅I8YƫY˃���Pm���ْ����a�U�`}7�Rt�h�t�]KƢS���Z]�uEӚXэ�9k6�|N�6���+��ʥ�͊����GbԞ�[��p����W +�o�e��8��5~���h���:܅��XB����Maf���zw�q�F��V��`b9���i'b��w��sZ�&�R�s�6��h�S�5{�>/�B9�8w^���W̸�?q����W���U�v�e����:x�ϴ3�A���{��y厁Dbv_��ݒj�8�N��|�S��f ��"���@���2�pzЭwa�%}�)\�)�{}?"��PԄN|��h�M<�3��spneJb���ҥ1�-ZNe�cNU����##��0Wߴ�u�%�s�rm��V^�)?�����fm[,�%� �Nib�Ϧ�xߏ�c��uX������Dv�y��F3�6UJy��w�Y�(�F!l��>=���/;UX�zA�G�fa%
*�7N� �U�jޛ�é�M}���;b�d1�l���E��̋O�f�3�r��,�7�@4H�M����#����x��n�����$�S�(6�!���_Rt4P�0R��_4�J����A	bj�Q.`���=Þ3�K�9$,Fc��������H��ɲI��W�!��.]�� X�8_S0����{:sv$Qz�>�z���и(���b�%ѷt�*Yz����1l:��I7eKP��B�@g� ;{��~hD.�̥�G��а��|�7��!�<�W�UB�f�ǭ9 ��(���]��&���V���e�ٕ�JY�[5x����Ֆ��hx��5����Co���<�q�$������0�z�PG9^c k�\~紉�徥�j�!�����wތh��HF�I�,���B� �d��r�O����5�b;�ⴥCJ̼'�X���	j��`qF���<�V���48`M��������?��m�e�Ҙv!k��D�5HH�����
'���1Z�Ò������pm���1����(��m�]��<��[ ��N�ɾ%)p��.(��3�a��E�W6���(;0�(c��\�M�4�?��.C硬nZG����c��@!�O�,������D��L[�'�C��p���;m�]8��#d�T�'+�4F"���)]uL+�;�y$8-�T�G;C�����ѻ�!L�x��
�jR3��V�W&GT��qR��4,u���D,��� �\޴4��5
��|%v;~�b@�G�oS4�ĵ^��K�5��E��7�w�A�NÍ��6�!՟��<���4���z��M��G*��U�u���v=q��8^��JXZG�bf�+�#�I�p���e�J���5}��� L�uHV�#�gr�	d�8w��G\p���?�;{���C2�.���L\�.�NMS#�]��,�j7�l��*�F�2�r��	�5��K�3���F�L��n�t��!���x�O=+K0+"ۢh�1i@*�p暶��@OB�@;-qN{�j����vqBH�w���C��6hK�~-=
�:�_��Z�s�.>����joO���5�}�+�U�ע�8(�ә[�:5[�+���	�ʴ`�w/��W�/�Dt��֡�;b��2��˟��14T*HĖM���H�ݯ��1/ުs�0QD7;͛���>(9�<�5�|�K�.�ډ�۰�+M�n]}�~��� �}*ʄ��H�Icoًt��U�\%L��Wn*�l�lt}kA2M�e���tT0� LB�}m�zIx{�J2��j)�-R��Ɋ|sDW�� � �?(�`+i�J���**N様�.8u �B����i�Ĭ<frS�W[4�Ʉ̐1���4��hFq�� ^t���I���/�d9��'���,<���z>�`��d{�6�\���M�"����! U�ܻP\fO�	�sR����NPA�uT�0�u�&B� �����\I�KX0��4�6p����B7�^ᤧ!i�U��BP�D쟏��Q1��m/�,fCY6��P�x�� sa�Tt8��WF��}��Y�;�����\��;�RE9
�uT�#���gp�ܯ���y�2n�:��W�I�2��t;��k��D}�k!�:��y�tL��͝�yƳNkh�Ӷs܎ō'�~	mMf�QsL}T"a��r�����v(f�f��}%��^�ܮd�i��hd(�[ܓN0����ѯ	h˄}���09!ug��D<���z4���4QF�B�7��n ��><Th�� ꦟ�<+S��?��,�J��D����['�f̈́��tǲ+A�?Ʌ�Ʀ��k����"����j�W��w�\�8c���T�|~����?���q\Td�Z�N���}��JB"�(=���B��7��b�xh�/��Fc�Z��p"��������x�{o�ao�4#�i����K0�!{8���Q�/}�|���K׺N��Po(���P*�$+nyhˏ�;�����_�$�3Db�*s���ۂ0�&z�Fu��>�YN���0G�ٛiÆ;�2��fŒ�:ه�[��T
|:���^+�hU�NKp8C^
�����R�����ޑ��Y<��|���+]�����̎�<o���@�C�Y�CL߈��q�dŤwV`��٩���B�8FZ�#�q�p� �*�H��K�c�Rvq�G|�jU�E�>�<����|̳~}�xߤ'�z��}�.@�_���%d؏"���4��x�օ0�%]��m���/�n6�aFp95��߼�!|hݼA��ЎQPY�G9��o�Z�N�0v,��"(�c��4�.{�7��\���i�mڴ�u��B���pz �o[�NN ��Ok*7��_4���w[�hgJE$[�ULlJ��WNQ,h��xϾ6G��IlN�t�65T�n�ĝS��"��t�L�"l!O����ܨ����p `B\#�ݑm�f�	+@��{Y����)�&�D�Fk'��]�)'�Y~|ǐ�,��y�E��j}�_�t�m��Sh�'f���=UBmi�K9ȸ�NG�Z�?����f"��l�z��@]�6�M81���T&���y����}B�lW���)���Mr4,�c�0'�6���;�Z'�b���m���30�Gy}
�v0+`�B�̈́��6�6�|�S\=N�έ�vʔ�/g�p]E�Sp�O��f������E�����7Z���>v�ah��{4��1h�t���:',�9������S>���G��jc��Ө����NØp{aC��Xa���7s�3Ԥz
S��Y�H��)�3^Г�J&�8��34�/�
)���\ʚIs^or��.��h�b�c>ܸ�)�����>
v�4��v����{#'?c�,�<���R�����3�z�q����@F��p]�"��>y���!N��K��j"�/\?��I��%<^Fd��(S�����&�n�[B���綊y���S0��Pk�X]��s��r���*Ň��6A�h��9�H�;���?>'d���?�*�2�č�d��g?ے�w�Js�-Ȣ�;���k�Fv��h˹��.�限��:t��Nqmգ��hv3�>ŋ#+��G޻��`
����Ut<�ω�v���5/#I��T�9�CbHhL����؍�h�����]BU�Dl��	�����O�>Mcis��f1��W��ʈ����;ˤ[�k!�#�4}�uJ9���V}Sn����B��H��8blk�RF�i���^����C���&����8<�՗{

�6s,��ݗJ3����2g�6��	�DfDgKM*zA9Ei	z5:�U�{{�uwA�C�{��h������9,��Av���%�ZsY���K�h����� &K>^��½������ҹ��i�I�y�߳���	��^x�)9/��p0w(���T'��٫�pۃn��B�g.ŭ����f��y��2����`���w`*���ז�#|��#��nѬ	����w�e������ >��Ey����s�h�<U�/��32��=���s� l5���S�)���ھ�l�V0F�f]��m��FL:GB��m{]r9!���/ᜒ�F�aX���vNLK�\�$ �vzj���_��5�[���l#����*��[F"&=�"�5u	��l�d�fUg�@.�%�`���M�w񠴢��~7�l�-��8<���d��_DE|&���h��[[u$�]6�a���g�cl�����$�H�<l�q�O���U�nQ��$��qG;���<�KhB)H��=���m��9O��3��������������W�4:�t�3�e8�UU�p�o��Qv�^���� ��Kp��GPc�1�1MF`�x3������7(3�?�ז8����8�Г@��'Q�����a�
p =טs�" ��C3�},;I�>���c�vFx�Ɩ&�(�t�����E�m5�!e�1'�n�Ϙ�;�ŧ<��l.4��C���q������0~
_�оؙݙ��{�w��u���*��s�C?�G%YX����-/�\°�D�:��河���Ff����3����ӆ+��>�b��/�� ST�)�#	�)��7���t�FzMdI��\j�	��G۲O"��xE����WS����|���c�R���+��c��ܿ���r�1�N�����(� |�2kcL_~G�(4�'-<��Q��C�=�gi���=���Fo�ZH�a�Ѣnx���G%��P���$�ˉ���m̜���4x�� �Wp���b�Z8�o�+B�F%�����;d�>+"��Xg	�{��u{-��g_� 	^y��ɢ��I��Z�4�Q3D�r�T(��oݦ�2ٹ'i1�熁�y";���3��l�m}W����e�|��a�ͨ��xH�ߍ`^A@\:w�1�O�u� Xۯj�ۃ��
�U 9�|�0�����t�����񍩇���ݵ����j
��t�r` I�5���D`�%�pLǔ��V�Wïv)ծ2��_+fz�$�{�v�}2�1X#�bv+�#���X��=�{�N��9t�qv������p�o �܀�i�:V^����z����s�Kʼ�H�*Hr���^����`�����D ��=�g]����BZw y�ž��r/�ٰ��qQ���!?�T�hz�W�7����� x��p�g�s�M��O*+�7��%�j��ѹ$�7d�gP�!�U���<�V���.�7*[�IE�z����l{T�3���7e�㡟K�nF�Ǚ}�6Ś��Q%�B��{$���6 ����Ջ�z$
F%��TW�X�4i�h���9�v�ɨ~���4�f��*�~4F�JR�!X��
�8
�+�
k�̶�`��lBmJL^���j:����*hX�D�4׉ꎵ{Tf�$�Ec������m�?BpSc��c8�t�E��i���њo�E��E���h;\.FQټ�C60Wp��n�Z���)��y)P3�N��&��to"(��T����q�T27.��j�|���ڳ'Pg�J!�~8	k����o�ɧ��$ڿ��5�-���+�E��>~ԵǊ6(xRg]����+n�K����(�E(2��eJ5Q4��-Ց��9ĺ|��/���yi]��}�G�O�����R�|��G��s�a;I�n���F���D ��o�n�窅tč��G �bjH�tAЈ�����{�h���*�-��֯�n��p0
o�Fd``FS	�A�7����$�����)I�Ä��y���J�_?T�*���⭶���g���ށ6��tuCv�F�Ϡu����"�cݢr�$5gylz�a��]��d9O4�~�2?]o�(
������Cz��Ş͏}��=5|�c�z������M�ɩ�t�l2s%GHk��&�"5@{�vؔ�>�Ȱ�cp�q�t�r���������6��YL��x�l��Gha���F �ou�ڲ!Y��2K:6��$d^⮭<����;67��E���r�|ߒ0���{�A)�~޸G�)�b��ӟlZ�����S��`ݎ���=�R��ۿ{��@=�^�Md=`������S֓�Jx��׼ �{��y�'��'{@O��T�O�RoC�ڍ��6����ձ�M�L�����>�:Bz��N�#�o�������e���2�z�����[*%��^��+���n#i~�M(�.�h��&൭��)�b��UG3�&u����es�|`o�p��ы�[j���k�$7UƗ�x��CL��O���Bzls��Q�!�*�Ν�/�|�T.���j���Z�Њ������!�{	�`*���1X.z��k�o[AӚ���p%t�_��o�,�#n�&�!_�27`�	`����}�uR7�ˏ C%r=�������'S߶�|E�u�I�n1�!�<n
���+��sD�����[���4� ���$��PiuJ���	�����\&Xh	๽9R���Xu��(��q��������f��֎2�7���E�A�k|�w���俉Ϗ�Q'��
���)mF����ŤR$�7�I�jm��Y��t�@�}DV�:7��Y�Nv��܂a�h�~
q�Z�?��P�ޕ$ɯ}��ݺi�c5�~�x�J�vd6xB|��Y��U� O�05C��PZ8�L�-ц��Wa�3�m���i�������Pҏ���Ό�j�f��v����T-g.c'�Z���hZ��(w��G�4��~�L�UHE��( v�������-�ooi��lK�U�>o�����&l�����yb��:�Z<9N��=�~�k��ި�h���� � )I�7塐TK�qƕ�i������*m[%[c�c��gϞN���K��a�A��sCs45�sQ����B����{>���5ƛ{�[����7i�����/rP6���
7�
�NW�Z�h��]q�XfJ'�M�W	Ä���[Mǒ,��EK#�Lz@���=4W�Œ�
�"t�i�������<������0H���f�l�]���~���Ev!�[i�f�=��N��=zP�-��,UzE��߱�vBp�B�f�y��+X��m�Xl�~�f� �Ǔ<Bکj��D�&���]��	e�ݔOc�I��s���U�${��f�M����o���q�R��VOE��"Q��1���L�1��tw���Ĺo��e�C�����#y�݉	��N����ɇ	��������q|+L4���5��G	��l{��_���RWRY�5g�W3�s�����'`-P�?޷N�R?�K�Xp���yA�һC����,D+�{*�*����t�Krf���f͞m��-B}6� �#�C_r�3��'C�������O�cY���X�e	xC{5�\�UP��K�yu5t/ż�ݕhad���?]f���f�`�Wքʞr��}}.�|��s�(HcԒ�q�R�W숛/Xazt���\IO�a�a3-�@G�8���gQ6^� ���Y��|i�ѕ���໫��5��w���3���8,�K,��a�s�$�Q�r�DB�>@F0Y+P޶���m�?$�ɢ���V�>m[$��4W�`����)��GLV�O����*�%��e�88J�<ݹ!�
�e�g.D�L�k5��Yo ��7��t�R}�����tkC@/`{�z<Gc}����/NW�S�]�R)��M��+�faVN��7��|�0�S��}ޒl2G�6$��ou@S#7/rir6�Fn�'�^���عR��ho�+���K,~Pa����t�P5��tfɃ��u��MyR�P �:'~)96������8vsR4���\A����SУ��ߴiϻo
�����iB����f>��O�^-8:Ϩ=�'��9j2W&�LoE~�f|ɘ��E�'��Xs�������=�����_?<y/G`o�\0�+��ǯ��1��fq�;�>e�غޏ �'R��J4�x?t��r��Mz�d&:���`l��6`��[H�님�����<�~����Ҕ�x�:���3dB��S7Ά���FQ�|C��t��P(rˤ���O
rZ���;td����o�O������}��t��L�� �%��p+(�U����0A)�+�4Ѹ�)w�^�i�-��%�%z���2��g�S��B��PS�ER�*�|6W�����GW'u��]�_�Y�� z�]h���$
�߯\�Dg�S4?w�����ݎgZRDy>f� ����Q��)���Y,��,v��Tf�`V[�C��c�6��+*J�U��e�x�o �\�5�,���*p�x����I����K2G�ٳ��z�R�v�um�����1$t�'|o�#Ve��\J�ؠVC�3�k
���U��U���=6�B��3�I�N�	˽��B��&X��d��iA�6O��/.Af�/�,ib弭 x��é�xQ��)3�:sN=��y2��H�j�{�M%#֕J���,�a6Z�!��0(����l)�����aπ���:4����c�h��#��H\�$J_�؆�m��'����&o&6)3��E�ظ��zƯQ���5pF�ZuiN�D�3��^+��v]�6bF�k/�9�Ӟ�ʷn�\�}{�7N[��[Y�ANC�N��zS=��ΰ�X���vXT�8�`ZA:�n�u�l��4�X��M���جE����E�NNw}�K,�s���u�*���#�`%3¢O�M�HQ��\~�k1�
k�u��7�H����0�TI\�+e|�7�IQ�|�M��B員��C�"���I��?�ÁE�p3^����[)�'�G9�}kb�qb�FT�^Bq�H^��a�Ǘ�	tD���V�58l%+�?�On����r����X4zM��?C�D��"���꒙#S���O�C&�@Q�=B ����:|���ij��YN8\�qH��(�p<<YI"�S A��N~��"!I�B}�@u%P�>X���n��l�ob�hkF����v\��^TQ�:i<�S�e>U�R� uoG�d^���ͱ����ٰ�܊�"h���#c���@F���1�(���ʨ.��0��D�O���� ���'�tJk�c����Y��x.?"j�cRK��i�����5�|O�q���{��r�dt�`_�K�L�kC�MQˠg(�d���a�vE}<5��`�ô��ZMO�SϏ-E�=�W����F@|�Q�6�ۼ���!㷥k�@�W�z��t~�����z-ؾ]g��s.�R�D�A1�%5���J�>S� '����p��j+<?�u��og�&!�9e2��}1k�r=�����(ް�lB8[�Cb�5^`z6�Y��JA�LB�Waw�J�ͼ�/=�O[�� e�%v�r�]��5��Wi���`���
o�%��E��;(,��ACJ��(�+e�y��o|�)�q9a7+�em�@ �A݆WN�w
����9i�Ǖ��]x	鶲F�����S]=&�(�Bp�#�ۈ�/���-v�@��q�*�7y�	��h�Jf����x�}r�~F𒰿��?�A`P�IC����]�g�W�5Y H���T���q��H��B
�j���v����a�l�30�~���m?s^�u�nI�h�h��Z��MuЂ�����	7�LV��x�'P���G��A�Of�u`�bʐUI ��X�4^t^�v�N'Hh��n�*=�N�h��_*�:08��R"�F���bO!D��F�/��B���\��ۊ� ^@���s8��K����~D��\�G�&|Z������U�}+`7;��Zg,��x�@��p�Z2�B���
./r�������(ft��"���F�ŧ{4��Ш�%��tu�eؕW*/��{%��9��s5+�x�$->Eu�m�>0��z�3�3g�#�wO�?p0:r��h� a'���,��?� V���S���84��l�NVv�V��@��"��`+@��)-˃��E:����1���(--�- �X�����;<��'�M/v_�BC������W���QO�3���U���Jg�>O���B�=H�2�-��>�-.g��[#W�X!����R��7 ����`Ƞ�T�d}o���� �S��:5?�0��Im1)W#hn����z���<�TD�]�m�\\XU:�Zu���@���0o��Y������j0k�����j��w���exSO�fϙ�~8�p�yk91u���e�R�x҅���_�'p��^XZCY�y��i��
_����ޮ��^�r*�Lྌ�� �7�q2U��f�S�#��<o������Q�:ri(�(�E����4t*(�����[����8N8O��� �V�Bȷ��,�v�ʏMF-EHP]ʐҽeg��)�YM�t�r�ߊ ��=o������i�@��Af�$�˼������P/{A������0����(V���j�6�ckLck9�À��3�����9W�.V0�u�Z�X���~,0�$"r�+���'�9� �����Ul7���twJ|�^4�����������]�]�ٳ��K���U�O�+�ß�k�|�-v��9�99��	�E���)�[�}���4z�U�����m����K�|hzpPc䴤9���Tq�:xX��єm!�!3�'�m4���A�q(�*�����q��_a���vbo�Q	�����k�{C�痑�t��	�'D�ف���h	���vt��X�AN M(�t�S�z�F��f�Q���6��S%�N����t��GY��U�aM�ߝ�H�δ`'c✏�5�$�Da�����O���(f�>-������˖@��1j���MڣU+kӅ�Q����z��Fݱ�(��D���]��͘�(g�"..E�ǳ��rLw?��	����z8c##i�b�����O� TRڂ�7���%N���7�ذ��Uz��#��~G�w���i�V90��SU*q�]��-��!j����#��Q�&?ǭ��+w9�Hd�=��8o(u!
����Z�G����6	])}i'�C˝�&�/�"B��8F�0��@%zd��������J�`$�e?Z$��-\��)peS�Y���&�"X���#��]�"`WrĀ��n�?�߳��23�-C1%�O:���!X�2�N��P��ߢ�;�|w��1�����r�r��G��{n�/{�ؤA����e��S�)Ψ����h@}1(����q��;�LF��E����L1�J�Ɵ���z_ cU఍G͡/�S����A�R�-�+�ӌ\J۰g{BG�N70�jc�7�y@�m����Zpx��mJ�4g�����'8�cN�����%�,��I�C��e�CA�U��-=�UP������ �1��}&� G�0��*�@�ȣ�1	NRWw����<"��Z�ɇ� 2�g�#��\%"�l�98ZX�mjz����ذa:�..Ʊw��Q�:!���4.���f���U[��W9���g�"��.z����j*�0՜2*��pI{s��E@�PI���X�#�������r܎C0�1����?3߸�,�=�`(��7��]�&�Y��݆�\�vz��~#ֆ!:�$�4��8g>~�G3ex��ON���
0�C|,�jʖ����1�{V��{S���E�@@,O��H�{� �\��&`�����P߼�q8��G�I�IEǬ��D#�e��%����Q�%�)�����W:�b,����_(}��
���e@��;?�΄�T��?j�I�������[L�%����~�����q5�h�~�Ӈ���M��*�*W��{���Lv#�n:d��	Wg��ِI���	yj��/��H�8���L�������U�P���A��V�6k���)ύv�ح����Q��F� ig�F��>!�a�!$�H>,}u5�*8@�d��5�8��6n�媅L"�	�zI�i6׋���AkB���/�Y1�����PS��'̥�4j����4�#�W/�ң�,:��X�`z1~���Q#��l��{0�	)�'q������q�қp�JK5�_F@�x]�m��٩��a-����u�V���( ?&#*�2�O�(x��*��0�f'���	�Td6?͖�W��W]ba�Bw2b���,�$U�����ۂ׮;����6Ӳ��-ں�f8i��b�b��������Pđ~�!\UxErǳ\��-��Dw�x�y,K<3Ĉ����]���	��R疫�R�
3Y+���H�zr�5q���{��#t@���z:8�[)�?)��.2�.dg1:����b�����>����L�X|�|��Zl-*%�*˩�ZSVj��gb���{܌e��"��o�H#��N�Er(L�&�{��s�?� �Qт_�*'�_JN5Q4�P`����+�����R���y0G��ϙ닑%���T��n�o�.�[�6@�d,�f7�.zڒP��+_��S�zA/#���	-sQ�=�.ƲH��'#�9��r�:> ��HskLv1�޷8}=�6Y��7Z'�[`!���c]��\C���vF�B���~w)�-�G�q2Q]�>F��Ob1�p���4װ3j��1Տ@MF
3wι��I��J��A��z<2��f�T9�����H��2�7���F�v�mKD�L�7+�K�H�2߿�uNi'�JfB1��\B���$�d_0�i�Lw�����W1z̽��xO9�6`C�4Z:;9]yF.��:���JԻ���\à@�b��ob\�C�ތW�[1��X���[b|�7����+Q��͢"�j��=-;�ߒv�m&qȇx��1���+�����j��K��9��̯�h��v��� v�Q�L�o��^�[/������e	������@f|��F�c|'�4V�ڽ����7�����Tl�&M��\#��Mq$j猈���GT��FF�ݬ I؍�V��@�P`���\�t`0�|� �����n(�|p e&���؛ƴ;�Ɲ�k�䴒!㲈-�r�It�G)+N�ƞHr���p����y9�i�h�� ����)����R��Q�I�>����
���bS�7��0 �)�oaǣ�y��w��C�̐P1T�ی���l�G�_��#,G{;g�j�5Zes�V]pL3D�o��4�S!���7�� �<���4�)`���t:z�6�Q%s��A��|�B�H�0�%��xJ#��I�0<���of�'��E�nK���\����:^�ߤ�s���:~��;����FU�La�-#ޏI;[}*�<��_�AD[
�M=|�a�WD�Fe�]�DR�+u�hy��M��]i�\��?�$M\���~���%�dG�7i?K�f����C��Y�`����-~^A������������f��,�����l�E�B��r&��j���#J�	�>0ݲc٤v/�ᱳA_��/�OQ��)��{���7$2���zB�=|�w�ܕ�l�*R��˲CY�R���}��"��$�4:���Ktk�IlCX6���Y��)O� T$R�T�#�t�Q�\+��M�i��!��q������G��$ t�N���<x��|�J}.]������ى\-���M/�3� �]6�i
N@kD�B�����(�	|]M`Ke)n��E�� �8���P�LK�_����<�6D� �[P�l�x��}�,�E�)S"΀i�hH9�Z��٥Ž�R	:DkRp�SB��;�E\2�v�"��u@.HvA趁���>�흹pw��;�;�`��ƽiz���v1Q�}=�pW�R��,.`�F̂�o�Zƺ��$�����T%>�����9Bj���L#�+���~���c5���Y�$���tϞb���s�Xd)�QYr���Wo�lW��['�_XRE���F@}�yت��B4dj�_�t�5���.PV���h�� ��z����I�]���(����Hw{�H@���`��I) J#)�{S��귚>�P�e�Kq���R�f1NiTJM�Tɚ�I�M(�as�Z�'�#�l���4GOi]F6Jqߎ�Ӑ�Lמ:��<^����,�{.��SV ��ֻ���_��2�`�Ҳ3�
Ԙ���݈�# !�xT����a�y���@Hg�P��ɩ�T�z��_n\嚥��U��g�L�pC�����F�@�\� ��9��c6wC�����D��&J̱��� �B0ʗ_��5םPP�8�C��y6�h*��O��aVVc��nZ &�ִ����0T-K^ä ?�E�;2�	�;|[��w9��b2$��
�Wm0�@���y�{���J�@*�"�Y|(֧�Ҁ�/���s�������L!��(#����=@=��p32% ��u�bݎ6ܪ₦LY{�y~9������B���<���!����"��g�3W�k�[�2�2� ���[�ܪ2:�<���ﲩ���A�w7��({���pq"WK�FE�`�;��l�vZf���D����q��"��P��<*{(=_UܣœU�:>R@;�	W���L<6� T��%nk�EYa��o�Z���08�R���l/F
U���U2�6@�xA"$��6
��X3�Lj͹G��x��ԋ4��6����~w%>����Zu;%�&�#p�&5t�	�����m��V�%�r�xX�f�_(M>�V!'�O�x������?K~-�+��X^��8 uci�~:;��I(�η���N�8r�y������N��;/"..Vtcȃ�dН,�tgL6�d�Z�y�+������ ���%������ASX0nm�I:}e���(���	�4�X��K�E%�7�A>!�m����p���(|�I0��Q$��2K�7��V5n��tèV��:'^s7p�����A�&T ������~�:��0�+��AN	o%Wű��Bh�^r�]���v����j=�K�	���}�F�\0D6�jQ4�@��W\�}�*�����%��S�$
g��������$�)�L��C�f�|S�֛�r;C�S�aLC��pK��N8���_��+���3n���E"�����Z��ǍEo�����w]6H�F�"O��������A@Bo&��)�u�إ'����L�`\���'`&J_�>LjK�H[�w)��r�.���x�/[\X�ā�X��M}�i�h��!$h�6h�3���y�$̘�u<���6~g�W/a����>�'\���7��C+ s��~n�Ϧ���~3����]�g��S��9 ���� �< F�W��wl�d�Ps9��Ap8Χ�����6����mP:��ccE�#�`���3x���p�DⱗЦ��v�-��s6��<0;N�����U]кMd�d�i���אC�>���}'"ʕ\�KC ��c�1��JԌ	�fn& ^���KϹ�^:[��Kp���{���ѨV���;���@<
!� �>�����A}�&���ǅt�a�F]�a`�Ҟ�-��~6g_�S3s�E]+K$,~�f���oG�2sS�M���?]wP�] ���UW�T� Rk?�h�����;
�e�����͒�G��0�H����c������G(6K�L�憮Q�{�cZ����d��_�J���Kqԕ�������n��7�껭�x����M!ߠp��1��w��֜���/���L�J��G���"����b�2�z�9CcBϟo��Z����;$���Ԏ,m��2M�$|��s0O$�
G������̝x�w
����:���8��VXG6+�h��5NR-�����-KY�1|y��e.�s�Za��F��L^��'����3�S��ȕ��7@h��d��/���OBO)H*[F.ӓ��Y(<�5:�������0e"_��Q���[T[����	_�.l+��_Sǂ�"Y�[k��m����g�j%,���| �(�$�&������f�^�	�2������ɰ_F�{Ilm�Q��+���h��z�?�;�k�Q�2Z"Q˳��.Tࠕm����o�T~{�6�w�������zʜh%*d)i�:�QLHA/�S	O&E(u�k�:�#2���=	�p�t@�f�iyY�T�Д�D�(h��a����#���/k'����T��bD�v`F:4���U>(���n�6���莣z\x ��8�@A��]9��Q�q5�m�SY�q02	|��)w���k韵��ʅ��'N_rCX6EO)8����L�.�oW�!����}Q�F�mU�X%��>�<�g���C�Z��a�7<��s�x�ڰ�e>IGd�*��$�R��/��d}�|��"�x��}��7!����xƒ'ё�7-�'�Q��pj�7���o���fW��/Kf�����qY�j-�H�C��;º<�'�7��O�y6�����������N�?E�u�	�>�r4�Sλ�����A�����x'���Q����H-��ﰽ�r.4����:t���.ܔx�ʌ;�[�̏ë������j�B��#y��$��\�A=�_cz����M�����,R�1������D�ڰ�����BQT�\�h/���1�Nw����T�G@	�@�X�*�T�ӠQ��wk<}�4ؔ�/]��t��icz�50�,�m<`S��6��[�Ѝ�t@���5J��n
���\G���j��`C7�7�A�X��[�beE3�(��j��c��Wkه_;��gϿR��J #��[�Uַ��&{�;�Lz�^�Ut�B���лhX���0��*
a�1Tr)��1�zr*�vCD���O���Թ�%�l��	������66;�{�g��@�#����ޠSE�`��v�7��b 1�b��ݓd;H�Ec+o��<�Q�$�V���'�,�I_Md����u�U�<&�
u���虌�m�'�w(Ս38�2U�~<z\�)�
���W��9,��&��c�D��=j�+���v��_�B5i����	���tt��@�%y��ɸ&��?�!�3C�ԯz{�=u.#����}���f$r_?1��{����q@qK�ě��Y�9t>���g"�#�X�a��q[֫�Á��q� 9o��9�Ǳ�T��q�NvE�ܓBSt�+��i�n<G�U���w�<UN������l��Fb���������(��:��#w%���t��b�ǌ�s'�<4��>e�v��L��j#���֧{��ij0�'� ���~���4�8��M�"i�G�9��.XV9����/>�/m�j>N�9����M�`ޯ�T��-���g*_2�bgYF�r��Y^����g��,�!�і�]F�X~	�,�鹯�� �$G�d��s��ʃ��9�ΗI�;��ž��>;^ᣇ�@�ʿ
6���tZGY|pHP�Ekk��.����P�j��IC�b�I��:l��N�3w�j��ԡ��M}>j1��^����>'��a��H�Lg����͈�#�L>�)x*�g�Q����{�b�-R��O%M�����A*��%�^�c�M3�:(�a�|��f����p>&����|蟽�E1�.��`6��O������*�3y�3��E\;sw�4������4w.�qȝ&P�Ґ}�ԓen�R�E�=��'��� �Hroځ��7�Ёێ]������q����X�j���:9,����s&�O�pƠ��k?�K!5{�O.��&��,��N�P�+��I���`m8	;	�y�ͫ?+��1i�=t��e�o}Qk�]r~t�	3�Ri&�~��<ځ�QH�5��W��wangL�#nF��Nll;bq�j!Vm/�Ω�e<VR.�N��җ��9u1���������jC�-�!J�ۼ�&^E�������O^���� ���Vƍ#즨b�����?b��O�/�	O�f�ͽ�p��(���X�$��H�����Կ��VN�k��X�\@|�fYwV������܆���� ��bB5	��h#���a�эo}���ݑ��I%�hHǅ$��oo��z��G��ʹZ�Av�٧��b.���ʅ\��fC;�i3Ө�o�œ�sZ"g���s ����m{;.*�m�D��5y'R��Q^0.eĿ-D�+-�%4:{�-�R�d�_l�"%����_�@�	Xɪ��HTF0�����˱���]IE�'CԀ�+Mv���@��^&73�f���xp���`vE�*�e��v4�mc�ý@Q�A��!���x�6u�3�/�O>Z�RaH�Ӝ��{�_#}k�6�/w/"��fT��B��l�N�W�l~�?̊Vf�����*�����6�0���k��p�;�wS��EWX֠�x��	�����c"���
�Y�^ߒ����Pp�M�ɲk��B��K��1S�(����_>�O�<G�$�_o� #�d����3��T^֜jx�^\�x�����{)��/�=X���p�p[��k��dK�wN�i���"O`����������2 �<*�x#�E'k�  �~n��6�C�-����Z�{Y�k��y���
w��V�wz��=�cSL�x�Ր����݂�ly'���Q�s7i1�����/U�	��2�&Ѵ�, 1*�~:F}Q����c�&�|����J�U��N�a'�9�ݨ�3{y��갳���sr�(�Ye�b���Mh�ԗD0�;F�QR�	7��]��t߮���#W��o��i��Wˢ6Szɇ��H�t�j����KN�z�4�gXv��������w������zE�:�>熯�k ;�5��4���=��[��~��E��(�E�.���w\Q�4'@��p��&B��0]>I�`�����Q#��6ӆ��� �B�d;�N�\P��=��BI��X4}.*����H&��=��(����rB���)��˽�˝Y�B���m��#���l !�c�O����N۪#]����J!�����G�E��rߎ������n��Qh+q��QT!��L�u�P�ld��&����@3�|*bP�Wk�Lx'B�̆@�=� #) � ���W	�j�u���yÈ�C�j��0�Ú�;0��2��5�7�~k9��K_+���	��	�?�F�.���r�N���&�&<N�Y�k��<x�Vr�+�-�7?�	@��P�:ՠ�]^�6_ɘ�C�Y���`}y��/a�ؗ'A��]����4n��qz���f�����իřM��4�o�1qhDfѲS�-���W�������;?aI��0�8gқJ@�4V�P��5h�o�T�#����?dB\Ƥ����-�?0<~��C5�9'-���F�7�q�wYY�3w��ʬ��*t���O�8X�i�/����&��J)+7�����M�x���'���؏��,%��W7��v�+|Q-�l�脳]k3����!�7w�����A$�D�,���X�NޤUZ��y
>'�[�Ni>�j-�r�ꖩ47Ci2I���̼��Ε^@��_��d��l��pDY����8!�^�p U��}m��|�h�XQ\ڛjWǈ~X� ������t��j��(����c��@���.�O�_"�;&�ɗV.?A�OE�Cn����8]%�
������xI[T��1Yt_�d�.��������È:� �ηW��G���!ʹ 抒�����$��-ER͏�m$7",�rf���3�:jB
f�լ�ڟ�^
:K�#��6$_��q8�Jtr$�2b����I��T�E��ߌv?�X�c��1AD2���F�?~`*�s�N
�����e���Ϝ��� +&75����W$������Lh T�%�p��"�o���<�'o����cN�vC@5?e����Nv�V�
)�Yg&Ce������KҖ~�кF�Ԇ�����v����0�o)'����O*^pu�<v!�s*r7�F���5Y2?�g��^�c� �fެ�a mO������V�
:v��މ�:�3�W�W�Wf�G���Y�4�&(Ώ*2�ý�3@��g���!����k�ƥ
3�՞N����>�q�Vwm�Ư9 #���W���#X*�k���� dlLlGu����kȐ�<v-������0\ѧʐ��ŉ�lb�´K���#'�L���NqĿQ���J�_�����|0�e�G����M��#��9O���>�����2vvd����,�/C� �u��]m�RE�ˋ��W&�azZ����?w�`j�e{L	W�j��%Q�F*]��c��l>�k�5W;�朋�%L-����@P:�R�%�LBD:E��/@L��a;��Iq{����I+gj4޽���m.\��.c�[�����j�@G{
8vS]�1��X�4[�}�[�E-HV9�+U�ȿ�@����"Ar�F2�Ǖv�T������l� �/��a@��cɫ�5��� ˢxc�ܿ���j.���v��UH�ڜF�D�:)�P#U�ɉ�X���zc��R6��Z�=.���!��K{֝v�P�,�i�{�@�xz���:P�Y�ڟ�S��`%m�A���{!i��D��V�J�d����Gk�y!��a�0R`�mŞ#�=���7Med3���9cN��p2.^���;�9M����C,�+�G�HTV.��_��;�p���=F����lf�җ��Y@�&f=��)�0����8{j/�T���f[5��L����d�էg�ƄJ���8i���w��K��X'���ƤP���h]�~h�{��S� �����R����E ��ȺUPO9��R�X~�0� ���a���Y"݇����i�刣júq	;��(�p��&4��8X�ck/�7L��WHJi��AYb

�	�C�Jn���mB�:���H@�3��yk�j�ї�$7)BY{4�AI�ї�7��V�}wS�%�_z'(4��Db��ȟ��^T�W���m:aq�t4X/�|�T���s�SB�_	�J	�	�^KLfNy�c��P�x+�������#B�EdXh���t�r8���=O���Gg����Z�Ґ%;�R��¯�b����>������Y����_`�@����&��}�;�tE�eoد���^�]��d�mrI交�S.ȷfɅ/^~�I���/�P�+�oE�^���N��\�MoA�H���Ul��H!4�3�>AD�˛Du�@������ܝ]	w��#Q�6xF(]6�)�s���~c_W�U	��^����D�zj��>����f�c~n_�kI�Ej����j#�/�����| �j��j�)N{<���D+��{�?��tE�K��$܌|�{/�t����1�^��^D�����P�Ղ��sp$��%�Z8(�O)2>�.[�1��*�wS���Zx�2��q��ҧA���3��H�cE��i��v��a�
�D3g©$�AJ�x��_nUQ���Ч��cg��oOY�<���lwm:�)C' M}�m���;3�od�!BZ	 �y�;�����wkp�F�b9�����U���x��� Խ�?��9��i%�o�Vf2t�8^1 ��Cu�e��.���F��Q�
�#f���.Í���~�ȸ��x��m��^~�o%��c�n�7� F���B$�C��{�$�>Ɠz�t^���G�d�A���Ǝ�����$͸�'0���a7�vi8��F�:�-jȉ��O lh��21u�c"��Cfip6L�����r��޽��HA+���?�q6죑���H}��n+��x.���-�2J۩|��m��h?�D���%vKR�Ӵc�dI�v�80��fQm|��RS2�?������C�ڻ�c;�yY@V�I����8Щ�g�m��EƋ��ൂɏ������^N��|Y�'����ُ{�����(}�Q���1nK��V2˔J�Î �2#ւ��X�o����T���t�0H�zm������j-�\(��=6L��F"�E��p��}�s �w�m+����Ѳ�W��*E�u�mo
�ϸ��K.=�OC	'�X�����U��Y�uGRb�����s��ɐ�U��y���/����8�O�"�
�Ua<�"�lt,����$g��ї���#,6?���`�R3b��rk�7Y{�S� t$�|���|�	���1��A����Ʉvte� 	A�k��8��������~��\c��V�Rj���FLG�a����ïdަaT��d������!4vO���_E��Dh��WQ?l� *FgYw�Q���O�ρh�="�c�΢�gM�Ć�<��_I2Ͱ�I[j~�,4Қ�A1ڵ#���S���N�76��3_m�Y�U\{;��Ս_�?] ��ML�3e�rVCY��Fz�yӷ�['/�����	���ID(��e���D3�ۈ�� $�R��`��Wey�\�A6^�+����������0bo� fbV���6����R_�"��2Ef�E.n���H�˃o����1�(+���� O�6�>��]Pl��)NX̩��>��Ŵg�@�B�Ȅ]I�H��p����!��S�l�\S5�b;��W��#�X��ֶu���r�����eG��K���d��x��+�O`���\<H�����8�x���px�fj�z��:>3 $l����f}�Z�=�RC��Pw�<���*���iPRI��Z��١�b�E�5�~�V{9��,�C��F���xb�d�oī[Z����+��O�p�_#�cg$A$�5Y/����m�W�{*f�#i�b磼QPJVLMk|iV�V�2R��e.%
��_.�}I�C� ����V�����>�k�+^9�(q��Q<�m吿[�9R'�=eX��?$��Ȱ���p����^z�SO-���kϵhhC�}4�wA����X�o��S�J�X0U���ٳ��<fr�řb�,u�E�:�q�.�D����9��0Mu����c��#[b^�U��\�9aC5Q|�%R~震�'��s&>�'o�嬕\�C�q����^�P�	��mcl�����q�8d�hqv�Z�����A$�InײԜ��|��6�M���e� ����,/�+�&��qlB	�0�.��P�����e��DG�*��m�v���[�!�I�50v*.�-r>�gk���[������6�Tس{
�KQDH�d�3D�ۥ#�ޘp�
Pw�|��1dز�h�8<�-�U�7n��!�V�+NT �c:հ%9���+�'�F�DD�����3���ȶ��s�7�Zș"�Ԟ��F댲	û�+�P�Te�GU�6��WS�7�.����tdI��e9ٳ"��D���W[i��v��15pC��ԣ�t-�~��q��x؞ؠ�l��>(*�8�<��R��=5��wO��ϐo:Y�q��9���U���w��WK7��� A5���7,y��t|���4����n%��ɪq ��;i�9�K����#��K��z�9C#��h�����ͩD��+���ǣ���A���6��5o����P0��m�hN�dq,�*��@fl�$���Z�����7��>���I0�[�QSr�	-( %�f���\�uK�M���v��ԛ#|�"-�&c4��䉴�Ysb�5��4L�3~�u�_���vsY%���	�<�\��i���\̆�5�Ț�T�d��=���&_MG{j��C��EJ��|��*T9�(zΏ��C���g�,���&�VW�$K&P�h<���ؖOr&j�p�ӱ�w^�&{MtY��ݙ��ؐ�f��^��8�*��E
�p}TU����݀fa�S�z�UuPĢ�Hύ��ĵU26�Nx/�4NF�/"zS�eè3?/�~��8�1v*DI&�ԗ3󔽎�Z���ڇ��]}��E�!5EZ�7�.0��ҦF�_�E��EdRN�b0��1T���Ƚ �Y�~-��
�Mt��U��#TEcq�P�+}�ueM���(��1V13Q!�~�)�6`m(_L����ޢ����h�"@9OHuw��*��{_P���V4�g��q�n���H}`z�+��h8�iZ�u߸�	���?`o(�l�GN��?�e��*|�������J�����YT9�b ��A�~�U4�+f�U"T���wgX���<�o­ǕwKC#*�1Кt��cqv��jp�Ppë�;Y*Kͩ��f�����A�0K�D7=�Vz��:��2k���t�J�s��A�1p�����֐p�[	�l����\���A4�H����j�xt�A��c��"�4bn����#�Y���4��ֆ�p��4��I���o{�
���D�]�r��I�� `X�1ڤQY1~��ҝ
������c4a�a'"Yܤ#��"�;��ؗ�a�?�k��+9?����lʨKF4��@3���t_8���PL�6�I��B�6���@�K%�s �Kk�X�������=y�  	�} �3�Bx����޽i��YR�J1�|:编^0�li�h���'X�m�T0�����LA�b�C}ʌ��a�ɑ���9�2�>�wu��L2U�J��H w17����Cj�J�:���~"N�F���[��j�;!�O�B�qײR�r`:(���Nv��I]�]��H��!
X�@9\�k��6���e\ȁ�҆�0�00���qq(M��ї�Ơ���F������ۋ�eR��Dp ��̹�9kI�`�5��}�;Q%�6�HMW=q���P�7o/��W�>fKP�(��[��D��ǫ��t�t� �Q��r���+�	nӠ�M�E�	�}VP��Q6�4Ѡ��8J�������a�f�0r��j���$��0�d����Sm/ T ���u�!����n�^(� �٨��	a]
���˔*-q�JqЈ��R3���|�d�G����H���L�N��+��&� i�Xَ���ׁ	�Hݷs��e��"T��\<ys�kZ	��R�e8��J�	"����g��d��{*FcP��%a��"E)�o���#�t0��)� P��6p���hp�Z)~�	Ո�����Úي]����+�q�g�H�	f���燣�7�����ٓMO��-����/Jx��kn��>�7I^���3:�!"�1��֟��V�y
�j�L�����;�.%64�r^bQ���?�))�4��۞�n�V������R���%Acu�P��;��8���t��J1��������k=�1��/�$����ݯ�
U����W�1k�-�m�ŅT7~�.�л#���!4F$���K�Q��@�ê�����c	�0Kw�$M�]A�x�ga.�t76DT�.*�M�OS[\��!����W�'��ϧ����1"l����4�$e�zX�tպY.s�A'��-�,�,�WG;GZ�K���+��}e�;W��w/h������t8����U�7�{����CS=t�,��p|%�N1�#<����=&�9&�J~@��ee�la��(Q��O讠�K�^t�r����C��霢 �����;=%��{���b	n����f��L�a,le�G�і�*?8���{�O�yG�/�u	��/3L��zX��5�9�7t��d���M�������W��V׍���~>cp���Q��޿��y�Ǥ�F��D��)���p0t�LGh����_)���T׼:"�|�����>ʛQ�B����Y�V�~G�w���A7h�`ާ�:�lu��V�#d}*���a���[��+[��\dۻ�d9������p"��Y��IL0��E<|������=W��~pk��|j�F�`�
4;䙅���	6�is�����`/(
A��/���Shu�B����`�_�����2��P���Y�urI[E�r�*�7�#���_A�x[:�hӔhp�]2>�Z$w�2�Xp�+`�����V'j�Vܐ�퉾�L�l�W����D�|tnb8	P�VOB�8w짵y|�:}� �v^�v�L�
P~eiA�0�,us���n�.cz��K��B��ˀ�T(�̲��H���kM�3�����_+HD����}M9��=6fH~��բ=���|.�So��e��_�V	Q�Pi�/2�-]B��֪�#�Bk�710��K%g���w�u�-����e�	�/I�g��%�4�f�Nʿ��]N�=���������xEtb@5��ͭa�&cp��c�P� K�A��������7�F�Y�$�@#���|v:�<��<^g��s6�ya���N�����>��K2_���������eua�w2�\#�xV�h���:X�+Q�F��m\�01���<E��B��"�@�`���Kh˺��-"�< ~�[%������p(��Let�.�'Ѥ)�է�y�v�7��t�0_�ZJ���q�' ����}�|a����ý�����Gr�k�.M\�1�1_ں|ڎ�C��;����vsg��<<�k�	+=���������8��j�Q�hA�P�� /~X��
\�d<�$�=����V�7?�O��۰��U磩o�Y�iwW̲���ih��&xQ4��ꐍ�?p��G�g[�L�d�����(���q�x��-�4�x�u-|�.�aY�tu�(P��e�en32<�ή�0`Bl<�M��d�LU�0�yҒk�Qx���4-~1��D�g9��{�B�+nT9��s�[�8淚R|�G�N~��
W_��˽zإ�G�����,������+6�T�J��{�J���[���q+G��;\y��h���Sv��]��a�Ÿ1�a>]�q���i�T���Pέ{x�p91杺ʏꕮU�,�ńLjQ��� 5ghd��g����_)�s�(�e�^����+ �5Sai!����k�=�z-"߶�E�n2�c0[׌��&,P��Ϫb�F�gn��د���X2�$�=�$u�R�������y�!]�"���"����ˇ@�|!*�L_ŝh��- �
F��.W�>h!������J����Yz�|d]w�KI1s�����s�NY����E���}�{R�?6��ε�@�W#zn\^�Ű�0�;�u��NqQ$�+Y���d\��8��}�M���Q�ml� r�j�G4�8�u\��0u�z�5��L5�f1hk��_��"M��2�_���~y��j*o_Vi$`/�	��x�q/ڙ��?n ��R5�B�Ef,��`�2̗��ln_E~֟7^��m����8��m<��͐~�u7�B�q�3�G�@ya��V���La�>#4<����`c뤡
!���|kà������6��x��a �5��iLB����T��,�4I�����R�U�1�uرL(��i��p��5I���;�>r �
��+T�A����{|��D�!�F��։��7R$Ԑ$��j��)��|��U;���[>��)P�����Hb�Brv�{�V���V�(uE����r���O��r� :#��2'y��
�,��|�Z���أkӱ'��B �������{U���N�4}b�tE�Sh�§�iLK㾤�V��s	).���#������.���>q���#?\�;o��N;��8M���;���=������(ي���l����`�М��������DL��u���/ߚZ�A{ˎ\q#!�T��W��Z�w�]U�M���}ɪ���[6�&+��.]|o���)��rL.V.��p��#���szi�v�u���!���;��V���y������7x���Ղ�itɍ"�ԞV�ʗ���5�����Li�9Fv��Ԑ�������9�w�w�_UD��.��S|�+G˱�kkOІ�Mʹ2Π�b�9aAV�Wu`�M^.��<7buUy��d�s(Y�R�����h�"�ƍ��NЊD��#\Z��qb���ཞC��D��r̍}��ש@��kM�����>�B��E��N��6�����b�E�Ӝ>+w�*W��Κx�!���%o[H��}��ۀ��#Au�1JC�P"��p�����W���gC	�a��G�T�b~qt�wBSR�Kl�`5/}��c��v����H�L��Z��{:r��sr�}D��e_��%���N���]��*_;MJ����$x������7���{��n�(��r~��vя�l��P��g�ބ�_�mf�aJq��.��vk)�ä_�n�D�;��̋�$.��d%X�F�3KB%�h/)摘���9���$��T�`���D�M�#��z�k�3��m���̝򭘤 ^��ф(;����@��Z�E
4��!\K�1���e�]=Q9�)�,��f7�p�3n|扙�j��ی"i.�~��KF�L06��£�N�ʆT8h��W�I"�9#4��|�$]���c&o�n�u�8Y���a5W�,����@��Q�~h��'&�'���C1ϦM��
���]iA�X���9��M�"�0����F�Wt~�؆X��@�}G�Z8��?�+����ߙ9R�q�g+���.&�PM� v�� �9Z{j�B�7n�����s�	Gi9����0���q+_t [M�`�㐰�>�)�����t٩��x?7��>���4�- m jS)f�W�"ε���J��'RB�����-	�U��aɫX �0����Z�d���/�T ����5���=]PK�	���ʩ�Qh�n�ho�j`��e�C=Z��b�k����	Tɾ���5W7���(m~�WU��a���XG�!�­�i>\\�] <6�]�P��~�����^�r]�|3�5V5nM�>$]�!Q�epР O{l�<��Y**�=��C�(�&E�.?�'��k3p+���V���9���1��f�c������v}�8#vT�Z� �q����gd��WT�w롭�H�1�ų-�������wx�����a�$תi=P����~����,��-��]pU? u���i��ʈ�J*�c'�;��8���Kg�#��(M|'
�?�[&�b�4��������A��%�a��+�C���v�>.���ۤ�_S:�u�/�"[���ͤC=E�퓾־J�}��t8���D�Ϸ�D�/��Sʶ]A%��!�Nh�4�ӫr4?�Bn�~4m��n�V8���62Ul%�R���W	�#U�Ғd��4��9z�����t��'�8C�#���q�#h�S�M�8�\ח��1x@v�vg�ؐ�O��|��4��W/!4��%���)�>[HM��C��ez�l���l(�Z�C��l�D�xjrķ8��{!$&��o�n��m;��F�׽��6�%���B�����#n�q�����y��$�kT�����pћX)�/��ѣ�)�;S9�yTq4��V�T����"x�\o�4�F?6�e��'��Y ����=$���q��K����7p9c�g�fQ(E0��1V���ZȢw[��WD��ܯ'��ۙ�������QQ5X�$q�'\"� رa�+Q���G +�J�"n�.�m>�Q*�va(+gj���C=Ř!G9�ɨ~���I�8�������vG�+�Q�͎A�D��֊cf�� ��^
ä��n$�}{�*pw
��i��rE`�$W��Y���4�K���U��3l�Xb���c](^���Z���1�����>��B	��c#�Rxū���D!�z��E�S]�^��ٽ�P�^��#�E*�_����ˆ����c��S��M�s�	�+����� �F�SsO��l"��(��2���H�ݻƤ��ƖfS�1w���p��v8>�lN��Ѧ��\�����ΰ�׹/ede�89�.lw�3�2�oX^߮r#��-�k ����{�¶P��*�#��r3¨��Y񸡃Xw�����$ȸ �!� � ��~�/V'Dr�)^A�
 �WY����U(�m/��U�եLCj���	N�}~���U��GI�*4�N1S�s���@�����5A�6�l�.�R�P�؟
89�)����$W�������	��Hl�Zh�;Q���cB�Lm�^�Oq�e�t�� �'���n�w$RR
5"�(��z�.}@v!U,9��,S�A�a����P��a�J�ʉeY`��S��g����i;�pr^�]M֚��:e�I�X�)p�NT�K%v,.� ��'!.�u�"�J��x�[/L�]s;#-p�;W=&�]�&�ā�2�=��,�$vׅ4���R���l��N�*w�x�Slڿ��R+�5�"f1T� ����S��B˃��a��k�����;Wу���@�<5�b"\ܡ��GD�VJ��fd՗ �����,�J
��յ�-�%�g5��qYz<pk�_���w��$�����	Z ����.���\��ç���;��IM4��a���N�b���Ƙ�!\UT]�eB��{qw1�x���"O�"�/�{:N�I
w��� 4��!BՖ�EP���%��p����h9�A_&�7t��G�����([��ݝ#�2GY��6�,���~��_a�� j飱H��g�
���an�:w�{��િ+I�ٗ4up^(mQ,.�%Ǘ�Fx=w���	l�-Cy(��9���j�mc����8g�k�2�`�g�^}B6��3��Pہ�F��q�
�1�����S�(�%r���^�Ξ��x��R�=�����#5V1H�S��r	�h��(Vş�!��,�� _sr=l�ʪ ��~x�|��R���S��ه�y�O�v��Hxp�E�J�%,��7S�����(�z�!6���]͸��Y�1�ơ�R�iEW�D&Q&Q3��,��	-wT<u@�3ئ�u�a.�,�'�^)+Jx+o3S��g��W�ڊ'Z�[B���L%����M��>��7����M��J	Jq$w�\� 0�D��-D�]� ���oW^����l��|�?0�16K �^D�fU4.���1!���3D���A��J�Y ��n(�j�@��/Q�g
Ϋ�0�k�$���23tA,�����!2D�3�n��	v����2���<�]��13�+%��\FV�T)N���`u:�o���e�h�◊�L��xI*��B��I�f)YD�ܿ�勴���Omg�=Ǚ�x�����ZX>�$���h����>x*���5�jzi*Kq�ԝo�c٪�\���ٺ(����)?�	o9ˡ�*}f�xy9:B�x=I� hp�uVD��m���ȍ
=�QG�+F�I[ԃC�p������r�j���9'�_j
��:F�ga<��g���C��S�M��!Ď:���L/4{�B;�-�M�494�R�Č�$����&`�;Ԋ��/L;�mw]ƙ/���,nz;#It?[u!�_EE���S���y���S��I# \�g�2�W[�1��:I����1�U����TՅ.�Yr�UT�C�wN5n�����,�ST`�N黲U�\}Z�U0�7g�Ռ$)��s�&�<�K��j�ϝ��1� �����3� T������"���L�v*�4~:�����`p��n w�.f���3%���c�|J��V>Dց��ދ�h��Ỽ������A)�z���
A-��b�H��~, ~ʞ?�����/3�/���<�V�G�5@Z1�v�ث�A*I�/�.{b�m b�ᐼ_J3Ұ�s�p�|��=�"։
��/Vھ.)n�̂���^D�y?s�ޑ����9��oy�A��m}�sZW���@�sG_��.�����J���!�3�	m���n�#�L{?�J�i��Q�%����SINGTѫ.���}[YD�z���$1�u�YB|��p QN�<^}����5(��<a�i~��	/u�o&uJ[0�_����Q.OG���ڐ,�.���v�P����H,?��`����N--|��ڏ]�O�۳��m�=��'b_��4��K�0gL���_֛����4~�m���;N�uC�~�I��	�7�"�����<�PRK_�T��=�W�����@K�`nF���fA���D>Hf�y�ͥ��`[�ʗ"M�������'w�-l:sGu��M
��n���|I�rR�@�H��(����H�EI�{��߇��r���'ϯ�	�2����Q6�K>]4�֕�����d;��l�A�p%����ŜdxA��cX��{p�(V��<F@犱y��6
E:��TgF�V s(X_8���{�������@	�.6d�z��v�/s.�-ђ*S��i݋����D��37���T�)�G˨���l;����;`���j��3i��;���Y�p�+�ꡡ��a�]HqcJ�f���8�d�n�-H��I5���y[\�l햑�&�u�k�m����.��=O�]�����]o�T��d)�db�oP;в�:5d�6��cc�OmM|{�
N*̕��d,�x[Β|gMi`O@�jc����a�a5���B��8 ��л�S��Ͷ! �hPȄ�Y���[t~z���"[�;53�^��D5����\�hX/�3��[��Z��V�)(��_%ɯ�����n�f�l�v�:1����D7	��a~5�,���Ԁ���<3��a��.Y��[L�.���C�B��ƲY<i-�Z(]
v.��Z������Sga[�l������v�:�ڜ~�XO�a#�����eh�%Ǥ��>,gA�o����稼�$H������_����o�ʓ9=���H53l�U!+�Mb#���r<E�����"J�6A2VP͚ͥ���	÷Ɲ��WE�Z�Z�pb��o��!o�A���C^���u:E�H�v=%#jٶ��5����/	a�ʇ�p�^Gk��ex��_�!��~5Y��͕S<���5�K&s~=�&x�u�i?��yYl���E*�O�=��
��o�kn0���p���8'e���Y�s�T��+P����$�f�,�ŠM�Gkޭ� �V���=G|��G܋l�7;'��w�n�=�t�q�,N��ߩt�/�W1��eV?{��@!%yޏ}��R3��E��,0�g�F��-]z�vmj׀v��_���_���yGi��L1�]v��ϿOVr$<�݂f\�s�1��_<����Es���Yƾ����?�s�w1 k@���n��X���5�IS�B{u��z��=U�D���)_e���O*����T��M��b�5?_��$v�%��� Hn?��c����$�Tdd�@�ZTuY��j��1� _�9��V�Z�r@q��0�ҵ�
���`&���eKb�e&|Ϋ���.���|�����,����7�VM��kڤ��]�~��.�sť
�L��L�p
�A�:��᮳��=4������T�@�YX?��|Z�:]��p�$��ԫ�� m"����s��)��/��N�:L�B+�L���i�a�3a���E������W H��[0��7�N�U!C�΁�l;��OӸ�Pr�ع���@�6U�j���1u���!��%.�yv��|ڮC� �\��F�Ǉ���lĒ��/�n�[�.0�&�D�⮙Go��=/ZA�u�.�����|�YV��WUͣ�))f"rm4Q��±��g����[����5��I����y��B$��� �Zĥ��C��Ge�e<Q���󬀬)�
�'�Y�wQ�:��Y�������'x�}�C�{�]�6��<n<Vi�j.��Z�PE�r��ꂺ�T�ǳ���tP�ûa	�����|%[�(1�2�h�0�!܈���B�wS������+�{ڠ���t���Nc�����][A�wm�F��r�~VC�	 �O�:��2	>�KLS�9�m�֥�.1�HVx��6�)�%0���Hfgt�:����� r�q���
lG�X�k��.Q�մE���l�j��3B��c�����8�3r�T7�$$����M�>$�4��h����)�4�� �ţ8.�CN���l�r�wz��Zʂ)-�Ő�/�A�"$㌏$	T1H�1zjN�i�9$��'ΈK��2�'�W?W�L"��Ħ`����jU�鸆�;ћP��(�p���^y��eE�_�d����rנB��ϑ	�T�~��V�/�!�P�@1�˖5��4��4�HFV��������q���ok���5�OT���z
�6XB.l{��$��@
4��h0U��fK�������7�?�|U<N�XA���#I����oʰi��4"��@5��?�3�x�|��qt-���?�C�p�,���;�iמG/���z��}Zڅ=K�I(�8g���i���_�����^�Q�!�p��֥�$�ǜ�i=�Z�!Nͤ?��)�8�4�wO�D��Bub����N�^�G��2[��{����5���JX��pJ��D�?���r���{�b��Er���v73lC����em��=$M�Q�[����'+}ڟN��\�qd�Z�~�9�fADU�1�&� ��`h�  ����3&p}�oy�S�~tv,8�s%�Ԁ�*%�k{�i���XmI���D >�q\��g�';��+� ��m�o����~���bgY�V���u4��D���`���Ё�n����~����=Rni���Τ࿪R�4��yX7��u-���������*$�W{�W�PT���J�Jo�M�0��74�T�a2$\&��?��h�T�g�$;�:FWpK����Ը��L�M���|���7�SB�ƨ��aE�g����M�g�R�cl�{C����pABu�D�&�|�A5)U�� QN��}�<�΂n��c�if��¹(
ޠ�_���cvԿo�w��|(���h�7/m �%I�!�5{[J���d��<��0k�0�jy"I7�*�?)�Y�E���`���Z�l!w����LV�r��f�g�}�s����D�����69�|';.��Z�׳"����@N{�M����h6�H�N���<ޱsbQ�P^���i��.W��r�S���_����G�Z�x�8�R��!ȸ�Z����}�եs m���A PF���ԐQ#��ج:�<�p��O  r�� ������
�f&�� g��'�t<����ŝ�,�Me��ז_ؑ�.*i3��ۙ]��cId�#��phu���v�@�s3�BL�ٰR-�rw���!�K�b���q���e�Xx68ܣ-s���O5
Xs�L�:�%�{!!��b8���\I�1�W��S�V
�Q�	}�+���\� m�~1e$<�8k�*�}{��Q�`�/ ����>ck/:�g����r;)r�e�3�ȇ�����t�<;�4���������w��=�,af������W݌xK�/k���j�v��}�Vk-��QA3W�HO����1�ױ���Ζ
��Xh�+�_u��ʬV(�� �d�ê���E/�(�yx�u�8��]��^�o*;�b�A�|f��?�}�ĥNC�/-*+���X]�c|V�@����`�}�32Д<O�Fk~�	�O���ڷ�x՜�+����ctԊ�8�����������*��9�!�%Tһ)���f|7�is�����*�e_a�'���5[���ćȡ��t�HJҺ�a^m2��&h�E0�2fS�!��Ì;8�|k
8�:��oW�/<(��о�3�"m�L?�`���,ʎ��`X�C�p,F�nGV���1��s��V�
C�Pfú���;����%ZL�d�9K�^m�Ɨ֪v���H���[*?03~�{���%}���!�US�+���G#��g�Hؑ�檝�,����] ym��	���;%���82�E}��gN�^�����N���E�Zbk+x�d�Wᑎ��l��w��\N�?�z	x��hխf��A��4	e0���d����v��?e��J"3�U����4c��ktZ�yu"��v+�1��l��!W�s3j����p^�ɲ�M�42 �-J�Օ��I���p�	�pܞ�6��$��:q(s���~����o$p{�Z̃�t�J� Y�r-����+�]�X=����ˍ���eB��o�N"�Y���p�C�%��;!��ԏ�����i�ۦ���S*��ZAj`�K^1�
@p�CD[�I�0��>=N*�d5�T?�W��ԭ�_]����� lć��4�F2�$�[��Q�ER��p�����r�z}a��<}�.��Q;@�?�bX�TZ��1W��T�]���_��C{L����e��`צƩ�1��#��X�Q�H*�KQ����\/�HPU����[��LB���ѓ���I�v/���tO��<S�hh�h�f|�l➩�v�hM��m�_���RkO��ܾ?�Hכ�~c �n�!��i����~C�ҡ��wu�E���uV�*��[(�0�e���m0�9*�s�nUʫ�LA�]זו�D+a�����-q0=�.��~ydؚ���IQJu�bo�$}B����0o'}�\�kU���',(�L�fT�/Х�R-��i�l_�J�7/rE̹�4��b�S3�D��j���#�y.WA���$N�P��鱭?6[�;C��z﷌�Vp�5��e��>����:.��,�!-�����ܑl�*�Z�C����4�?}�g�~+9�L��=z3"xl'SK�����Z�н��{��=��0�w�����'����N�3�� 6%
@u��2L̙U�n��ҁ�I��wh�#�W��QT���Ƅd��D�a7�P0�S�a��S�k�χ�->X!{ϼq�9�G�T~��9:"#*���ع����X�W�Ĩ��8���:ku�TV��]�7�sn鐚����Ƴ�q�����/fb�*�Ɣ��͜)�N��1�������G�"^�<�!#ɓzn&���/�eਤ<��WV��` ��٨�ו��>��7��!�cr�@+��(h5��Tw�>3��b�h[1����>�`�,�'��^�����>v������4�=���<0@�
DN0��9P�1��d0_O���
3f]��ڻK���i%d�N����}r>BT��hp��]]`�U����0@�+�����o�N��Ҵ ӡ?wt�+��*H���l��
*7�n��ܵ5�7oʮZ-䲈�O�Qozk#�"]�����=(�3����{Y��i
ԃ^W��p4�t�
\�򹠑Ӭ���^$�J�3@����Ԁ#\��ߚL�;��-G��ry�������ş�a��3 3��x��a:������n�}LZm�B����t��!)�ۄ��v|u��RQt�:�*3a��Bg�L���� �{Oż�%]:���)���p���h���2�����3LVRŦ���x~.�u��r�Ʉ7L!7i=3M�l��)4��I�6'_�k��;�:<�V����R�#f)D�\�btH^ғ`Y�*���$-���	�R��������-��\����0�Ԭ`����g��|�L[�g��:���CO	j{�ce��NIXe�p�����(�W����R�ȃ�$�`ס�KZ�d�]���n�(ǆu�JIF�Q'1�I��nt��Lf�P�^���Ő�\���Ò��'%{�%�AyNHN������%y���v.fa6�-k���M���t�4�����Y�86!��988�x�����rx��J��Ȯ�������T?",�L����7�LdZ�P��� W�|'*�4b��u^o]������ ~[r�ؑ�~�'���{��Q	iI����8�gH�����}X�3���}���h�7K���լ'�J:�U�f���㚈��;3��Ր]*<�-e����!��d�rR-�7��M��r�f%sF 9�qR�<�����H&&�54����Y�ZG�j$Xr��E�e���Ȃ�|��ܽ�(�c�)�T����Po�f�����Q{�������v-��$b�2���َ�����M�sq
f��_�l�v��*�z�F��!�J꽙hn7X�&A? HL��rĚ��-&	OF;?�p8Ş��i"����h���z�}�Dq}��QNū��Avu�0D����z���?��e��w0�=��
�g�=de�>��o!x0�?�+ɇ�<O7�����;-��%~��v�W��N>3�\;�78�]}��!��/t{K��#Ǡ?*\Z���!k	��=�*����b�`Z*�|#Nvt����s<}M��_�����B�+u<b,�0> XH~4��[=�liGTj��g���g�z��I����r�ٙ^�x}l���G�L|���,��O�A8;�*B��R�p?u����.p'��,9����@���Lu2^ۑܢ}f��k�G��u��7�e'X�5(0�JXM$��Et�h���2��;h��O*�(M?�u'�ՙ�5���Ԫ�����^�B�)4\PVS�	��wf�f��Q�ƌM��xܠ}�h	��x�,���Z#���rs+�`)M�~:�F�mt�1L9a�0�b��q�q�����y�d��>h�2N�Z\X�~qG+򸉬ol��Q��K2�m3�2���~u��J�F2���Y��55�p��i>e�I�}�D�p�B�I��O�y�*�e&*��,��5�fh_�� �$����w�Q�h�S�;?�?= ��l|)޳�=����E.!>�kaDo���h�r.W�*�xsڄ��t� �<d����/ҳ�'i=	�sbD芫�T��(�lǾ_�z�`6�O�o��'�M��������e�/
,��v/�W���b7LU�} ��
�FM��9%?v�G���1�bkj��ǣ�n���N6��)�Ň^�
@C"#w�A ��?Ql����UU�8�i;��bn�e�S+��ɻ+J������p��
��������m�;`^��������X�*�e+s��¦��h!�ڈ诅�8��8�1�A��l-�W��r����":����>� <X�%�?�1�MNU^Udi7(����e�{
Ν{J��x!�D�?EZ�@�O�W���d�*|0�]��9'���|ơ������j��;�Q����đ�){��F�+�k%��ܓV �K�k�A�u)ۺ�lY@�{�R{�n�}�z���BE¤��anqZW[�v���u�vg4L�[�v���O�a�����'���<�Dp���q�#Y�$��c�°2���A)t�뻥������ ��z� m�s��f�&���Պ=�{��ITO�GnI����B�6B�Hã����mc(�W��g�� ���Bp�|*}�$��I��gst{!{*�F	��s��n������F^�,�]�Xf�l��bU�)��jR3���&�7� �jv��I�&&�@�������E}�'�iu�'v�]y��R��sɤ�KA�2�ISW͂ �\Ɩ;b��b����x���X_u���]i�����/-���\z	�[+�z�c�K(�Y>g���o�O6��̝��0�f��: D���tQ��o)59�&�ER_y�����b܆!���Y�,.�#�aY�p��\P��yCڴ��&:n��\�uAd���cw�b�>p�y(|*����m�|�y+�XJ����������+�w�>���ٛ|��Ԟ_%�b4�#�!�H��zdq����.$٣�	��ßu���G�C�d=��O��Ӊ*�}����6;W�(%�) y'�һ �����!f3�xʾ%C��]��+�	��s�\�����Z
%$O�lƔ����V��6MG�j&`�9�L����K0"�G�q[��٦��{LH�HfJB�S/��uwG/C��ۗ;��q��H�"���%=�"&οsg>�����9���:
r�=�/����Oʍ���$"������c�
=s���݃�X4&��e�G���hD֓��n��۵������]�-Ԕp�@�F�م(�Gv%K[��M��H�,�Z����I�֢~:��m��H�q	�$�ऍ+�1�=�2K����<�@*10CW�xBB���VVM!'�sd�3���Drw6ep����\b�6ܵ�q��Z@��	��B������_z�h�EW`�e�ЖY�G]{�䶆��@*�K��{[[�-�]�K}��1o^�\1���MP퇵=�NXĔ�7Hgl��I �dI�p�4��	�ם�k����~�0��dϼG�P�ȻK�Q�}���Z#��L0����*eqGpZu4���r���A�'�C���ih���s���ſRwx%��qUK��_���P�����3s���I���w�����K������!���(]�!��c��YG��kK�nY�ƊI�Z=�j�]>ic�"l��)����P�<@G���`ǃ�M���UÈkXFL'3GT�a���۩���qA:5h�i$aT��͞W=t�#����!�Zm18�CvڗB�hO��o᪀�Ve���dZȮ��H��i�������QzopxN<n�rQ҆-�@�߹�Y�WЍ�S�W��q6j~���W��BN�?�#�J������D��D����Mpq��շ���0�78� E�"s6i���f	a3��6�i~#�_�����|��Y�S8��j�tY���dW�o�2wÎ$����~CL�ͧ ����0R���HJ"��5�>��2}��}==/�D�a�+})�	Ԍ�[���j鹆��p[c è�X�N�����i�E���{������ՁD�;��UW��� ��1�/���r� 7���U�p(ua�4��my/�x������%���jW�(i�B��f�xd��j���5dϘmN
~Mr��F�%]�ځ�����P̈9˦^���6Ku�U�1���W}�4J\��s -vs�	�Gs���:K��sHey�*_��`���6vX��#s��B޺���4�9O�G#;�����҆D�77gCe}��0�AB#[ށ9r�z�l���J����I�|��)CmauQԲ��g�b���HtsK�)���I�>�� ���q�C+�l^��]Daih�g��v�3�p���Hx�c��G��G�8XS����)�E�(��uz�K��q�30��E	���Hm�3���Qʝ�m���~��w�v�%��R���ο�Ĕ6��m�}�I����w�{�E��VJ��?�ul+�2 ��x!%���T5B!'i<���di<.`��D�6�y9�� ���g0���j��c�@:�5d}�L�޾�Y�*���M��42�ur%�ϰm�;i�8�N��7Ս���0�v���6u��48�Dwh�E�*�����JOي��.��q�ˑ}6�r��>�8El��<�E������ )���/��1P%��W����Go����.��b�����R眱i���x�>H�T���ũh<R��m(b�fA��M����&�8�����@�B�8]j��bh�U��9�ރG���ǺI��F���UЃ8��_�����q1o�������B\���8hx� ��`hs�)w57��ͳ�/�tH(�W���J��VߠR,q�>���\[q�[f�+�D��`Qg�{�6���W��U�aiz�>��'K�u=R�M��]�oy]O���P����FZO�"�F��:L��0g�L;��Q��>o�e�A��&���=�J��3f)���U9���=Nܳ戮ONFg"�n��ok6VS٦88'6]�OvY���֓4K���9W�p<<'!Ϣۈw�*���L6���;�x�^��]��JF/�^�A5X�����Z��}h������H��+P��U��M����Υv���r��ႀ룋u�Od��m�BA�]�^�R������vyɀg�y��M��T��n�XU�4�ͳ,%T�)pG�TȇÁ!�$��0����y�e�N�gg���7(�J7��8I#;�Y�YqT��`0o{Z�gt#%�7��X�6��u+�i�l���z��4a#T>�v���fV�0c��N�PĮ;�����Xس��۫;\�֛4�o��J�Ȼ�]9B!-~9|��/�����O͖�9C-�ޞ�)����u��
Lz���1/qS���xθ���x�$��)�4�@$av ��:���1���%#����}�DP�_���tG!j��ϕW�;�e�E#7���6 �[���Ф/��'�GO�VLBj�u���J90(��IG�U��@��K���@��Ufν��D��'a&ǥF�]\3�r�i���U�ڂ����A[���*<uMj�oj�I��ZA-O��"e�ɿ��ydB$J2N�:�v�e�(���2(:+Լ��39�Ed����N��)Ǧ%=�m�5b��y�ެ
���1&>85N�b*H�0W��	���O8<q��H�!S� ��f�[��yc�4#����<N�����d�R������֣W��Ԑ������ �uM�q"GQ�L�0B�.�&%u���TѺP�^�t�q���9Z,-S	�4]{�}�غd��]� �X�p���c��1-��aƜ����2z��a���#j��e��Tb0�!,e�q�f�#���9�8 @ D��_�'�6�,lj�Ε��F�s.^;�ǁu��·�A��s�:-��07���4��|<�#�t�Or+���B�e>, �i�g�������h�����1��M�������{n�*h��OB�� �<z���}Y�,\/�B�*�o':]U(o�� ]7�kU��>]�~�Tm���?r����O-������^Bk#�^s��Djm9�I5�*N��en�Dc m�Z�|�$L���!��J+�9��������d0.�L��!�@]�������u��<+�V�IV��9#	,݄����~?��u���Vڏ̥C�]�jGoWPrS�׫a�b4�Xѵ��Ҝͮ^,���X �u�ӽLך�j�Vj�𳺕gH�+�5��Ss��ڠ#�/xy�Y�ѿ�vsXYWQH�v�v.��֩s���K�T��\��	%�F{Ii~�/��#��Ѹ�Ɲ�8 f��-~d�=v�V�������r�I�Wv�#�4uXw	Fv�Glt2�`������|��8���8��7���弬�C��,�t��Ń�r�����P���AƊ}�-0�n�d��c��a�P�2Ci�t~{d�pv�:�X�q�9vJn��J>��Թ�sx�j�;�R��5�(IW:�Y�28��P����9	���4�h��)�`}���gm?��t�;g��aT���K�a�����]*j&X�w��<����ٕ���0��n�qZ�M��#'��Il&��Yq�k/t���o�>}���js!!a���1Ů1w�]5F�(AЄ\¢��7k�Шs�;�c(1� ��$I,66���NrC������p�|�R�Nj����'�ї(���'�Z����By:�m��50e��H%�w	�Q���b[�v~��_ .j~�Dz@f}����1����������N�Mui�������D�`��:,r� v��Y��Y^��w��U��O��v�5?�b����i��g���R�B?g	'0���{�\�f}�Ĵ���s�"w�~p��>�U�SY]x:k��s+�O��?�qb(b��\K�?�C�o�X,�BiG�П�Pv��� Oo�����˔��)D3vڍr����c�%O��yܤZ���g�/W<��\ ���T�4,���������8��V��w��@9M����"�a�C!�S&��2PJ�
���+B��8j�	2�#��� �1�Û���M��d��˩�MH��L�7C��'��ĉ<�� !�t�}�Z�&צ�s�K�B�lq�w��ۀ��EzuO[�{ǹ�O���o�Y�H*/!�#�j��.hTe�/�(֐�\��GG��U�����sV�_��z,��A �t*�;@�^��t�U���v� w�Y�Xύ�e?l7�*��aZ�����|?Ԏ3@[���z�3�Ӏ�� $����>������Y�._�B�4Źmh�s펔��qy�y���1)`�PRM�Ǉ�i���4���{J�f
qAZr����!�;��!� �M��K�����"�r��N��/Ҁ�f���9Es�_��Uj��aH�?{v���������L� �4y,�e�Fܬ���e�K�؞�ُ���a!W2�CO}��\�����	8�0P]բpy�@k�[������uM��<y�R�<D#φz��,�s�S�f�$�08���
}Z^���Kt6N�٘Au��h��<�E4~KNn�Dp�����y�?f�I4��P?,�g������.Z�����n�8%c�3���4�1�����1D��tV;�@���U�r��5M\^���I@��n&�zK?����9X�O�{+`�E�b�2�Z|r�c��'�dԭʓ	�Tgk������E�88g��w�f&����G���S録8���v
���rw�V����y!ƅk��{��ąՒ&����;���l܉���,��H�
���f���<��x��#��rC 
D������.��K�����ԓ�m�U ����)_��f��*ي5W��D`ճ���Q;L5m؏I�O�a�~�f���PV��%�.B�/�������.���ɩ���qа�V�e�y3�d�;3�_��䖗�T�Y����;�?O�s��FzO�PZ��iA>���y�H!v2U��[������}"�}�dCZ�!?���?�V�B&G����u��)����j����z�*3�F0�ְ�&��Q�K�I�'�ˁX$O�Q�h����=���ňNP2؉i�ښ�+��96@a����&b�Mw���&q&R�A 5i�N>�1��BZ�~�
�f�Ux�� ���!I���b�c:��{��R�:jٖG��k�x���]ϰC,:Q�nTY
�oh�ܣ�U�*^J72���8�@_T�}+d�x_M�RLy=}�}a���6�!R)	��gEq�����:��[0�"��h"��c�z���kx7�ҵg\glp؉�y;����$j�(!�H�Ё�[3�O���{�X2�C�6 �A{�5�({��Hi/�Tɻ#�^.�/E���B���l�b��֖��Y2}�f#���[����?fN թ�}�
��Ïm�0�4s^�u��	�y�nM5T ��J7��<Ӷ7`sS��"b-�ra	>�������d�[����t�Ga��ȋU���n`Ӑ�����R��l D����&�0�:X����C:�Ճ�4���.�b���fiZ%A�����_��c�C���!��Ryz(	����c�S��Hoyk� �S�(����
�����	G�|@[�f!�t�,�N�m�ύrƠ;X74����f�)~��c�i��"~Z ;�@��4�C��C���×�����|�p�i�2�W�4�$#/q؊�|�4ܝT�@�Ih��)��\���7����=�.�� ��� }��e�W�t�Y��Fka6��'v�-��y�n�<���G���
t�
Z$8I?�V�>F<&P������E��@�h��O|���A8�Bace���o)o;y�t��G�eLy�o����ˁI�9m:��y��l�ib���$�S�:������Ԡ|��تĆ��'�g�iH��r�����h���!�/,�zˆj��	��>װ	�l��,����O }f ���=XF�4�ր�4N�-*׆�ʩ����"�1?����X��Qo��8��n~G� W�#��Ͷ��$�l��Rv}Nbщ��WE~'�I=��Q�x�T��P:��=ɪ��4K3�c�3�e�OOTM3�dnIc�2~����X�W��*���o'2)#����i�ҼKZe���|Y��+�/�t$�=�#�m�#�*eن<�4���h�.���u׹��_j�� ���F���
$Nț���b�_�i���X������D�X�8&-��N3��b���D}��p~9I�~=����zr����j9c DF�������F�d��v:U6��!�}���J�����;Lp3��k(��+�j�k�B�n�-��:�Xc7:���ړN"�2qZ@[ǲ���J�7$rU����PE��x2Kc/�?�ü�흖ʴ��`���m[Q��)��A�R�z���Kz�+��(ǻ�gՀ��5�)7 ���p��:��4�oNr���ȃ�Z�'.Z��qȖ3u�A	m���c�o�e������^� 	���㝌`~D����}�E�Y�����q1��	��LCH@�m�m
eE��dA�r�13��Bo#SE��d�t�}��:�o����Q]
���V��^L��u���C���\�@�4���qߦ���M����YM`@�������0�	�`�^��d\�Fo�BV���ZtR�����f��k���K��-�O���9�J�'�)��ْ-:MZ�-����򹬽�^��$q�����3�/��J1����\�?1�u��r��43�JIխ�9��es�T�`�co�#eb�,B�wcW��@�^�趝u5'J�^���-GN<�O���q�V
�m%G\�Z/��b�y'V'�k_�=!�����cbhzH�h���� 2�b�|#�d3S��b�R�V��\KB���H�e�9R ��Խ�j��r�;Y �M���lFu�ⅴ���|�$���4�8�;��|�.5��Bv���� ց6��MJ�5m10q\���}�e_1]E�RK�J���:��kPK%42�)�E��;�Z�XmA��,'�E��� ��ň#�C�xk��K�o0����x�v�k�:&�V�������C1���pߒ���~����M9�+��՗�Sx�0%Z�����I6a��T2�I]NM� }|1�K�!s�3�'��� Ç]�M���!�@w�m8�$���
F��~pe��D�.u�B�Au�M�E�&��x�	l�v�66^hg������Q$C�~Ox����o�wC�o{�RB�Y���U����}� Q8�H�͡����X<1�a��L�X�g�U�W��޿�T^�ve>?~a����V��D��h�$�t ֑+S��Zi���bb�������
�����Je����+�7��zM�@G0�S� �� \<��\��1u@��\M��)��z{[�Ў: -�C!���!3k���D���%'<�����{5!�+��3��v4�w�3H�1O���S�_����K��zD��f���h�-����B��^���nqvll<	Z�Ӌ!�������GL7� E��1�T`���xޗBA��`�'ī�hK!s:,�������]]�w^��4�[�����?�}M�д�#��f!�ԑ��l�g��:,-���F����DZ��g/x��_�|��ON��t>�^R�x�Ug'~�|b�-�H��;1��v�������ɼ۲��`���G�����98�q��2�NB��b��td>r�$M�%���D�q���s��,�޺~_��c�2h%U���{eO ];���I��hf�ٝ9�$[Obl�>����u�V��7u��H�����;��Eµ��M"��S�G����F���QY0�2:��}�8��4&��{4��
c���TC�E�+�����p�[/��7���jTyZ
w͏�C���[��G�u�%�-z	"��3�@+/߅^$S鈴Zv�5�U	��I�XL�6����V=y]�5/ː��}6�Jh1kW���R'/q�l��{l�눩�������Q6�/���_��?��`s�$=�H������Kb/#0�PR5b$d|(	|iU�e�F`6����]n3����M���b�Nꎿm:~�k��i�SB�ǹrc���.1�Ny{�:E������捋�n�w��x���jU�xV��^]��.V-oM\��?̓4���{�$�mG~��Z��_�J�zm��4���A�!Y�|�zg��Fv(0͠ �ѕ�Mkd�~�II�&� ���݃�8��d�sǟ�_��h��Ro���%l�D�6�ݿ��K�h(�r"��-�|#&D���BR)�E`�e�ȯ�9�%��������u��Xoem�5	���H��8'�@'؍�4|�N�;~m��]U�e���wl��jz��S��&�	��ÁdGj���P_-[kޝ�z�½�#�����@�_Vi�KjN��r5������Sf=1Ia�Xhӕ���G�g�x��ΫO��!��}���^��2Gd�(_\�V5��.�︦@0J��#+� �����Oq!'�PGAQT��z��Gʉbg�s�P�C�dT�[����(�O��y����,�U��ho�W�k����&��xr��OXU��!9O���^ڬ,*h1�Ҷ��^����3콌_�#q�$�gv��x�5�?�+x*���mu�h�]A��|��3;���f_��O����O�k��)%��V���6da�"��K�@�:t\��`p6kc�"���ͤ���p���!�^R��Y��c=*��mg��R9b���ׂ��{c;����	��bk���bG�'8I�(��\K�I��:9�#u��o�:|е�\_����髦=����=����
�q�����E��4�h!]q���G��Wf1U����T������^��[�c:p�@Y�G�i�����K��$�1�Ej���*{a���,Y��1���k
�mI���|��W�qk��t�����Es��T#x��2X�z��c9�d� �7<� a�<�����]>k]����aX��r����W�'�$����X��X(���(�@>�`C���L_^;��o�C��H�қ@���M�d�Meo�o�yߎ	2��Vw��F6��t��A�4-Q���_`�~��>#��9X:���l��(#���vE*�F�Bߏ���u�;�j8M����oV](��@c�\�����	�m���L����ln�Z�\	�aT߆��B���%�SŜv-Tϙ�h��9(k�}�S.�ӗ�.�+JV�+60�>b�g�CجppC�\��t|\�L����|�����a
��Ќ]��\��/�5D��-U3�<	���p����n�3�YFìоs�w�>,������$�쒒�����|M�p��vx!)	���JSz�l(H8.%I�ݦU�{Cg�}0�u�fL�g�ZA�0�֗������"j*qKxXt��i�WWX=��H:b��j��e
� �V����t�p�_|��1���i�
QpKg�P%#F��Ʋ���6{���R�4�U�\M���}liq�WP@��cyC'���O��9��(��NM�:&��o�<�c_�QŪ{�kd��uϋqN� ɺ��t�A�ʸ����ECٶ]��`"�!BC��9l-�Â�AC����">``�[�v%���rMv4;	�5L�-F��hfe�bx��.�4��"W��@uA�&�Ȇ�4��'����GM�³ia�[�y�$}�A�%}��5��:
m�Ma$���U�kк��!b���D�,2�0ͺ����u�o�Д�|���rq��oΝ�l���Ȣ؞Y���9Y���0��tM|��T{H&ᑜ*�~^���͇���$��y*o=��e�16g�փ]�誃`dٓ��71�>�X&(MW>@v���t�=�=8M:	���>L�}���ߘ2�����x��ܧ��{ʌ�0��%��!��Z�2�#Ċ���Ȼ�T����m�^�z|q��������9���h��#�H?ո�ŕ�D7�?�[	X?�L�Č�{�1���T^��Jc|���[ ���Kn[I$�N��!C�~j\4����^��	�$�I��b(?U$�f�@j���H�|<����+�[�l��3p�I[oԻ"���a"%��ĩ:Λ�����?��q��A\�I���xE/D�8�y���]ׁ��D ��8 ���#ek7�/�U�<<�[�g��0�|������{.]��)�m�໔x���o��J�ZY_�Y�X�K���[�(xi-���W�f�fXm��ysH�>�8��g��/��e��i��׬��K&m�-�f��0����>}�Ħ$�f�3wg�EIK�o��R.bu�x��*?�> �P�M ��m�įf���^Pw�"W�Ȼ�2ڔ2f����j�'���#� EAF�63��F~&�[G%���|۸���;�D,f�+�ó)�ݔi������N>ob{f��6�ɚ�kl2�]R�Gw�\�l��PS*�������\J+(�s(�@Ymʊ@��L��),K�{X?��8ʅf�HA�`���va�S�"�N��QJ}�Ĕv�qy��)����!,Md������8�@��VR"^y!�_��vlb�*�c�j���>���E�֫X�<W8�2����I\�&IG�U5���t�f0�5�!���ވ���pW�	F-Yгt�9��B�*��1�Vx,�N�"Z�����g��|f����AZ�D��<�f�P��8�ɗ�w���}&�d4͸��]Fh0����률q��\�<w93��AŢFnR�(6�
EG�<����UA�����~�>�oˁ9�g��\�g�����<ζ���L�[�r<c��,�	��hN��$?�E��&��u��F��R�{H'_�����S|���3
�����b�y�-
t�
���+7��L��opm�iom����O�C��>��V�������ou(�yl���'�ty;�Cx1���C�P��}�� �ŸG�1��q�5i����%v2���I��h��
%�������e �|"`��w����j#�㪩�iǢs�ĴH�^�y�\���+Q�[��h�X)&X��K�{��^0E$�i�*��8-0(��2�p����e �S{}�W>����=ߓT.1U=|<��1w%:��ݭ�'�vU:3Ҳ���-����'��i/%WNB0�/��XO#7SP�@��
t�'$tw�Y�{3Y�P�R�Z2��w�1ǋ�"7����"�4��ټ T�V�]vt���FD�kv�t0H�E7פ�F�.��V�/p-��øa��MŶ�'�h�cQ f-��#�Ӝ�"]��@�(�GNܘ�33�����J�|ޟ��&y�]e)&�S	���+�L�U�	q�by�	2*"	t|J)��YѠ�ٚw5�B�>!�%
�r�̟��V�� �PXrM/{W�#W�S����,����yQߍש0��F�#��T��x�����$����C �ɐ�,rB#���e���pr���l��k,<�=�_V�aT>��~��GKD#�ɦ�
��`H��ӓ_0rڠ���R���TZ�y`�oI2�`�|����P�^+�MV�{z�ŪL�m�E�^�}�B�����x/�8Af|:O��gOMT^��Y��s�|W���i�o��9
���=��� ��_ �1�2�ѩ��%BP�\A�x��;-�����_�����T��vlx�w���; ����yQ�x4� h�@a��:�ch�=����k�o|R@�'�wO	�v:!���.�ع��������zO�j��A���	I@�1p`e�۔)ܲ]��u�Q�
�N�4�)֎��
��+X$�`�:%˪z�Q����Q���ӽ��L�35T�v�}�$��L�@��C�?�����o�x=8��.�G3{�L?�@�� 925`���!e�jF�֒�����O?}�ũ#5c�T�! ʓ���lք	@�(|WB�~��Yc�$�������b����DOԍ�Qh��&��"���s�e�����	�m	�
��B�4]r3G�fC*�7�"�]kQ|%u!������;�3� �k�F���[{#g+y���b����#Ы_?�B��C�#��������J޲uH�|�dj�?L��9�u=}t�	S~p\������r��xQZt�򬋊�/)T���,AiS+X�m13�����K�k�S�y�#[{��}�ףt�+��l�(r-_���V��}��[|����j�#���{��1�;}��$pL�Cp�w�� 9��vs�.�3�D3��������b^Ak�[�ҵ14Dܪ*�r��9�������!����+W;� �#��
��l""���]'�R�#)�q\B�m�y�Ɠ���6&G�e7�Կ4�i�o+�S4��M29�;�h9�D�%��N��ܟ;���H�]�޿B:�L�,�-H���"(v�q}_��
<A�h�Cy���F���=��=�m2��å@�e�2�->�9�3� X��]�r���A��Y� �ĩ=t�&�z?���b�/�y+$w��y�;���i~#h�p�4#B�{�_��1�"�!/mK{��������3�7���%�j�nb�9�~�q�
,��YK��"7��a����cER=4��Q�J�ޤ	���L��ֵb�	��j�Ks���]�q(U�?W��!o=n�t�/�������c��f��xd��yܮQ�N���A��8Կ+���>R�4������٠�g�$'��>� -?m&�|�Q�f�cseN��'$�]��8S &#��'p�E~��o��R��AH�+�����Mk���KWX{Wy�R��|�"�˃�>/���mSjs��i��B9{k&�%q�߂�b��x��`:�.����/u�!��z̓4��P�}�98�z�<ֹge?c���f�����x5zU�K��F�IZ�khJ��	5���]���90Q�9.�Ú����e�B�]��J���_�#�j�����x�|�0C����o_�7���w�l_!��#0�V"���,�Ny���A ��S:����b>:L��d�~.@J7/�ʼ�F>�"�ʣ�(�b��9��
ݽQM}A��G87薶,��,�K�����l�=��+���.
+��I!C�m��4��փ��V��Rv�e�@G�gn����*,�a���0X�0�	 ���|qF㔟@���p{(#��W����2�� ������1i��X����\�w�s�����Nô����и�53�D
w�]£V��H�>N�7ծ0<Dr�	ƶڕ��&m�}o���v�[Ŧ�Ӧl��w�(�Z����t��d�ef�4o��$�˄����L�zh�:`�0�s'��!Aʕ'K��p�_RҴ�B��	F)`����R)�y�%Q�Fx<7y�R��?&8z����l��*?�8�4@�����?���s����t"��ޖ � ;�D�c�������^��̙Z˛�C������'��@!��L�3�r�%�O�Mwj����J�ֹ^����G�X����@�a��k��-�����\��A�#/�����/.�}�4� K��ڍ����
Fޅ�4��@�xe��f~뇾*Ȓ�k/�Ñu�oWЅ�0���9���z4Ϋ��:�ѡ��؍'��BV��xw6�-c!3`�e�A3�ѓJ�x�y�7D��B�}�g?��	>��8����u��Tk���0\�y�E��H�3��4����a��;nҹG��fh��ׇt�u�a�S�$tz���v� �%�l0�
�5��Ol��a�F�l,�;t��}p�gO��$�7�����ԫ!�Ի���ʪ҆TIөvv�I����|ʴ�{]���?~���h�X �jy��+j����DF�����!�[T�m3?{+z,M1.���ׇ����\a� �Z:6��ZB�e�˒�up�O;>aɣ0��#�B>�5)l>��CL̢�vvS#�ʦ&��w�0j���M8�/�����fłXS��c4��PKQ�6��� ��;�p?Vy��(6l����QIC�ɬ"�ċ`I��?��es��Q�/Jm��Š�?��v�N��<h�h/X����]��m��P�
eI.���ּ��I��W;b~8�{}����A��(�`8*����$2�a��B �ߺ��	�2�mGl���>!b�z����p��!��s�g�T�
��#~��M+L{Vz l��BpOXo8y���{�ZV��*%M���۬����8����#`b��q��l���i�'���
+N�UMC�hH�U�Z�+ ��[��K�{��'C�hF����%�"-BR:�����j�^����(0G�~6�+�������^����Nި���'۝����AB.�آ ~��c88��p.S�5��ӻMK�9���ԣ��퓤2�d��SsM��
��1mK���/ݲi�c,�7Kǰ�R���	ϠPGA�/�;��P����IUx�*��R��������Cao=�#K�~u+RR��o�!S���o�?j����"�N,��O|ղ��Y��&�2=.S�[�Yu*m��P}d�r�ҩ;�&����;�Jx#r�k=X8 �ڧU3�Y�O~��Xg.�����!m��$`��"�a�~�?�r0Q.|���+}s|ru.o,ս��}B.����Y����VnB.@��4�Z���nZ+7O��'
�c�<;A���y���dIUD�z�=��ކxȹ�[�s�e��
��c&�N�R��������,َ\���i�A�Ie
5�&>����ӻ�'���Ŗؤy^�������ӛs ����R�|_��o������R�������6܀�]j] ��=v����-$/%kH���/QCH.��}�Р�r��x�֭A������?��Hag5���B|RQ�8"�_������F��W/i����H���΍m
ȣ�X�)u��\�V������� ��z�\�_1b�ۦ��dkEN6٣�ʂk;XHd�3���t2�B�����R,���*�C��uiE�]��l�y���R��r�$�8�,���˨4�yY^�td��z�g��e�̬tNt�Z�n���k#D���wD�oR��5r�� �����2� �d)�:P�G�P�m1m����MІJ���9<Y{.���f^9�,=}	��Y�������C�옷r��w�i[G�8^ĕ��IQ&m���]�=᎑�<zLփ���S�h�ޟWs�pVBT}
Y�����֥�������w�������hL,A���T�������$Hc�*�n,�\�1F����F��_��B�e�!�y�����oVm*��W�NU��&����=��꯽�L����`1����h�<;�z�%���(*<�Y�%�d�2'Ëu-�oѪ˰	D�<$5�b���jop�d^yD嚮zψ��i��@?κ߉���,�Cc{����;�l�A�C��>��T��!��ޢ�W��6,l��U�b�u3��0L�T}}-����c���ɪ�Q�{�6�Ŀc}Ԍ	�M��᫪������Za&O蔗a�����)l�Ƌcf��8q�,[����%=zl��^/(<�p��e)����X�b��$J�!!�v�q^*���(f�qy%���6WP��h��z4E�@=�h�}Wb����8C���<�;�0!����0�r2YFf������!��2�R�i�P7��T4_���i��q�$�ڈ[zR�46���&��b��e�2��ۜs����ZF\���wk�G?���Խ"����T����p_�jZ,ЄC���A�<Rׄ�6�ɺ�LL�!_�!+��bv224�U�@rs"R�̔fʑ�gK�u���� ��U��Ԯ�?�\NE�H����t.{9��	P0P�A�8�������"}�q0�`ٗ�f����������eyN���=���F!&�����CP/����
��0�+8��0^�!Y>O��]ύ�᜾�$�Yp�z2'��X+y0��FG��So���$e���A�ϑ٦͎����PF�~慾Rq�話����	Y��I��t��rԨDz�!�3�Lӏ��:(u�?yt�=��)(�+�9J��Ζ-�8d�={��"k� o�'s�^&�5��HA$:�:���l@YU@���Ә�(`����XBV(ai~�ݒ��1G�~sO�+��M#� ��E;I.�Ek��l�Du ����A���2M[���ן~
.+�Ts�g�ϔ<Rvf�dSȾJ�� ����m�C�Z��P\lM$�9��J�ƹ{����m���2�Xό�0h�#	�O�/�]	����~�n,X�*�&獘����g�O��#5<�p��B5���Ec��4
�;�Y�}�8X��܉��.%N��	n�����V�i�W��u�樑l�'���=� <�a&��N��N&��!��4�!í\������i�S\U�[ɶ�d�H�{ ����=pWV���n0(AV���4��*eVG�Ƚ�'-��i��>&��c�>���#��,�X�Hs����䒳�UI*fw�����nu
�ǃ���,���BP�$�59�]�9l��T��� �����Ì�W������Z.��xl�_�M�U�n�
�����E1������q �v�	c$x�ZJu�Ϥ�{��bB���ꜰ��������]Q�^qW��l���/GgF���\���]���n�يWH��Agֽ�X��5��[�l?�O����s��h{Q�횵!�X�ߊ�S�%���/��������������5ŀ��=T�֏��C�Mi&�m '�ތ�b��q�m��z��uk:HE����>����R������|nL8� Ϫ��X\�Q���'Le�ם|��$����
�nU۠]���Y�t4�-o�Z���wL1(���.�W�a&�����ۯYR����S~��q�NQ"s���'�6�]b+t�c/���|3~�}�L}g�r �V�r�
�c��W����H?��i�Q
CJ�\����=���*�N�A���?�a͒����ь���æ)��C�~���iV!�! �J:*�;�g�nL��@�7�ͦ�\�{{BCe����u34m�*f����,�@;�bPC���ӑa�l��^������ga�7�R�\�v���	�u	��p���ѕ�WD��~���<kOF���#��$q�Q��3ĭ�-���>��7!�%���H�����L�ܢ�@�uַ�6��Bj�&]0{2���?*
о�J�/�ȓ4FgMLlSd��;�2CJi�) F�r6���_���8?�UO8z��b��;Jt�8�4����94�!�G�@[�\J\���ے#�9�ejs��)�J,�}�-M����W��`��,5�%hDSAun���� ��=1pm��ګ���|�J�>������E��ʭ�n=���y@���z�@܎�"����(���P`�e��O2�t=��T�f!��f���m�77��	MQ��.��6��翻��:�n( !&�΁ m3��g�R�@�!X�v]竦л��[���-��T�vO\`D��6z0�^���GO���HRF��n,CKFP����k%��D ���嵑Ax��S����;ߦ�u�[5�/��V���t��}�z
��-�b�3�c٢"qO^x��=���*�v:v(���7�iV��<���6d�>W���#���Ӹ��3ʮ'3�=8}��د]>>M��E��Y�{���m	49)]�H��%0m�Xfa�t�oK������~h���'N�]��S�L���C����ǛJw�ٶPJw�z�돽���<2��Y���ף�7f�b�TA�eqР6Ă~�]����]��E����E)b�\�-S'��O���[��O��%d��Q�Ԍ�ޞڠq��ܞ��[׾�M�|�*�	�7lIδo������e\�SQTt��^�,�Ykk������]�����~-�c�Vz�/pf��8} ]Y�_RaĪ�h"7���]�y��'�������I����C��7�����m��?�xUP�%�녋��LPK�A<v�M;������5u�̃uO�IA�Ȍ7��ms�'�8�3�h�K�5_�y���¸3*�K	:X�O�Z:�����c�Xx֌t��Z��oUs�~��lN���"�C��r$�J?���(L�.��酦����Qn=�̣
�TO��D���g�b�ܰ�K�ϯ����A�r� C��K��d�M�s����1�#}>R	ӣ��(h��b�qБ7�X��&��#G�'>4֊�A��0Y��nDy� ]6Oj�_9�1�54�g*�<�"��%C��d����t%�<(���QO ?���� �����4'�to�H
����#����=�a����I]M�ݷį{�����\EBM/�
��욝��ӫ��,����ǘ�<�L��� 1ȰY�F�<����U)��7d$�����!���vw�dX�m��x���=~�|>����Er�`����8��vqö��t-K�1����LW`��*���{�.\��F�&
�����GT�Y;����]�qt�!U?�µ���c�:��|(EC���mS�S�l�3����`��w�7�n�Ш�L~̥?�K3��4��
�������Xْs��JuG,��B�u�7�dm8$��@�W�g<6S4�_,���Z˵X�>�1z��Ɠ�����\X��l��[�7f�G�.�w�be����d���@9�mJ��!� �(8$����"[f[�ڟ��-��cѸN�d&��J鯪�8P�@�
�z�wtS����?�&��D`4HO%KJ�m�� X�I49e�>jL����ɀ�l�0���`��A��	9[H����K�F16Wj�!ؿV�$��ɏ?I�@�'pc�_�7`$A��q�m٘Æ,f��'�W"�ɥ��{gܒ�����g%.�Y�� z��gwN���@U�D�*\Ӄ*��3���<:FICE'~A���M����jI.�k-�7%����-6�r�J9֥�2���A@Ï?@��
 o�͠�:�]�Ɠ�����/���8�xo3�m��ӎ���EH���Ad5�am�JW���B��@8�h.�3&���G���"I����GA srx|�F���ʫ8:�Q=1|�q�sH��"B����#�O����=xL�.�t�O��E<�}$��,��T�	��aN:p���ŀ��m�a�#ɸg�7Ԧhk%�~rm4}X�tl�f�&#�v��s��/2+��B��ТL�9����T�A#�x2�$2o#b�sx�R�>)j2���x%h~}����Y�7���l�N9�|9չ�a/��'Z!#��5
B�gE#����N��D�*�kJ��������_�If�J8��0��)ʺ&�D��V�qO��l>M��7	[@>�9v�\
qF���|e�	0�E:-�(.?a�tA����³N�i�b`���E-C�ND�fg�������ȭgD��2'���)�)cH���&�*Mq\ˏ�\b2�G���	�9hjdx!u�2 )�e�ƽ�.S�j�h��m�	(���\B�lZ��w�9@��H��:	^��yAtPDǟ m�3�X�Q���Tz�v �L����>rObgn��I��s]�7�P!S/���,I���R��Y�t!��
Ż� ��	˃W`��* 5���%���A5Q���q�/n� DCӒ.����k��UފAg7�ao@Y1R.d����Ox�l����m
�@J߽��������=�q$�p��_64�e8��5���Vu��Ni;���-@˄��0Hl�f��^��F�N��g�\8Z��ۋ�\<�'�,�K兽w*�_%,�� ]	jαK���,�Oͣ��
L�>�`�c#Ɲ�lky|�K��s~�JL�������C���6[�����'A���Q�X]�{_�E�`����\�56��1s�K����������m��;b�=Fw�X��k��xp�<���o��1D-��$$��k���7�II@�`xN�9��U�8�*yY�����5jي*�L���Z����xe'��4�^w��V�yH:�!4�.v�]�e��\��a�_�kBg��[�c*U�L5�Z�߂R����VEө�V��{�D	_.υ�6��F�X�3�XI"f�W���]�;��\d�����5(MkC�o���=����w��������� #�3&�]u��Sb�£�8���c�9�'��M���^�9�C6 Y��6M�b���w�Ӆ��(�����C���9�T���dx�j��u@��֘�gzS\�����O�ݐ���K!=l�%k��zݟ���qhO-�k�)KM!ue�f��^@�[bȘ����4���b�8�[�� ��y��(��T���,B7d�ȃ-�?�������rh�1 ;������)s֜���%	��VO$�wN���w���݅��4������(��.!z�VH���t&�ÃZ/mHUoL�-�N�"��B�c�9�a$Ѐ4�+��#d��m���Fm�G�>�A�HUw*\ ����[�,���(�_�ez�VUE;�wx��� �2zC1~D�k5����N���5����@����7Wm��X^�g."N��Cx���$�<Q5�vq���悦�����E����+�ӯY���]"�}!�V�/�Q��ֿ��q���}.���ګZHoY�`�j��&�<��x�@U6�c巏X2�-�D�4�g�T�}E�$|�ݛQ\!1��'�I�G�����/�Y�#�o��j�w�ꁞw5;��k���$U-�C����vT��WMF^�z��5������K �6r�$D���f�1��;8��v��+a��-��bQ"z��'k2lH����͙� U(��Ou��S�?���S����|)��ξ���+��x��p���'E���uȼ�7����s�f���z�m7cN�K������R�tڝ*ұ����9�}q�gv"��E鷴˴X
��
%���}�\Ү&|�j'�G�{N���1g`k `s	�MūYw[�/��I�܎��>��i�VO� �0�����i�,|��1���=m�w�$��M��x�dl`3��h|q�6+P�R������n�h����Č���"^�uH7�胑�����@���\�>�'�A�2�ׄ��&���7�X�`~���b�N~顑�eC�*�����2��\NX� sZ�s<���EZ%YlL	��r�d��C-�T�?,�%^�Y�7Ԍ�8�Rd�m���}�gl(��qh+�@>~�O� ���ߖ�`G��t�9����.�q(JY��Z�$�D�O1`�)�z��$�R
c�,u���v��S4����7[Ϟ<��t����yŖ˛)=�0h��1~�%�K�qk��3^�� �u@HN��g��aO,	#j���pE?��qi��k����A�e�҃�wK�Cz;��h����ִ{�j�-���k��u�gKFD���b���u��QUi*	fWJ�� ���,(]�s�J*����M����۾�������)����ע�D~�ܒ�wh	�y/�����/�ϯ�r&&!��(��d��%*�eCT�i�.6S�DVz��ߍQb�L,kiy?��|�[20�)2:��U�:�$��pE�"0� +���m�M���#bI?��ҚWu���a(/t(\�r�偲X��b����5m���)�:ڷ�G
m�����&���6�F�;AB
:Lj�����-���Q�r*�40e�m��A��о��T�9���٠�Bke�?WND���� m�[�W�U�3T.��UK��=���w��΂�N�Q�IVtx#��k�F��
|�ɗ���Ɲ�`�T�������.�����q��bk�b��Y�Yd.�������"��K�����  Ep2'��8�g.JG�Mt����UԒn3�`z��a�e���+W��6ƭ?
���� �v-���	9%�"m�I%/D���E��HqTH!O�d�/_Y�dv�� �DoJl��+t�jʀ�2��ᚵ�GM'���3��[�(:�~i�Ĺ���qqT��5�2�x��1�װ�>�u����h�X�6Zn�j�� ƉPl�ʾ����(��K@�'Ջ�����*�(q��po$��S줝}ĳ̭*��<$�b��)���=~��Ϸ�'��A��5�}�Ix�.
��_M�|%�͋C�D�/i��U���~6l,��?���YfS.k\&A&��"�uz^�q-54��������+J�ٖ�p����ȿ���-e>o����u�1��j��Z;��Yv��� /���͗�,�JN��(/�Y"�#xy�(���;\��<-�$��s��Q���q�az`~�Ot�ڦ���U�U�mC�)�u��y���4��T����qM�EɢIa�cW�*g���If�TF�hgR���me�;�CT
%Ԅ���ȳ�4�G8�q�Bځ��JC����y�~�0H�Zݵ�0 4T(~��?�?\}��&�ݫ$����=�Pk�*��,�)p[����p=��n�dWK��b\�i��#c<̳ܢ6�9�|��\���|3�1�[1�U�Jr��o���5d��jжM�U�8��������*�]o�_^����3�=�%ٖoS����w>j�Kr�Z6���LFx�4vӤ�8x�28ҁ;�E_s�2�I��c^R顿%"��2�������Tr�(���rEc���S[k�ki�Z�3��@��V��Bj�s�!d�î�"j��Py��� �\��Ǡ�2؊���e��K@%F�t���FӻY��8>-�S�R�N��+�6�m�S����3w���� FU��r�6ZIS �:��C	�w�;�9�"�b�5������FJ�A�&����}�[Cޮ�[�ۼ����1ſ���j�Aa<���\r/�����!91{l�9��ܙ�S���z����2�U]jW��� ��Qv�O�X�
~=u�F@�r���#fz,���.e�Ά��;��*��}d�R�L4h�`�WԲ���z���,�O�[$����uz%��W��G��h��<f�5PEy��&@^����V3���5,2L(q d�PF �H#�C�4��}j�zD�sB�s9KM1���C4��Xn��Q[Y����cޡ)ޅ-ǊU��K���o�fP<On�RN��ы���l)�#<)�9��1��������ͽ"���+�e.Nэ�n$h�xN��a��1p��B��!dX�޻��&����+˺�T�f�w95��g"�4���Ƕ~�u����nRl��zt��ڹmi�"1�Mҟ��*�6S��ZEhI)K�lE!�>��N�+�EY����L�g��V��`�7H%W�g�[��v�l�{��V �e[*�	p�]����rX�8ţ���٣��B�=�m��wˇU'�$�q��݋}I$��8��t������&�V�,]8��uiX�d L�Y}�w�h�k�������:�e9�����}����:��u�f>T�!�>1��Y��cS�1���[Q^���a&�F�F��F������	����Cџ"�I�m��w3�lEs#1�-Zt�Bu޳��89� #	9� �ćB��l����1s�%�Ռ�
H��1}E#�6��)��y������������VA	!����C�k}�߶G�(��\Y�u������wB����Д��ؤ��H�S �����1J�ڐ�,�� <����\�R�R��bać	?�[o��c�LQw����܂W�ڠx�(���c�q��0w��f��M��5�Py_c�<U�p����|9�$��C���N��A*#9vW�>n�ߓ�EQ[�`~v;#��=�(���&4�/%s:�_�X�����0^�D���X���G�(Z�+�O�I%\O,z�A�!wJ*�#'d���@���;q0'�-����,A�7i�.yU�NUf�'p{��͟��q�����d�WkfZ���D"5�3�J���U"v��?�]í}����ȓ��h,�%z�Wa��Q~7�ӗM�,PM�pWf�=Tǃ@8�A�Qi/�
݆^�H�R&�v�Z5��~:�h���B�b뛼W���N|���[<+7#z���QGx�[>�,сa��-(�:s|0
�ց@?�HG�i��
������&8����q-��~�+@d�_*eg�wFZ{3��Sq�,�\!'D^	%���oL%+ϴ6L�C�J&��<�E�/F�r񀥯�Nu��e��q��d�s!��cT��������<�?[^X�5#T�"p(���zC�	�I!^�·=��~�3�Ɇ�h�F��e����R��~lW�wRQ��U�V�b����"��E�Z5*��n��n�~�5�4#3��к2ٖ�Ӥg�Z�<g�f���TL���Ǔ	@ C֫�X�K���)��Ko��0�7���A�kY�C��Ő�&�c�_DX.�j�=���k��z��z����e�p�'�*�	���Gi�˭���5H�̣,�n���)����& !��|m54��9G�sqB�w�P�5�Ի<Z���)��IRق�}\��5�\8�WKU[G���|��w���H�@p~�9�� 7�ymFF]�VC{�FZ��c�:���c��R����hd����U�lr�Ui�-poB�G�Փb��/sA��I����U@�o�*�N> �!+��|�(RĘ�!��S̖���{����'�M�̬���&�f�S�<��*k`�;�d^�ew�,[������-�J��?\sH�P�>����Ӽ.NS`NYڗ��h��i��q�n{�3���J���[��x�a'6�2�5��m����r�ą�婫�R��2Z�`�#m~�h�[6H�����|C�wD }P�f(@x)��M ~��U��@Mչл�6˧]��MGEcǅЊ3oiL�v�{�t|��«��� )����4��ظ0|CK��j� ��i��MO@O��"�y>��TK�A����J���;8��U�a1̦���[g��j�9EY��a�p�W�o�d�N�"�2���xO��Zu	Lb4Oy�a�F߮��P�9&9a��$��W�+�9��=n�m�R$�H���u;+���X9Sx��@~U�OϢ����:(}|�+u!O�(��Q3P]��<��0�&��j�rd�B��G�2N�nk��a���a.�? yR���3��FIP��D-`� ��&��[l����9�P��:�H{���=�"J;�ٶ��j��%V���M�Nc��; ��6U�@κ.qc�����
�b1U(�d��^ţ�?��:�#�� ��*��-p�*hJj7ҳ�?��cIT�&�'�WN����X��	��5����xb� �(P�=�81]�d䡛95���o����J�����5+"��ڏ�5{�%��ZM�ԲbY����J;)��xh�[�����G��r��U�&o�=���G�e�Nڼ裋t0s""HٹE�x���N�q����ԭese����K�9���g��X�Ftp�P�#j'�j���e�����*��o��0���Qj����"��oYb�5h�f)��H��`sjc����9���&X�ͥg�%�Ǒ��H�n��)��bP*�ܾ��M�n�n������Q/SLoT ��%��9�Wa�4���s�;K����EL�0i��'����A�*
Gi��z�����*��Y�H�8�X���ܽ.����a� ؔW'�	�B@��P�"�i����#4�1nS�����J���N ��S;՞�E�t�Lx}��S��nF�2�K��Vl�,+��D�}$�,��i���FD�[�a+1��(LS�+$��O�X�����k:�q���!����e}YҵpN4�k5gC�#��8Jӓ\����MO�힣-�I-�bE�z�����X~�r������ؐ����n�L�䠡̮�u���Xd�g���iˣGZ�jc�HCd�0X�=҅�qi�����heʞ;�l��R �,�����!��r��K5�IG��m~��n7jJ��h�Y�n���ӆ$t����[:�͓��VG�[��x@{i��Uc�h��u������F�̐s)ʞ� �fK��o�ӝ��;p9�癀3-���|����x�����&DP�� A�p�Ǚ�2L��C-h���"���(��k�8d⻎b'r�X�7�V�nZ�h�g_���.��un�y| ���`��1���-7��$6���U2|FN�\7��a���8�:��K�7�����5/�F���h-�ZI�`�������1�����3��τ��U�9��6g���h?�Y�4��Ɠ �n��Y��c�9Z��Bկ�a�ʧ�0(�?۬�=ƪ􀇁��>�	
	22n���:��FU=H��>��?�D?#0�oV��q�3ډџd������ߋ�դ�j��t����i�x�c����6���Ax^���᜷�&����Jپ��˗�F���-좃!�;�F�;�6�WQ�1n�$���a�os�㓺������ 1��xI����w�zT�����y�L��m�I	��&��5\/��~�_<�����aO�������
�R&�5���X�p)�3_l�O�+��Q�O��h�y4�@^]P��Q���%���<;h�g=�I��ɻ'�n�\#75��~2V��jč{��$(����'���їZ+#��zi�(Q5 �z V+����	8w�7�L�{�8���Lr�˪P�ʁYp"�k~��Q>���F�iW���,n�'��B�c�D�j+F�kOH}�����E���-ڈ���Ӯ^�Mf������?F+�
�ߐ�E�a�Fæ�|�rTgzu�h�e��9n�?܆$V�2�z�ӷ��˗��7gg�B��/�����D1ʀ��uJ�ۉ	�w8��&mPN�o�9z�m�9c���,���2���	��|iaf��O�N�G��\�K0����(K�����,�9N\$؇�.`F�]��V7=���ph�8r�	��f��95޿���W[^sT&I�$Gu�l�/G�n��i"Pu^!�u�09��6�cN��Z*����K4�I��Ė
)?�|­ɵb��OW����V����f\bd.��wc����-!0c�w� i#1��o�b�]�*Sʮ��>	a8JH�y.}Y# �M#leu_��í��}��˅��l���4�̵g�v��궑t��j����Q�ଃ�>�XH~�m��f���CZ&{xu���03]�9�3ʠ6w�{"\�S�QKy_���2��ᓠ�l����:dv"8���Ց�8��F ����Ҹ(�j��2ҽ��ݒ~�ֶO�0�c*^[����Y���$w7�� �ٲ�
z�����Ʀ���c���>�g�)��>�&�t����ⶂ���kK�3�9۵��C�bju��Y��&����{4ʽl������S�8ӭ0�6�
Y�������Ԣ�<t�V�5�k��K�8%���w؟&.W��~/�x�7��EGx�������9�Ilٌ[�$@��rۏ��������|��|ةO4Np���2�-�Io��6F�����f��q'M)�AL/s��aq������S/s}mr F�~����g�=!������X����8dX�6�W$�]��`�7�?y��s1�`�O���A��7��s��X*ݗ󏟿a-.N_�ɤE�|o�x���Q'	�Ʉ � F�bi94��|��+-o}V7�wq�)?[�_P;
|m��t?�E~�D�sg֙��A���'��ɫ��EOl�5Q���W��q ���ȞI�\c��b]�>>�W�UAy�.��y��3%0�C�x�HG�oZ���f6\|6D<�:���4��Bg�i]���Mˈ�}��ˑQ�|�ڶ<n���n��6!��_i-�<x�;�Sx+��:�o�;�err�:��7�Ѭ�'9�0�0fT����}#�\.�4��'@5['Y������s�r���Vk���}��qA�@L� "u��C��8�3Y��GV�8y��
�1�z�lg����!���I���,1k ?�;��m$�&�'�ԯ�����a��4���C�7l|atA���|o���F;�4����ɻ��4���C��T�u�l�{)V�"s_e�GL1�Y�8z4���5���o��7JkJ��wHt�����*�0?��`IXl�HJV��5c@P�f����(����P���`v	�N}<��Nƹ,5˛���ݦ��OX���5�w��&G�H74D-rv�A^��{��R�hѣ�F�f��p�v�;95I�= ����c�I�ui�&�]�^I���ڷ2���,·��'��rc���B'3�E����O��E,)��f��4�(��8D0� ��&��������5�"��ެ&@�r�eU�ݟ�����QR.�{Q'�^Q$}��N�m�$ ����Č�&�/:�pUU6�V���h�3�>�CaI�������5��\�hC��gmK;{X�w�:'j��܇=���`������圁�U�B�
����\U^\;8�Ŧ��+�����m
H8`	�m�/���"������k2�Oi=��	��X�뛸��E�h4i9p%����0!qN`z�GF��~i��
�,~�a�{�����x��l�[��uM1M���/�7)&Jg����B؀�f��i����P*� C/::���<�<p��%+�Ş�8��%�^$놦*��j`@�EQ.,t�S��oGh�ؽҌ��b��aܴ�F� 9I�:�&���lU���^A�K��l�?�|9�ܚ�e�g�����( ѓE��V�ᗅ��޷�i6t�����c���<m�1�Z�a#u�*FѴ6�ҫ��a� �?�J�&V�Dr9T�_��8���Ȟ2T�w��o�e~��>b &��6�8���Zi�k��5�ۥFgR���x�C�`��+\��X��+0E�y+,���6���\��j<'���i;֕�!�glQ���[0�����$\X��ZX�i�:�8�A1R���l���'IKk���ͺ3��v�Pv�?��qAB���Q~`���m�rԷnn���p�h���us��)�^���M��lh�G�.�	W�$�>�N����M�Td�K��5��Su�.�=cO�j��$�v1����{�Y��Y�3Q���q}�F8�sx�:7Qj����	;I�YH�C��[�G�7�݊�%��Z̗���{���?�$��f��ȸ��Ro�#
1���;*u=؅=Zӽ.�<xz���(�13L�̂$��Q*�L1�-���n�\�2b����L��n4��ɱ
)�W��SX��4��>c��uv���޻�`���!s[��)_wQ~�������B�T��/��v��c��'F�<tC��>t��!�����X�� B~7Ұ����H`zj7�(g�Ӭ�9R�qUR^g$��5b^u��L>��Y��V��¬lݢ��I���B1�׺�,k7^2�l�M��a�h �({.<�2�%*�[��\,����pn��_֕�r0�6���&es������-x��댣|oςm@�R�����#���&����R���g��`�g����twf��ǉ H��)��F��1��R�S�gјW#C_�}�v�T%��M+^��b�%i	o�#����r/'H���@��$��^�j�;z+B�����pi��-�����:�����!�D���,(Mvbz��}��ɑ�v��g�6���/XY���?�
�Oc���� �Q5L��Ep&�fNޖ�? ��'9>��h<K�F�M�=71%�9NE�yM��i5`e��Ec}���V~|�זּ-O$!Ĥ�v0�'~T�O~r�q��;G�1��������~v�ӊ��X����K�n�\�SP3�!έ���8��@TK���>MK�Q���5���V}�#��#N�8��oĝ�٬�S=�S v��"@ɰL nb��5�6W��e���|O���Y8��Rlo
����UеIe����4�s���~п�VF*P��6��3Z�?=�d�V $�(�v��n�sc���[ӏa^ZV�7̟3�wF��-4����W�݉Dv#%��'�C�A�$9�H=�#���s;����q��Ы�Y4,�x��;4�}��b5�v�״���K�97����N��/�{���ܲ�y�g��)t�b�εW�a�� �3�6�k����2�;/��5���^���>�T��~|��:���jJ��Ԥh�.�L`�%���Q��)�kQ�Ŭ�׍���~#w�wd�A_{��,���v��`��x�=�:K@��r���)�N��Ig�
�z�uX�-���>Cմ͚�؁f�ԘD���|���1��݂ۮΰ���w	��d�8H`�Zڢƀ��/Ǐ��'��!��'s��ErHvr� �c�l`�&`�86l32��;9's��o�2\���L��L�z�Q, E��hhA�zԹ	J�3o9gd_V�i"VSzy���C��*�^�@�2����o�^≮0T�f��?�
z֘�Gkn?X���. K֖kķ$\�e�s�P$�����w!��X�Xm��O�v��'b�r�57V�U ��36"y��7R.9�u1����*��kpj�%�e0D��l�'[�,��Q�Qn�Y��d�O���ٷ�:ll�!I�[K c� F�m!�Tx�6����(�U���'�%�ǌ���G�mF�����,\̖�T�x�ُ��Yq30���X,�t46�8�O ���{d^D*�=���E"���8�{֟�y��]�h�F�F	��� �67��H��[���c�>Bk�\�ȧ�4e9�InHCj�HƷ�QCh��!�~�>��[m���! K�����e��A����bE#5�%�+�<)f�V�q�$��1�5��K��*�,xt��geW���ʢ�WE�4a�	ڜ��##
G��lmU�~(�'�c?>�6B_�ݸ$y9���9�c���x�ӑ6�0v���eo�����w�7�ILyw�C��&�'6<-���;X�1q��Rb����&�Q�< � �ΕzG���3Z�,88WK�����c��U�%(�H�/ӟ��͢r���������(���A�������֫z���G�K�[^�|P��$�~��T�6�{)�e����^�ބw�L�%_0Ջ	}2d�Z륎����{T_��u�57<���"h��K��ec	;-���@#����?�9~���K}�}YvU4J���h� ��Z��p��8�!2u��.����C��:m�Jⲿbc6��s� #"��k=���IP Q��>qN��-4�<�K��8��e��{.9�狘o��x�=>K�@p�j�umYIO~�>fIʎ�g������)�������VؘGF�$;�*L�ڦ\m3�JF#h���T��F�pTz��$�z�߁�I��ë�*:O����CO�Sc��-�{��?���e�a<I�׸Z��O�uΜ	.�C��B��i�
õ؈5�&F`V�څ�����sE����,s���Ѭ��}&O�\i|v�<�7���oka�H����7��Y�6�G����N�-Y�h��Z���b^�����I��pW�т��z�%#�ZN����諶Q �y%Zy�%����e;�x���!���fk�F���\~��/�9��YhK׸��䒟e>�o��|V5���<�����)�"�+�Ac�1����Y5L�^|Oz��J�o�r��J4�9���g��S |ޓ)=,��q��QGZD�Gxd����^�d��A�?��C�#`>��g}�ٿ�8*�[r5p&M!���4S����8��Q�"d7��;�����Lrw��_ԑ�wCvu��_��_��6'���Oa�T:��S��pg��*G���3�H������zW4��ao�˼
LK�h��"m�t��q�C3.S�}:�L4��D�㣘Y�`�Q>3�11��jh�d ��A�a��C��R��̦���o�Q2�S��qINaM>!���Q�R(T����*�G��'�D���4�^,l�iL7O�"��1��Pq��z�b݁5��6j��!i�D1g�rs�������F��dq亾.74�d��G����D�L2VvvO
Kr�q�P��P���&2D�ĵ1s�Yk��J��#�y��8ۆ{��p�.����م�Ơ0|E�aQ��e�:W�:koU_A#ҊO���cu2w��Sz?��_c���F�W�a�FZ�WGh{Aw��i7E�~��3�L�����M�h���]fI=�a����Y_�I{�jͯ4_��~6���cu�>��`�����$������a)Hx-�g��E���%�������C��M+u�*����H5i�^3���򎆵�vƇ�@V��*��Ӡ�t���� �.4JP�J�4�����8
ɗ���s��������3�?�u8/�0��S����0P`#��P�n�ϙǠ�HM"A�"��x�f�<�Ϛ��Ҡgk敪y��L�	����	�s��a�YA�+�������4.��q��_�j~��ݾ���p%�d��Hu�ש��\���K�"H��-6���Ե��GJ�k�oç���R��i�mIC;BЇxu{�x��o���?k���XJx����y������TV;���|�ZV�l��Or������u%�nzw6�ˬ
jQ�uY���ް�b���~��`m[{���gˉR �f�2� �9��J���#P�����ϣ�yW�p������ߵijPy�PS�U��^q#k�� S%"�O���C ��!�ç\5�����&SH��t~'���CBo8F}���[��cp���l��L�����NMJ�#X���{�U!�]j��P�m"���ђUYa�#\Q�s�gr��2��]mY�x�	"	:]e�� ��Qr���s���omͯV�scv13r�4��s�YgLo>b�,�`xB+�A�)���gx���´�0��~��^����\�?i��ݖ`�W�V,�_�(�����'͚	�]!> }�h-�б����5;A#�#��0����#����E�v�4��Z��@��W�e�t�m��Yc�,!�Z�V�7�L���ٚ` ��w,<�V�q0D46}@���"�J�R�����b��G�s3��Ul�~�-V��'QtX����g]�,r?4��艅�?o��r顰�%c����B��z�㥾��QA�Xȓ�������B���'�ю��ے�/Rץ����)7P7,����7Ԉϲ��no���=��G3�F�����m�<5�<��sD }��h�8����%����k��3�D��s���[�5�u�����ː�kB�st�P�}��V �_��%˔ӆ+���0�꟠��[zX�b�:�Q�x�ș[�����r�s(��v�V�4���]|:�~e"YʜǶN1��}��I�̾�'Fmuo_��i;QË�.���������ż%������dd�8q�g'��8��W��u�R;i�Uf�f�L⊘˧\��I�.�[�ߥ�sN����;�Gʉ%���U�0�x8�-�Z`�3�e�� @�Ͽ�C0tu`��}��n�	MM���(�W�i�p�Y#u�C�����^YY3�:֧��"�����)��$>]n(o^�˳ ���y���ej|��<'�\&��n�R8b�J���g�b�puՏn6�d��׽0lL��F�~�-(�0�/[k:_�K�jh1�p+В��g)H�p*^��������N�2�VA���M'9�!���>���ȁ���]W�т�1�ޣ{FӖ0<���=,�t ~�E|CJ�m��R}�Y�A�"���K�m�MN�-B�݀s�Kӫ�)��[�(ޤ eN9oo���Ê�V�Q�ţN�G�w�d(�Z�l��z�	�㴧ExCvHrw�8�,������i2tң4q��<�@�"?mL��@L2��I��(�K��w>r8�tY���x`)2I���*4��H"�I�U���e���D18��.JN��1�PQ_���ƌ�N�0�%|�Q���v��$�'ܜ������J��-�g��w�C��E��;�()����&�Dʕ�Ϲ�)^��y���q�17�	&Yl����Ûw���0��/**w;�.��8�I,_��7��hR�ƶ�w�av��6#(�[�B��ҁo�'��Nv޾�U�z]�|L�A�gi��"��I�%�f^�.�ͩ�{�hڷ&Y�x���U�灹Yy[m��Z��D���Z3���mX>�S9zB�AHNm�S�Rv��D���IB̞�]�d&d�>��L�'��㢦�I������gbS1�,7)�m�m�P�[q���C�UK��$�l��4ukӡe����I\e��=�-x	I�<z S��������`���W#�Q!���gcp��� �G�T�n(;�b�?����3�R^�n�TmI�k�:�&Y�ΐ����x@KK�B�[�;s���e���\E���� �R��d&��^n]Q7��ch�X)���Hc������V���>�`<G���9���'�����6�������SŢ��d����n����W���������>�O�������ߚ.����+�M8�_�0���d䒘���ߠ�ud廉��S��'�`�S�u����I
g�G4��K���8pZ�1���-pD��g�h��Cd要?�Z
�j����4�����	�����E���4Q�,���Ⱥb���N�dZ���5�O��p�����U��*���O�ڑ��Q��ױ�'3<��q��[i�߹��[����v�Q����Zh�~� -�soy��H�ݴ�m�(B-u��,Ճ4��.$� ,�l������ָ��O9�)5��O��#�Dr+�;!��r)�FRy(��p�NO�1!��us�i2ea�|�Q �+�U���\���&����g��Z��q'�F�D�G����a��g���|Ҋ&�=�Aܨ�("�v^���u�aR�,\/������.�;�A6��l���J����M��cԵ;/�-���a��������)�Ь���F�	b���"��2��%�����*��G����׆���'^+�o�[��ĕNLw�ؽ����H�������!�VK���f�X.�������'YϾ� ��`�ו����IC���(�:��E}E�-�ָ�@0�r�� H���!2�E��,�1�b���n�nY��o��djD��&^��c�>Nv��m��<R����X,,<N`�i7�wf�
O½��y�=٣�{[-��u�nk� �%���MN���k�ɿ!DA�o����I�ؕI��*�]"G�px�I����x��J�oe�����{e��p�gƤ���""��<)�0�b���!�E�m>��_�����8���:t���-=�a�J�Od�gu��]����V�JkJ�e�U���ȁƞ��0�[��+�տܢ��m�X�M�Z�������J%�4�#�rd��6'Ϣh��Ɋ�{"�z������ֳ�E��s�N�/����3˚��<p�A�q���Ş*�_[hI�<
Z��:-wJ��ħ�kڒ��x�S�5+K��I���E�fi� ?��>{���%���ϓ�O�'�h�����pk��!��vN�G���t�ɞR��_ey�4���ҪP��P95UK�_�O�\f1��_�.�ތ���1�Р<�O7;l��^�?Xɏ3P��d'�������>��6~S>���CU��b���Rɘ�/�k3/}�� ��y����Wye�BD�=Q	$°����c�G��y�|�R{�,�#]
���a�	��wKA�Pn�6*���ۑ��z�a�h?�>��ܑ
`���ę<֫��Ҩ���S~��`qHуj���צ2�d4�|�+�������R�ᱴ	>xE�B��{�$F�7�A�<��q^�����_%�{�	��=	�v��j�l��_��)�\��hҵ1
t�3�),b�k[���ι7�S�e�(��8����W��d�~�V�����J��=��A�c�6Wi3vT���|���5P ��N��|�$"d~f�a�.�`6#� �.X$'E��ҭ�|c��P�X�TҽȠ��7Z>���$Qh����('h�E���V����3 o<�̰o�!��f�ZAj.�j9�[E�i�ݷ���Ʊ>ьG� �y��^�l�8�'��2��i�P�M�Z�C[���X�nA|��f K-���:�S�q��KE?���c�m���g	�N��8Z$j4�Z)����p>��O�au�7�/0��d�^e��E�;�8|,��B���a9㞍��N�dW{N�q� g��c�rH���x&�7�76��I�r')n��Pك2.$Go8:��A4ϠYx���b���m�@���-�d�Pkީ-�Z8mZ$��=�}�d��W�1_�qh��S���V~ ���d�Χ����LmpF�\=ri᱋��ÚO=���&�5&I�j���p�F�R���~�?���*��������{�<�q"E/�n����ϩ� ���Y�1����JU�N˱�r�+?䰲�_�1��^!��ޚW��P���S>�*��(@ƴ��G&ɮ�lJb���h9�5Hnq�(�U��:C�w�=+��[ɋb�-����E�Xt��M3�� Y`g�C�Fr�)J�<����rV�!����-��|��ePy��D��zI��{B����!AB���kT�%�l9g@��A�H�S�yI��Ϋ"	Qe�>9J|��q9L�|M�Ar)�� Pݶ/�<aB-�4�!}X�cƫG
���s7���"h�좺�{��l#rۄ�,ᛧT2�9�d#7*�2��#��tzg0�}?Q�N������V�DʃwV�Α�����F��T�"%#����iLI�����F����L�nȚ�7��n��[������&/�)���!�I�~ݘ��ga��r�Q8��ր�=e��_QD�41x�d̛K4��Py��*p�k\Ɓ-����ЬE�����,|���`R����xZ*��R�d3��?#���Y��ʘ
��pG�	��I�IGt��+�br8;;��J� }�3T���c��-���K���&
X0��1+��͟Y9$����t"�@�*k�h�nA'�Pf�g����ላ�BC�-�34��}[yU*?�0f�P�ab���A>���'�������?�U��76�Ku*��ƪ���*�G�$h��B^=��,���������!�p\]�9�B �����>Zl�8���Mi/������o�+OZ�UG�Ne!,�����ԝ�X5`A�D�9����<���r0��>�!�:�eIp$�r����� �ۤW�
��ۄ�X�8|����q!�T�p+��i�r�dK��4A����a��D�c�t�%u0	�B
�Zq��Q���K�Z�mLEy��9?���&���t�����M,����1��o�N]���{���W��=��s������z�Q��b���[N$�� �a��`쐍�2y1r����!���LgZ�,f�/��>���4���>�ES:2�*M�$b�e��Cwm]9h[y���aHN��Ș��	e�����Vc��̊����p���F!ͽZOY9/ұ���O���6�4�.Ok��Q ��IC����!�p��#۞'��aF{xZTk3�\�K&��3-�aD�+JK����z��%�����X�ԛ�ϯx#��U��9�w��AR��U	�2h�F<*ׇC�!!����B<+'��Էh9mhT�\�)9�]H��6�f����3��fh�?�)X`�mN�����@��[���L�&��!.��w$���YZ�����!T���t�{��BB����.Y�63as� �}"NLrsN��K�%~f����[�lHMg;}��GT��"��^�N!� ��Ҿ����b����H:/��cP��-�3�Cq^#���[��Т�� v?ѽ��M�U$#�����MO�V�V)-�ؤ��)K����z"
@UF��b�v
��Z�uԴ��"&Z%�='>�m��V `�����.�z���H��8r�7��)nf��,�/>����L��{q�fQC�GU��TV�d���KvJ��ո?�i �7��/d�n�L�2�|v ægһ@(�,�3<1��L"�Y;Y��ɿ/M86�x������F��vǏ��_<�.�O?��=2
�/�źG3a��hEaC�`��C0�g�ݦk����ô�&k6V��CSp9�%�m�KD	���)�EL���b�]�o>N���c�'��[(P����M@2}Flރ��.����,)�i^f���<�/d�E�#�]��s��-.���[��@%�2E�+���3�ᐈ-Y��O��r=���"~��V���m=�� �%��fZc$��lI��%~|c��%�e�P�6�Ew+Dj�������U�C���J��:�)]�ل�Fy����Џ��%7L��R1.�mGzdX�d\��YrA~�eŅ��9G�U�I�/[Ӯ�=�����0<���ZX�PzƮ03hrT�n�2�*ιf�FL��PGi�2.R8�efV�`P�x�cY�0�4AG�
�uںw�d�A�N��n ���{��K功#��%5�����ʉ�����jв�ssϥ�J����}3gտޒ���1��C2�U���X� i�'��wr��}&��(�6��$o4v�]�L�;S/�oj��X��M��'����U��ѪG��ïmz�C!���S8s��Vk/#����7R���4��f=k����⚐��X����D����q���_���kdk�ݖ�t���ވw���� ��,&z����͏ӧ�Ֆ@����Po��S�t��11\$p-l |Av�5!c�;c})�ȧB;��ìѸ�%ǩ�� �r0-.n�s�:���5�[|��X>0�\ؽ��yx\/QkO9(V�B�!�a�Y�� <"�[o�jf�\!�b����ެ���N���}i�bh�^��1ٞM�5*=�ey�3 dggT��$�u������ת�$͜�<J�y�Ѕ�l�@�C�A�����r�>��x�8>x��@B����`:��A@^4�Vgk6u���Z��a�+����K�UK*��[��1�v�9�HA���!�~��fK����4��mb
��}�n
���>c;�:܅}��t�0�U{*(T1��#[�ͨ(p�h��D^��vN���Ҕ��W���x0)��X9K�ܥ�K�Hܯ��t�_Z��#�>9- T���|�yEg)�K1��Ч�z91�]a5���*ۘc#%0a��*�3������g�BA,�ڽ"�H�]-+%�g�[߸��5��_�����	|k.Af���8!U�˲���<xt7�f����̥�����&c��K���Q5�z� bH��+^�FI���RS�`]	N O�0 �i�E����������y��^�U4�4��#,UFmT���R���!�Yp�QQ��r�0)�'�me�����k�������I��0���Ju�����7g����'G��e� A�E-�çʸ�v:R ��\��G�-_>�����4�f`�4k2�	�wj�5�C��-5b��ΧE<��a�X����i{��ca�93~���bF�mzQg�
{���U��*uL9�u��}��[�'Џ5�nBA�񹒮�L�I"Qo�!`�C����E0����F�Ҙ�V��7B84��h��C�v���������=�����Co��
<��O}>������hnYo��7_k%�ʟW�Ɍ��9�	��*��JVܯ�]ڠ!�pZ� բ��)� �:���%���b�V�}gD+� �AL�S�7�+�l(;� uu8�7RHq~��YrP"B�?������D�����Sj�ty*R��Eu?�8l�&v3Xh��6	�[;�\��~��� ]�K�?4Ԗ�!�o�_�Tm����}����3�)�6߾��W�3�Bʮ����dx@_a��g:�~hy��Z���ӾU4��$af䙉q���s����T�g�[֢zub��6g.�UP��y���eh�-��&�#�
a�Nƪ��BHZw����k�V����I�v�����n}��ʡ�7R�|��TZSq���c2m�kN`匬�ޛ���Ƕ+9�v[����P�Е�C]4R��qR :�)�!�Y3�Qw��`\@��Jo�v����r)����Gs�ڏ�gA���	�����sn�>#���ŹJβWC�B�YU�pp��H���;^������P�$̸r1���C�}�@5��d����T�FU!����TrBX�Ө���/���\Lآ���ҷ/T���w�b_U���4 ���B�/}���W��V ��{K�ޗ2D#�'��<�l��3�_г׬E{5��Ĝn���!S�i]�M�L4�B��W���˳�K�8����(��v����5^vW�
��$e�3ZbQ�|y�N��r�<�*]R;Q�!ͣ�U>�`[X����y|M�����轚EE0l�uu��pn�Y|ܬI�!��ʾn�Ey�"*�!�Ph7�Ȣi������QY�] ;��	�PDWN��,~���j�el�9�����Q$����(�sp]�.��v���0�_ ����_A�hR]�ɮ#.D(����>��@h�qt�bE4ٰl$��<��r�}a�~�ſ}GʎŰE���W�,m�LT����G`-�8���,NM������6j�r��W'�D&���G�!��MIR�4m f����u5��U\U��/3g����f�<��;�yi}�xC2�3�i��Lt��+�D�Ǚ*�ۚMʤ�(�4	��)O�5��[,�̂j�φ��|����Q4��
�M+E�q8k[���N��k�u	)�IR���	�K��s)'@�J��t	����L�$*�L�}>/Y�FX�yǐT'�],�O�%�g��6vE���Oddc�x����,�	P�o�����޿������F�D&���9\� ���@	���*c�^o�,��x)�;ڵ$���Qt�Ur��]{?9-�:@;����k��:�R1kĶ��	���9_�[L�}SK�W�i�(�=D�������D��K#$���d�&���/����3�s3��VL�y��8U�=��q�M�\�N)	~�$�:��mj��O/�Png��	�z�̽�bH�Rʦg���S�M3O^ñu�R��QޯQΗ�C
)�k��W����waE��e�5�i0���d��=�{�C�V�1����%b�S��s^�̵zQI[���*�C����1P?pҋ�_ht�N1l|��J��Dh?K�vUai��Y?Ǥ"�D��lr�N�
�G�ޥo���cƋ�Q��J��b��P���b��5B
܉aom
�>烲�#C�ƈyɶ2�o���i�~�,z�a�W;�6~R�؈=���h%���ϟ}��!-|�@�[��&�[�,�z��Z9��(S�|�\�o�K}X��t���|W8���~[=נ�Щa��H}sд)H��\�W�������:���5EK4 ti�yc�ܶ�I��'j�9f�orU��<�B��&ƥbc'���X�WtWɇ!��M�vs(	�� �o�EF߅IB�o�K����U�`����
s��h��h@a@+f�uC�&�\�ܱ�&x�ǆ8J:ns���������eº�����4 ���*+��)��PM��ɼ���S����+�8.<ٛX�6���VN9��"@W�O(B*w�9�<�y�z�ceap���̧~�V�<�y$� ��ITz�^JÃ����y�I߷Tˊ������i���(z�>��;"�Dz�؛��G�*͖��7�^h����v����S�<h�"8N���GSٖ�ض�O�Uy,�W2=���v�H�m7��.%�B�z���� ����d��%����ڜoYy���R�s��#�D;�>EO��\TW{3a`	�)/�S�@�="Y(���	�|��Խ�J���	�]r�x�P�I�g)d�HQ'#NxJ�j� �����1 7�J;Ú��w�7yX�vP��,���e�L��+J��ڮ���1��=\������a��&�<ʿ��'
�K��c��v���
N�Jl�x����-(BL;�n�����s]�h���-�k9�y�+�a���-]0d����`	�.S����;?8��ajWҏ�ȏl��H������,�������P�z 9i��x��]^	��idM��KLy1��DM/��< 6֪mA�yX�c�
,�M�� ٽ�I؄:�R�t_ڔ�4\���)D�V擉��H�<����x1���Qh��|�Vw1U�}���<aSlaŪ%숇�ܬ��M��|u�'�8�9_�P�Cg~f�t�w�m�D mj!�ϰ����Z%E[!����^�����3o��_Z~�i	��a@*hq�kJ�M�H�<�+93�n)�D�yd�ؼ�:�Y�(K�ŷkC7˝���mkQ֬#�{Qo>4�jk<�������1�I�	"_�k]],�����g�<�>��@ʯ��KZ��$�x���a�9��G��ɀĊW��!�Ʈ���'0�s\�k�`|���a�7*��!5{,�Ұ��mK����#��w)5ܰ�v�-�o���8>��D�3�>��Bt3���@/�I�!�[���ɱ�mB�]._�V.�t�)�A�}��'g2(�0p
u�C~��i
�e2����#�ʊ�xMJ���q��������_�¬ɖ����#� �!D8rX-1;�ű4i���EJ���5(��7���m�xD}��Yދ'�7��$w=�f���+k�~�<cD>�i���²�1�\&��^�G�E?�"�tvY.��Xz��ub�sbb&th�����X�P�&�V����+��~g���a�T4��g�#%z�C����"���BtZ��"[�k��+WQp�`K�'ʪ<O.Z��>#�\j�O��L$��*�Iz�~+gi�%�����,�r	OT`P��W Zq�F��Qfo�C0��D�̈@|���}H7�8n{�����͕��CȇH�m���J�Ѷ��znWT�}���� g��3+7nƋWW݀���$���#4���tk7��X��h�Р�����N�Y�{�b{�,ڌ��!����R�˔&U���QJ�Q�����������B鑊>������ ����\�|��\&$B�R�wL�ά��Ǻ.#��dg���U5�/���3���F���}��|dT����NK��y9�&u}NxY��Eb)o���̰�-E{lϟƎ�"m��T��Z�&U�腳�Q�;xZ�k*�����$�9-�b'8��'�*a���w¼�$\c��R�p����I�\,�+ /M��Y����p������'���$�5�6�B*�r/��p������HrH�Cw� TD����1�.�(4H�����p����B4{�l��U�_5�m��F�S�w7�~id���d�T-����ǫ�)֔q�{T����0�)R4��@�����Ohl�Hp��3��5�[�?�}«�`Sa=C�܃#RFB�kym��r��-_O �"C��VB�e���MH�z���m�^�R�i��+����g4��M���Ρ�|���!Ҳ;~�nfs�jC�I�i�.�h-���"+�Kl��y�P4d�:an�`��w"�I�#����Z���j\$��j�4@�i�I��o,���So	�o���m�78J�l��?��W���%uYTU���0�Ň��#��a��(��{�(߾Z0s�α�Z��j�����+,"Bnz���J���3m�n|�������z/�}����&'N���VH8���Bf&#� q�c���؇)UaP�����������H�-���bNY3��l���|��|&ø�������>�6~*����qӟ`:*��GY���c�N۰��g龩]���E���r��Y���r
k���X�Nzl�֡Pq�F�@�\�,,2��\ I�+�nI��K����8ƾS��~,�+���S����:1�T\�Uk�1�������������R����Q�(ɛ�8�϶�r���׫sG۶�͈�W�k�N�Z��m�{j����+9 ��g0'as�~�N[��%i19�0諃վdr~]qmߞO��⻈@���T%9N�im�#�kaHz�R�r��Z�%��f��=Uw�!�G!H��Y65�0���܏@��D|�R�b,*�!�4��H����7� ���Q�T��$��U��$�sN��Ϩ?�GC�o�3x��eҞhz�u�P�����ߡ�vJH���m��]���xAB�^�Ѧ�Gu15��|l:sV��qϢ����Y$U�f|~�7}��D�0�T�깼�V��Ōe+Ư@$�M2wM�8�=YH�G��g��s�֟���R�����U�_y]s��i=m�ԋ�
5��0 K����[��E��Yc��l��V�o�v�	#T�� %�4jx��c�Y\��y�Ϲs�����.z���K��͑4Ƈ������-����q�����59�����p�D��6��/�����hGE�Jż'S�,�0��WE����)zߪ��&��n�ͬ�?$���r�eA5����&:Y�n��CY�@?�WoM� ��r�2�T� �
?JHn�dF�zKM�D>A��}��-1* ����]�_�ܻ�ӂlBv�;�KYn�9��;i<��F)��T����49�!����)k0,r����ql>�V�|?,t���Gք�vA�'_��������aΙa�	f�v��;��5��G��K/K[<�+�4��~w�K�錈.����V��$���mS�t����L�%&r���i��P�&r7rp�+�ȕ��6wmMf�4��𵱥+s�n��%3�)K�?��ؕ���6<IL�O�J��R.�(M�}QXʉ�y5Dz��Ԓ	�r̻�(:�.f[.���(�E�r��#]Mi4S"b�2��K�Yk:ޭ�
�-�C}(%�%�ߩQǸ[^N�W���b����`k ��������P���s���,�d�i�N^����g��E(�e�\��&��pv�u��߮����vMY`���Eff����49��]��l��Mά�D�*���K���AdF������ؘ�r0Xq�	�� i〟�$�w��m;Yy�7⁢�#�7`���P���ww�^�/O�"ax�ן���������Hl,+y��K���rٶ��f��Ct���#ƶ_$�b`���H��<L�fly�l�O�0�p�ʀܵ�kf���϶�uz|���s)��7�iQ���p��f�<:AS�g��4A�5�n��� �i`��"�T�D�mfb+i~]�/҆6��TQ�m*h�B�.�����-)��x�4��7�SS��#՞ZcGD�}���k�S7'-PЌ0�� �^R�H?�X���v�����C��b�	��~�� 	��� ?6���VXߔ�k	�m쩖5{lE��ح���J��M���+�ir �z,�����,�?H"��58�V�+���.B���0K�i)������J J�U�ѱ�q<>�t���I�1�V8
��8�����4��Goϛ�ad
��W7Q�]�#���%��"q\TL�f�0ot���OS�#�������~��J�]i$���ݝ��-/�%T��ܮ��p�p=�8�1����Η�[ST\���Rb*���0���>��=t��j�H�ഴ�+�U�j���yѲܶ�]@ڐ�0�A;�
��"_�Q��N��Ә������-�0̙"���M��fXH��xP�l���)�����: W7br�'.Q ��<]�u����vc#t��Uvw�*E��O����%׳�8�7 ݗ�K�*I�H�֙�Q���Y�B�T3�W�/]<P�(iG��G)�f��{�q�Ti�p,R�T&Y7o�`������D�DW��"���/�oJ�[�uhSQ�p���1@���)u�;X����n���f�u����"��+�_�ՄO�*�*�t�g�)JN���I�I�ɇ�%�{ ���JJ�(5����qM&tfS��%=�[�S�&����x6�9q3�섄-��I��sl^��8���p��	v!2���s�^���	�����m,�ɫK�B�(�k�ҷ�^�u�N��ֈ�!]�Sĳ 1��N�  2�aUx)�LIZ�f4���&JeJ�/L���ȟ�y�}�%��&�0�����_���I��?�S0�n}�Ҹ���C2�.�]��M�B6ܤ޶����@��+X���S�~x�eZ���7%`�R�I4:���B�r�('!�{�T��	#��+���yw��&��	ʥɸ��w��އ�TDy}���<P"x���g=�]�i��f9���b��V�7(�<��i����~���^X��$.�Rp-�hf�1�&�PHB�ǆtui}bCa�>j�&f�Ou��lvA�fb��Ԏ)�ә��|���a0�E��=��MC$��i�?�D���6�p���O�s��.4��Eo��f.O��"z{��M����a��/O~��f���2�!�L$�����_3\�-���M-�u���Əԋ5���~@����ݵ��5�9�4�y�Mh�� kh���~^�t�/�X�5/^�v�p^8��J�x��c��� .F���0���-���M��Ա�l�ho��L}�9� EԹ���u�I�U��^꿃���@��}���)���Z��z>D8#��w�ȫ�kL7<��sB��]��шAdT���\J�|H�v.57���<�#�6�l��L�L�/���/�b+`�/��r�Sԡ23	�M[��!Nt#���Q�B������3�0�@��'�:�ʽ��4ӑ�������4J�)�j|gbH����zt=�0s�����w!!K�?�v��FJ�E����+���Q��P�n�.�����q��mB��_B����a-9�cVt�\eWU@�5�N-����:K�x�]dMD@��f��}���&�p�:,w߇z

o��Ȃ�ln�e��G'����$��<�p���Q_�B^ �}��� �`k��Za�Ƅ���)�޶Yr=�Le�s�|��!f�̍���ϱ��b�-��s�i���@��A�Ɇ-����x]��)��?fχY���,/ A���H������\5�g�׹�̢���pة�u�h�|���o��7x����La���K�B,2�~B�yM�Gʃ����>��%�@�mbhX���mb9�������^���t�M{�;T���p\9E+t�{?���/�1��%�έrכ���'En��ō������f���S�Z���g��x����ǧ!����+FY&��u�r�Om݆ vޞ>L�Hs�ћ.G���V,~r������D�� +��ƴ�<ڄA�~T�1J���;30����&���^� ��c����p3�nz�aO,<?�Q��md�Mm�	4�#Z�Ĉ�:-�LM�qm�cŉ3^#��N�"��d�Nw@�ڠk4O�>�V��?��E+��h_fT�ݔ��VS���&cp<�ي4U���YJ�م�̫�q){��/�P_:v1.(��D�f�H���/��
�P��ͨ��&�`XR�����3��R�m��e	]�G�x�����i����Ⲻ�Z��usp�,�|O��)
�[R�]sM�
�Ɍrv
�E"�ͺ��s���n�pP�oKz���$)�:����kl�.�6\<�l�����?8�g�N�<�58����댩�-�6��p��A�6�V̲�E:�,�ܑ��KR�$Ƹ82px�J
���(���f�V&??5�1�?+&㯄U�d6M"���:e?ؒIȷ<�Ӟ��59"ҥ��l�P�c�E3��#��8db�i�I7j�\7i��}������0�y��~߁b&V6$o���F=��+d���m�l&NH��`�ᓝ�z�=	%������
'e��և���x��(����of��V@�Rb��bD�F����2YE��!�@��i��*�A>Ã�B&�GLwb�\J����_�f���^���G�6�w���	�k�/2�|�:�^�$�_��`Ev���6e�O ctѕ��?\�$�,tpg�q�Dq�gx�J����lr��4�}R��ǀ��G
9�a�=��m���x&�r��:��R�՝Ċ�$Ү��[# !z��X�@S$e���o��7��z}�������]t8"�/Gƫ����r;���Gz��f�~�o�n����R�Q�;I��۫ɔ����:���v�=��K>"��*} ���_�E�葉�8+�D��z ��p����\�
����%�}"�»8���C��p}'i�-��P�J��b:�w��d_m��#r���T�1H��\R��hv�r+���H��=�ݿ^O�'�Xs��$fc�2��qa�@��^��g;�^��b�e�{��]='��4˨ۙ�#��'F �2�d��#!p���#���#��5T�,����%����6��~�旔��%KÂ6���yQ��T�b��,3�X��r�~FQiQ$r��Nqh�@*���7|��#\ �-�@2,��B���9��w�,
�$��Z��d1j�Ø`/�w������<�9�\��Zk� ��kв�/��WVRYcȦ�Š���� �*��p*7�k�
(E�h�vΖk���s+b5�����<OGFV��L�x�R��u�o:��_2���yG_̫�k�n|r=��x�lB65.��qyx@/A�g 	f�pc^���Um-�ˇr�ޫ��wĵ���F���ݠ���@'��6o�4����j8q|��w�9�O�B�^Bڽd���$ bl[��+V޺� �&H���D#h�r��d���A�r�����ǵ���H��m���F�B��mv�RsJem-�&ĺ�9/�Kդ���J��f!:ڊ���e��T_M~)��� �5[��dP�@�%1A�C[�T+5"�]��� ���-�C�1].��L���h�$Ĕ�ʯ�y�K��K�`�r�K2rɝo���Tj�ߌ�\��g�t�Z�u��V��n������&y��ԝ��D�Ŕ�˰ �&8���!�8|� ��A�{mU6$���^�b�[�@a�s�ՠ�ôC�h��� N�*�N�8��uz�Csc��VȻ���2`�;�����_S�ia�VQ�omv2�iWzr.�����]�e���w�]x��'oX��"x?�z�80�;��_S)�\F���R样�ث�`S����]�S�z��Q��:"��F7��(Z�f�� 0�8�\�K���\,s0�/z�ȅ��ӳr㼈�r-f7\}؂��;��t�7|�o���X:-Y��,0�f��BX������1Y�6
���~CD`'0�r��z���Q�E����� t-y��+ڕH#���Kn�����5Q���<!SZ�I
]�7 ��2i�:C�=��)��V�pӰdx}N�ؓz����H�}�N`C��t�1�`��-)�Fx7�P����c�l�������'�HGGe?�!���p�9����q@25��&OL˥/��
v� ���J1��w�8=�<�d�BW]*�n�D�|&���bOk8�N���>�w����}[�����_v�_��?��ܡ*�rqZ���Ҙ�'@�Q�2VWyR=���{q��z�"��%4��P�6�!��E��^�5�%'�(�
!&pE���xv�7h�	�Ŀ��X/�N��F�����G~o͙K:I�^"'q���vw��d`0^��L-7�;f@*�D�W�G8$�mb䒃Q���:���@F�=+�Ӳ�.�s9O"A �>'Ύ�oFk�l�^Ŝ�k�J��,4�
���c$U8�2����Ys;�}��_�3 ,r.kb{�	Ze2�wH�p�NR����l���q(����%1�E���	� !�['x�I8i������]�>���1 �MEM�		�ڬ)o��\�-�����M׍X|�H�|/ߛ]�f�+o.[~(K�9�	��r9����"����\��.��%"��j���.F���Y�0���hui�,��V㇤��� �mZ�?�W T�2a�Ȱr��h�_W`}�����E�Y��!7{H2~����������[+��?�<������5CշQ�I�ĬH܄^cH��(ș�S%y��o��[V%�����&K̕<�չ���Xwvm���A��"*S�r�\���zGk`�͗k=
4�3��_��D�㘼���0`��=��ldF��)�{c�u������Zɪz�Q�o:8H��i_�r�gD��Q`U6���;��v�}���0
���pjRk�M���>���I_'���	ITG��G��� x���)�P�趇�f��؉Hy��z�|� 9Αv=���k�h_[1�x�GJ�vL.2V������������={!1:޴�N���|(��Ϯ+P9�l�	�3)��dׯ=����p$�c[���~�:|~(��8����1l���X����`S��$[!�T��PL� ��+��X|�i��#(�������!\Ѩ���e������8Ɇ��oA1����]��6���f�r�c���ӫW+Z�P�Uѭ^C�mWN�ބ�����mx���oA,!=�_�*��-2I[Q6W-1���P�jj�^��Ds{������]ݱ��4��y�/�v�G:�\��: \��PYEr$Ǳ$肼�qRZd�+����C݇M�G�:t�̋剏��;D���U��S��bF5M|��;}B��P��K�^��NDX��V������J�!?)���|9�=%�C�V�u3��WEi�L��պ��E3��1�s�=�P8���k��3<!��{�E܋�-�ކ]�ˮ���	�K(�tALFq9MC�m@����CD"H/���Js�2&�BZ^ʾV�ik�#͟��Bs��%�6��m|,�6,M:Ӭ�J�ER���dHdy�7�=��02�WXZ���W!�G�2$|RV�ġ,�$��5ݤ�g��_�\^�����#�ހ��U�38����*�8@���ex>}o�>bDC	�i�Й���y]8AǼ���T��|��2��"��c����4e�W�JF�C�,P�&�<0�0K�$F����X�9���%���Ԙ�i)�o�l8%ο���l��͵����� s/��W�T�{�W��Ey�ҕ���̞6
��jw�������[Ѓ��~� ���4�O^	�����mo�'v5��Z^�qC�{_��@G���]�W`N L��$*��Q1󽫽��6n�A5>͕���>^���s�����M!�7�|��Iu���7L̕E�sL+_=�4�j�ߩ$mkH�J������fV1�� :,�&�7�3�l
х���¶��Dn۔O.�RR96 �H���Lت5�2�{������Wm�:��i��2��Ų-�+ئ�v�\M\םLg8���0:P�kV��rN&
K@�t[
䛋^m���tɌ��/�R��s���p��z����;�D��I��yv�\O��9��A ��a��G��.�����v�	Q��}�uš����]�����i^󹖼�{CZNK�X��'�z�}�\�}�w.ӳ�w�@�,���o�((��0�ra�c�Fy�B1�ls��1�h��b�O�1<�U>��
��hۜ'�t���� ������ ���0%�Bs�z�Fq�i`�ǫ��e���b�T��[�ʊ��R�81�f�C��l�R'�� ��Y1��1{����Z�W�=�$N�f�z1č0�o���v�Jx������pP�"���zA��`w	�����m��(���5�ʔ�����#c,�DڑY* �k�Nv�_8Դ|x�lJ�+l�v�|	jAR�g���d���y�[u���(��_��Tb�JY�Ht���g�4&i��9�^��p�RI���>g�ݻ��L&�F�F�iM��rbiC<)/F�֌�p�Q.��G�z  @�ng���h�@�Cf�^����-E��U�a;�D+�����qm*�)����p�����ozOs*�b��0��0�{��sV�Io�g��|W�P���I�2��-���Ddf`;.�rިo��*�bS$ ���@!�<w(s��I�m9�:��T~�[�p�Dj������;�\��}��P����C8�O��Cơ�1�訁
����GM�6@��A1R(?>4�j������E5e���� ��e�_q�qQ����ùz���iDE �P�M	�CY����a�HU���n^eU��A��km��~<��;�����r��3l���X-���L���򭱱�B��+�/+��V*7�&=S���J�c�s���{*YhP
��h5��o]�Z�OK�T:�ƮX����9��[n)��7���2c��0��.�O�H������^O��V�̭��ΨW���I�Z�y�M�f���8�J���/e�lȯ�����������ƽ�8��v�Xy�7���Y�1��uwd�]"�o��#)���
)�>��R�B�#{�sZP�b�����4πA��)� �khy�Im��1,�_�*\���]�fFo��?���sT�Ld3wI��*�*Jzb��)���p�;�2�3x��?��藖��o��������%NE�x��k1R�͚�X3����*u��p��,w*��Av�b3+��H?��Oݸ������i��܂�@S�Y���V�w��T�&��L�8_纥`Fѷ?8S��������G?�:�>��;�W����15 ����GQ%�W1�Ρ�t�0f�	�].�*�rV,]���o���M��fqg�ޕ1
f�R�f��d���=d�B��PZNr����i9��;S�¯Zyb���40�w���k�p��a�,��5\f}Y�w3Xe���sC�e4�슁q,���R$͞�ޤ-��o��f��&d�q$��!�"������!��-D����#�R��ϛ�u��� -	}_�GyJe�ߍ��Pty�g�d��]7߭fz�t2�2V��%�I��d���$ҼeL��������8<�e%��u��ߦ�����lT���{���VO��!�X�pgI�R^?��Q��V}��'���X���rH��d7Q�PM�(�Ϟ^�]tv߻ͰDaヸ�qt�w����JFN�y,{�&PF����������v՞����c�3aG<�J�$o`��Ә�8;�Y+b��^E��CPk��j�D;0�B���͸�������ׂK H��2k�$:$A�����e-`�h���dPt2cD�X�o��1�C�ju�W	���M��Cی�K\g���z*�K�#,�,�4"鈑"4��9�d/ 8�d��&�Ġ}��$5u��U-'�.W�x��<ީ��*�r���Wذ�C�
j��'#�g�8A�}�i�y�a�W����	-��@��2˧�cm�!ކw�PG����<X��W��,"��[�n����Jp
���;;��z������B��Whm]/^�N����;=��+J/H���"i����+ *y��q��sy��*{���.����=�fl�]ea'��t�]4nZ#Ŧ�e�A���}"��_�g�����$e1&V���N��'��2��}
�r2�X�!6b�?��W� 6��$m33��ڴ�#�|4�5�c� 
��@s�FX�.4����9F�Ԑ�r!�t�K1�O��ȶ�˘�uɅ�ܓ��}+풐�\�2��9
��CЍ�>T!�ouJ�&���1[zt¢��|DTiB�'	�d�A��o�����E�"��O��b������}�7ܯ_���; �'��	���X|F���eVup�ʚ'��/#�U=�E �,[���x	�ݧW��nJ:<�zVF��h	��P��h>{�q��t��h���jyp��!�0Q(D���#�bd��yc�j9��%�dSͲ�Hpӯ�#�#�}�q��4m[�1.z�K�T�[�����/���}��S��vl�.��N��"o&�n��x
�ġ�0:l����H�K�_*yo����-}��"猈	[jq��N{���&�T���	M�^����6>D��y??Q3ǌ1������OX5z	�!A����0+I�����Z�k*mu��S�0?�ٸpO���	�h�� U���~Q��Oa�pפ�jP�`qY�1�|̛n(�P�{`�XL�M��:z�k�]ײhmJ�@����SD�}��M9�3޶*ӟu��d\��]��!~kV��@�9����8s_�Ky�(u�.F4��w-W�+c�-:`��
.�A�+^���(5�~Y�|��BedU,�dU��̼F�d���Y�+�ٶI��e���g��ٙ�O4<��{�ʜ�G=���0*�f��%����%�m$�W+8S�u�7xyy�;��;ݹgͧ6������c ��ݺ �d)22Y�#Õ��#��޴�F�B�H-w��P�&���E���.�9�;�W	�M��7��:�����&K�9��s���+`u�[�,y33��Y�����_��S��}�E>�z�e>?�x3���y� !���%C��]NY���#鿗��,i<���fE#=M԰Τ��*I�,Ȣ���O6%$�B(��*����?#��9싢&��V�x���e �c���y���|����c psՇE�.`q�m�+*�{�K���u12u���8��z��xw<��2=�:��/,���bV�	�Ѷ�o��+�nT{0 q�T6YX�G����o[�7��Q-R�9O}^�.�y���X��f�=�)HDs��n/�ږ&-�9=�����͆�	�����D�bJ�J�
CD��bOL-WU�>I�Y�3}�\S,0��l�V�I�3+χ�� ��Q����?�Y������]S'�ެwdAd�4i�6����,w�1�iFd;�Yf�`�%��I��;��lS�0*�iH�j����:=�G�<Gſ��k	qh)�Qz�S�P�7��&r�w��B���Bխ 
굨�V��(��GdW��y�r�9rP�3T�����2mEy=�Ck�R`[���8��L� ��,�_�{��9�o�V�ق�K�5�'6���2 �H�k[��h2�`*�]A�)��2��@9�K���I�ZE��8���W@��[?3�՜& }	�q��[H����/�!�i"zR��=�+��ጬ��E�����?�"P��[wY\y�p�fhi�
��ݳ~�l�	;���pq�f�L�{�0�v�����ZƇ�DMP��ܡ�4z����~���¶�㘪|y�D,��"�-T�K�)��i��
H� G�1�u�É7�����V�B�gH&��
*�X9[P#���$�l�H�l�.�Y��G�Y �;��ÆhD���^lT�Jj��r���2�*H�3���x0��w�F/x���	���"�3Č��8�<�6��],�瑌���_�����/�*3�$�O�_VE�U����Ҹ��P��7~����=c_�H|>i�R�\f���6������k�5�,6�ьrM�,!���S�[�[F�X�Ԑ����3w�ؓ��O8�r�g����JW�����66,BF
�N),2��m���̰�T�ur?SxW��tO�����=i�=0���k���*v�uGd S�AƯn�Z�3<�<O�烦�$�����V���:��CiԳ1q�/G@N!��Y#��N}�iH�D�Eм-0~xJf�ve�ܹ�����"kCqSP����F-^��eg�r�U�Z��D{�<t?��5�#vh�_HAx��\50As]�B�������_���r�W휲���ދ�d�k���Dv�����H���m�ap�W7�v��IH9�M���;vĲ$a������d���׿4�.��}���k�7��m��-T	ȩb���>�L��?�Z65�5�%(b��Q2���u��MC:<VM�Pfx����V����80�w�Y0(�����K.E�$�{�~��X�[�+��mɿ�{�git��0���s�#���2}�PPە-�|�>:��* �O�|�$-E�/��yo9� ��ӑ��z�X���L�?I��#"���v���tژ��A�Κګ�R�Hht�|�k|����7>�������:�"�Ew^��|aՇ�������D|xE2������� 	Xf�&,�g�&���~&���\7���t0����Ԙs�s!����D_Al�ŗ`���Ն����W �;�=�����|,��$���W׶G��z�#���_��<f�r��T���7LS����K���z\�L
���4w�X�T)@��j��7#;�#���#p����j%������%���ٿ=c��+d�+�跳�ϸ��{�(��J\�,��)ee�4�ypf��r)�cs��aC5ؖ0԰��~�% Ic��TsY(���As3�D�rlZI�#��1A�/�P���R��±;p(`���Nk����l�&�Օ���>��	/�$���=\���֭x�֏/:Ě�R��
	X�an�Q�B�Mu�P���ʖ�܋���<(����y��@M��d��$y�s4)��}Y��b��kk-�B�@�n�F�-��J��2zR�<Qs����8�S��S�XB��\
g�Ś��
��.x{��74��+l�=d�CV� ��;���<	(��[��@H,�0���T��(+����_��ŀ�OcO�4��Eu?���fW�=#��f�cH��u0��  ��w��t	6���l2ß�FkZ:3�3䖌Ӂ����n��+ع�ޏ<��\�Z	�`D��fMCJ�UW�w����w���o��ɷ����Y�]݃��cQ�>��%��c�p/!����/J��^@�$�d8�T)�u/�_V��"x#����i	|�m�}2�X�^���LѾx%jö��+�)e����F[�fJB5�#D�L�M�N���n�-�8�y�T���z@0��<�xm��r=�B\e��?��H�t�>��!�_���S�<�,��OL���)w�2���i�x@��J��&��h��Pw��,�n*�f����;����q<LQە�A��w�dP�ȮԞ�D&��5��%Dų�\v5p�:aoA��_�	i
~)�4���8�+F�fp~x��K��N�b2�ƾIt΃ht�NBȧ�54��z�ި�T�Rrק<�A����Vb�\BD{3D�Y=�?��_@�}ݽGh���m��b�S0P��G��>	�v�x^�Oa���k�����1Dt�4��G=�v�~$ǉ�C@��Z�r!D�U��a���Dgc_PH�ٰ_�?�+�j���r��{{��@tY`&Ff���7U,�lg��FI���Mf(���/���
M�sZN�xk�+F���_���i������0�yI41��g�k�Q�-��[>ϻ�t�cv��9ny��8�O����4+�9&qַ���y��f��K�Zҭԥ
�a�=��.�AJe��O�ę(>��B:τ�Y�	_<����ڐ�4�~]��W8��yȈ0�a(���k���/:�[Mҟr��nur� �//��鵅�]��}� ��O��� �FU��|Eh����"�@�cqUGUHuj?zRdI��^.�����p�T� pp� ���I煻Ni�-� �]�C���<�?z�P3l�rֳ�hq�"ىve�t��L�Kﻦ�O"?*��X	��XZy��A�Hs�6�u��Z=���^I��*�M�e�k�Ṩ?ʢ��� x
Ӭ�~5�\�
Ƒk����)��c�����y؃Ŋ�ngH'@\���c!��ȩ}�G��f)��M����s���H)�pf�|\�]	�O�,	��T���~�x���nX�ڂ���[UJ�!5�9\��ӹ/�'c[=��ji���̴��WK6�y��-�8� TvB,�����ZY�a1P<�G82f��0MO��_2���>b��'��wsVw7�w�p��"7��Y���ݣ�D��Ц�lͬ���VC2%苡��X����N��;ЁčA����$j�0�v�� 0M��$&�����%i��W�2��%��6�珑�'&G����k�i�.����zUV�cK$M��_oL�a�8B����q�A[�RǄ����?��P}��^l��!"��� �
i�uϨ:�����4�E�҅d�.q^�����˕B�-�>�S�k�#�c]�H{U�s<+ʗt�ܫ�D�w�DcCF��a5��07+x�D�m�z���qe9�]��sց�:�+y�c��� '!��6�m�}n>��x/P0�dj�����������1��D�[X�9���eP®�f�����=ۨ���>zJ ?� &�)L�A4�=�)T[ ��|�Y�^()�C? ��	T�D'*�v|�c,\%�0�i��+nT����h�VҘ���9g����$n��4�TR�I�H����е���������Bb��p��6�y_��V�ћ���2��I/a�M9�MȐ��z�)?��|�8q�"U\B�����&�%^�#��j�������q+��%��E=x覾\ʅFj}s��M�-(� mH�T8��_�5\�.��C_�O�s��!	�*�U�ɮЙ{��i˽���bi{��2h�:洳7w-�?_��j�ĵB���g34�QI��WQ��r�{��M�Lr�m2����}>��|��������e�oT���CP��'���f�X��vq�ұ��� o���ߢl�v�6�Y���σ�u��"$��~��ԑ����kIl��ՠ�T�6���<nr���01Ekߪ���x�"��"Qg<H���y� )�!6��e�(�(dUeK����a�P��OV27�'�Y��BG�����f�̍]�!�>-���������� �q�:��.�� 4��z5k� V�!�u=S�L�q�dO}�~�J?oe�4=�6��VW�'ml��Z=�[��y����j�T�Q�TL���G�X\��������!Z��?��d��y��-im��ۤHU�2��.L�z�u>ߏ8?2�Eak �vdV(����F�.�����M"��)>�ᙲB��_�Td/�R���~��H[HO��6�ۄ��!��#�Op��Ѹ��( �/ڪ���O���n��w:��2qbd\�}����E������G���{�`5�(��}k$G�"�>��6�8F%TsI<{�D/��!�����z?�I��T�W��,��[D;I���Ǣ�J㑝D�eD/����I���'q��j6���3a�	���6�fFZ�(�b�Zx(ӈo$(&��YW��Xİva�� bnk�NT����iCv^�]2˸����O�j������K�C���9��Hb���N�{���~��A��"����vǋ%jP$�����{�qZ{�	�$heQ��(�BH���Z$A⨛���MhoΈR5a�="�
V-O�j���eƐSǜF���3;�_J�≡����d��pQЉ\��2��B~�pήU�@O��0�����Q�LL�H`��˨�.�h)�J+X�l[��{\џ>�)^�P'n�W�ɼ騗������$������ �M#�n�tu��J�Ff�JU3O1g�11�tIN��@[K��8���gUT�&��v8�Dӈ:���Ŧ��-�ܥ�6j�S��K���R6m{�K,�����QU�0W��@/im�3p)����$+�/���hXJ�P�C���Ud��%��;�+o�~5C�ա��g>9��]�7ے�}�#� �	�G0*�	i���F�cx-aӡ�LBuH2c|�gt��1���3�~fh:��"8�8[����/�o��,����7��{�BJy����煬l�3��2��� ��+	�Ⱥ�~�-��@���J��h��mC�#9�%zĚ˘�'�'�9��q����n�T����,U�o�XԷV/������ũLp�ԉ�p��	X���f�����S@Ļ�(�{�B%��2�N}PJ>����V�Se�W�v)����p`�M,H� D�x2�`N����B�O�lKF�e����0{mLXv�4FcV�-��.T�:�+���I��������K�˽xeE�&��+�&�ɬ����,d�C�3:�R���'�ގ�-�C�\6{��m��f\�����'�}]�Aߦ�����B��tZ�8�}l�l��p�r��"C`rD*D$<�C;�0���O��6�>D֏e<
�ݜ�E�pʛ7�Eb��A�&���^����^�8��.{�k0X���{F	q_���5$�W7m�֏-�'�Y^�L�v��������e.e[�[�v����RX�s���~����j./��}�ک-�+B�,O�2[�8�6�5E0����26g̏v��`���J!J�>�V`�#�I�X����<��F��^z1z�|mK5��u��2l��%��QƟ��Ĺ{�������X�b����^����d�����e99�B7Z�+0����(c��u���D�G#�#�{v�*E�<�� ���������"+���m��+�)
�k%X^��'!x��N����u�!&��rt���˵�m�j��TW(T���C���\�O"]{���WB/��]���)��c<��vJ3��Ëyc�bD��l/~��ȻG��-$�d���d0����W�	�|�2+˶绀��e�B�dmW��ϫ�R�%��g˒g�ILyu��y��q/8�oi%��7��켶�'E��daI*��L11kA��F�}�s&cڊ�_ܵ����>ž�iQ��
T[��wvR������q�eM�=�G6Ǯ�:��B�{v�A�����#|HХ�$7#R#ҹ
��.Ana 5��\]4�Y��a��|f2^�y߿�g:q�s=94a��H��[pn�Uwo۟���-J�� B��
��H�
8U��
�����J�ڳ�G���,�(�~w��*M�uK�_q��kj�T�"��_s^9	ݱs��I��! ,�7��E�o��� LE��b_�v�R}F�x��� `���-E�ܛl��}���F���+�4b���վ���^,�q�_����`��>���7�c�ɝ8>�g���󻨱&��މ��8�?5 ����:M�"e��֝'٩��8I���5��ݣ)���`����  �l,�l���t{)��%v�F���y��i屧�|��x �K�).R��7Iࢸ@&>���8.�;�.�۷h	i~_��D#�t���G����U8�)4W��z>�uS�5)�߈%�����D�� ��� 2��A|�a�M|OM`�e#��g�q�p-��zZ<��q�jOxP��K
�9����������	4�1��g��7�Ƿ��5o�˺h��L��Fp�7!�SlnH�L��?��	�\T�hS?WuZ��m��X��K`�a�
H=J#>-_,Y�򶤄:y��XXl��:�*�86Ă�c������:.�#|�!@+"��w��i�Rt�81�98��ɠWZG��(7����
�KwPF�,�A��G����	��W�*��|d"�X�R��fiI�<.2��j#,1�$T0�#"��.ߎ:V��.��y�h#��Ms�(,�-d�ef)��Obt�x��G�	�)'�-����l���އ9S+�_�QF�"X	8c�w�Ϭ>��Ion���kI�֧�=��-�Z ?��M������۝Q�H�ۜ#�ؘF[㙿�Q�F���_3"1���/���"���W�܇�"2��;b���F+�	�{�>0N[�ry�L��2��"�TN-[�|?G�KW��Z��ޥ(��	���@Ƣ�h�������E9"���f��p+ݱ*q C\����!IUR����6��Ԩ�9��|�B|"e��}^�#S��l.yt��<*g��g3���'$?��gd��˳ل/^�^�����|@ `�5��ؽ�B. _*����tI��Ϯ(�-����x�>ÙT֮�sG��q��ũ[v����!sZJm��&�=Q�!�l	lvn�*͞�����A��ز��ݱػp�#��`����٥T�X�I�����'ot�Y-��B�/��zKzϕ=��g1GVv��[�'��:T-b�>�^�ː�8/��E������������3���H��V�����f{�O��;X��|3gy�0��UQ<,��
�
q��%��H�[wQ��/*��a�_��Ҝjdky������TDVBx�$^��FQ9�\�Zl�+�I�T����fa��5��a�K3���4[���������y3��������ϡ��]�DK�L}.0��>z�ʍ�ډYq��[lu!�8Z��r���j����4�β�f;N
�?��:H�^#,�����7� z�����1���n��H��m���#��WM�؛y��f�9vD�?dC��?p5���f!O. F~�)5�f�a6�~+Y���m��;�����T�����]���|�'T)�C&6?�0�˄���-��<��z�;��D����wz�TO��&��y|b�2d��|�=��-~P��B��8߉��͌��eT�<]-�mc��9�%=�HU| 6�7��;%s�;��ä��Y7ʘV�W�mEϮ] �����K%B�W-k̑'��Ia����}�ޒ�[mx�{b� Ξ��n�&XG�N��eS�򠽶�˭J[��]c�c�����Y؟k��3���%�
�ݨ�ІU���cy��-���K�X~��h���E�,� |�t���Ց�A7\���ui+B��+z���HL����)z�|����Y'a��lP
�%�"�UtީL�0�|�ʠ�D*��h�1��ݳa�Oc�^\:k����ʲ���f�/�8���1�u�fe��F߷`�FGr/Z2>U��,�����п<��M62�MF�o�k�qI.��_���P�'r.X�?ne�.N��ZSH��g6e�ɹ�a��<��[����\.O��#�����E�()sֳg��PU%�Y����02�M�y�9�"�cNڙm�A@�O�R��2���T���2p���2[�i���?T&��9X�!�6x��H��O@�e��ܝ�
R<I��E5%�~U��'U���qk�qo�r������@�e5!�=��8�x����hp�]�n����yith}����x9äGc��v�d�$�'�^���~�_�D��'��d��mj�X�ti����`F��2�������y��I�4��14d�p��G�Z�N�h�g\�|���B�K��wְ3�hM.j����߿�<,��w	���S�p[����\}hͪ=KEa� ���n�%t�+����7Ecɖ�Y�����â��c�*��|���p��1/�_py*�@��-���Ex�|1I �[R��~��WO��������� �6bf�����`
d��G
S�8a8�68%:3S~���0�s��e���h���$�F�У�+9�6�Q9��~G������"�ѡ-�U8��$Q�''���\��d�C�5�0|'������	��|��;(�p�H�r�q]�]]�<T��7tD��3�:c�Skk����T�lgڡ����3��%���4���b�x�u��4{n� װt)[^��p�}��Pz�*�q�հ��B{j�A�5&{ϲn{PZ����涼r�򍔛knM��3�HHi�詳�/���S�ހa£�V��U��ȯ�i_�vʱi����HP$ҏA�R&�	���`�β@���zų���ܵ��d���P�g~c�c9{4թ5)\�/��	���35���ۃ�o\�>�ģ�X;��.t\zHF'x�Z9��j���G$�S~PQ,12�{�����J��2\q�
����^� �H{d?]N`8n �9�s�Z�+T�.���?�pF��	�1�n���k�ެ3��B?m	�t��2� �� EUd(&�)�kۘ���΋fAMr{h#R�E~� ��$|���f~�+�2��l�s�N�m=���}σJcp�VJ` #�{�/)9b,ѥեNu	zY�;����G��X'a"��y�.��s��nj�Io�OAo��ol�(V�k��v�	E���+�w�l
PԋR�t�&Ԍ�6�������U�!�,p���a9��\)�f�r� �A��Hl��4�-QB�"�@�F�|�1����S���(�lB�{���8Ģ>$J�t�F�:Έ���޻�����^<��7P��7KX�����=��r3Fm���b��]��#o�5~LǕ�i�ђK��l����ۍ���L����R���v��-�Y�QS"��!+�7:⁇R���?pZ��M,�&t��(0�e�q��3`;���*/G��xNR�B"�Q{�kʰ~�*!)�]y[_"z���8_�P&E�L�I�D=91߅�O�.���+c��}^�R�Y�V�L���^y�~��W��o��?���{�w��Z� ��Ú��Se���a��Dp���lVX���z�Į�V�;v�&�|�z��,�:0Lފ��nF8Cf��'y&��*���������@8�<%*��O���xMJ��mXa��a?�l����\�K\_���������~
^ר����"}�I^FbLE���~�J��L��/ �7آ��e��'�M�`1��>��<9V(�;8���W5��m몿�Q�!���:?Cq�h�(�S3vbBc��.݃�z���
,�\��ٶk�����b� &{0��6e�g�r���ŷ�'Έ+p`� ��>�.uuT�ۍ��֓��a���͜��]�E�}��#j�5�J�y� Q7�-hgQ��� �V��iPk�T;��mc��ZDw�!L�͖G�k*}ֻ�i�׻I�E��/E���A�#*�����)�q�gO:"Ą��7m�Mro�}a�O���17/��VB���z�.�<�x���#��7(S�����uA�RB��+(�#��kZ|���v*r|�qK�PXտC] TQ��(r���џf�|���
Mq�m��7[����l�"��{A�b{Q5�wO+�	9W�h�I�b�M�^&�����fyJ�� ���͇�]��# �Ň���bs)�Ma����_њ3�s�3�-�05Ө�o�f���,(����¾E���p���bÖ�X����\%,�&�)G5���d�t������7�WdpQ ��i_&�!p�f����{�V��|{�0�:hᣆa��+�z���j����]`��5�GE8gOǢ�VL/�Q��(~�g+@�#G���{��o��]�D�QK����2�y	���<�	�+׈L�(FmK?�S��l��߅g9��j�W.1<����b�C幙���Q��j�d>,M���=�u�7fG[$x��X�Ȃ��\@Y�uA���"��^-lx_�?<`�$�@���:��y��A��z�m'�w�3�~g�i�<��@4��7;KI�
i6���W�fvc��= �f�~�+�C���z����0m���9�M�����q���|��H�=�����D�e���*��r��ϟH�4���z\�D�}��w� �v[y��|�E��d ףC�����K������8�Ev�p�Ԇ���޷��_)�a�Yz��vp��8ұ����Ƙ(X���(�IA�H��Q\�4>�o���ʢ�1�Q�yϺ�f�vu��IsR���DN��W���Ȏr��q�`�>WR���"�q���%g��Z��Lmc\%`�1	�Rv'y����PbJJ�w���&X�BYq}�&В~T-b:W�rAp8�R�\b[�Y��$Ի0o5�`�@�t{��Bm�4�2��L|'e ���$L�"�+��z��9�	=n�&�n��İ-8i������е�]p�!�5�?'���5?v�X��3JG4��S�n�/A�>5�%C�6ۨ59)/��&<�p�E��1y���$C���D���BǤ���E&��|c��~�Z����f�е�.L?z#z�|z��U>�uu��9����y�y^��^������%��4���G�Bvq3�i���L>btS3*;Fj_��h��оP�lS�U\�3�W�4��Z�.�#���ߨ-�A���s;��W� mC	�Z���M�p���|W)[Ct��t��U��SMo�
�-3�4��ɘ�d��m�3q]<�6M������m��Tӧ�-,�.���r,;����
w�D"� a�O:9��ĉw�B޵K'�㇔X�}���c9m6rt�}���Ȳj�q�/p]�ck;��^�(@Sn��A�5ߗ,���X��
�y���ku���m���6 f�´u�&��8�AM�^�:�iMs�7��PߒVe���tb�$�*1&���5�o��`V����r��X�)��91앾���,WS�4#d#���ܡ���|UX$�(^W�ڂ���c>-�W��ս/d�M�kz�/���t���o雄��������eZ���QvM�(�2���i��*��M0��M����LZ&�L7��~vjǅ�t�ʘ��<�]�A��n��q|˗dã	�m@�� u����W o�y�釠�N�uGV ��Nv$<y�X��YNS4�s����k��s����Us�0Y,�5�fz�D�;h�l�ѣ�?�k#�U����Yt���@����?�tx;ވ� lF���0�����h{�+s+�j�	B�C��t�Ϝ��5tzuw�Lg���Ʀl0*@�7F�빃6-z�-���@��@n�+��ʖ�����x����YYH&=Ҫx�=�-�چ*[�(u��k�(�'�0��^K���%����}��.քX�F�fj'kPP��u�+�S%�Q؋�Z%SȾJVD�>�r8�[�P�KT��<���
�gE�������:(p;V�ʞ�ǯs���Ĭ2|�!:4����yi��E�t�+��&��� 2$��e�e;T[|�!���9M=�wa�V�3�L����*�A��4�Y�r�N�&�k�h+^�(%�P�7v�4x�{��'��Z[jb�;����ɔ�ۨ��s�L"��0�sĽg ��Cp�zDy�?���B��xe�{l^6����%m���A��O�jx�G��� ��u�^����� Tܸg{۲@k@���Y����.���+��%�H� &*Ȣ�A];����|�M���2�l�{@[w��:@��g�u
yJ�,�R�i��g�y��uX�_11h��ƀ����.�	h�>�pau�K`�Aߥ���l��*��n��������BkڏL��@~������Rn]$�}Ia\6��x�ܑ�'6P%�:R-_!x�1L�����Ȭ��),�C8��Ss�$� ���{ϸ�J���]��;nx���9O
��;y"�pl�eeTNl�O{O���Br�^�^������͎`���O_�>��לB.D6����9�X���Ə M1z�b�]__�Ԁ����&�LMV����z��+#���9M����}�e���eoT�� ����X:���D
�1h��F��0�2 �ն�{��e3lft��Ë�_{�m�
Q(&R��c��@#[Z�ve��U�'>�?���H��H<��EV����ȓm�j_��bT7�H��� 		u���|M5�Xḇ�w!�{Z3��=�J�E��w�.�~	xk�l�KE�`�ߨ	�dV+D)�^��C����������ߩ�%b���2x�� ��"�Q%Hd^P�԰��q���%��vu��)LH�F^�C��v�f�{��$����;Dw i���#�%����2j��U�����k_�{Ú_�9z��4�6i����/ȷ�� �;�؝�����VNF�-S�Y;�[����n\����Ƿ2�0-�Pc+i��/���3����(Ms��`y0>����픲L���z�v2�h� F�RΝ�(�{u� q�P~���Q' �(`{qQN���a+�s��B+q���l9�7%��� �tF�ˇj�ۚg�.I�(ٓ����HNV��\'SPa2I���H���;Ŝ2��?�i�w�E��Rw���0��D�����0�b�t�$	�R�y�o=�N��bQ��IE:H
w��k��?��}W�%��R�/�JM)���N'�BR��&��o}�xvT;[v�&��������CyV~۵�+)�w���Z���3e��8U,f�ۖ,�f�{U��G2�CE|_��1���% I��۵iӑ�>i�ڻKq��Z���cs��=�0߲�b"NÉ$�I�H37P]��5LG#��i��<-=�1�8C?��0��D<tCU�р�#c�7������&$�0�!���4��Yr��z�2]y��tXl�2p�aq�V,�	s)3���Դ�Yӝ��� *����3v��:3��l��X�ڨ���)u���OQ����U�]7غtR��l�n�?��,j?�g�҄z�]b�4��	%�oӖ��V`4�'�.�̤������J��75I����v�N�P�N��[�]�{%���%�A���u�IbT)7#*��'"垖���t%����^'���y
]+��쉜�7>#��3m�g{��E�mH+,9x������#��Q�"�Hl$�jHP�5N���y�9)b��y;	��:sX���W[�̊^��+�|;g!���S�ǐ�gMl��=v�x[��p��
������,3A��{Օ�"�����AhJ�� ��d06z3䋵�xU&��p�+�� ��E���F���.YpJ�������*@�T��T�#&������"+ب�L��ve�7���N+���,�_���_�M��3�fiQ���J`�i�P���H�;ǳ̴�͵Ma	w���}�r2��f��km�*��v�op�f���=:3I�*ڮz�6+��^P������V1��,��"+�՝��zڳ��o�QX�!|�J�झm�qq8��������@?��t��q�$Ԡ�éx:F^������4':�h�<\��HV���|J�V۬M��[�s�,�`}�T)�`�Lc����K�QxG�V�f���L��ƚ�+Dr$=�e�y�zX�-`��	��5?�qLH\l`�2�^aa�ox��Ny�{��'f)�oh��@55c3�`6|��=�
+�'M�����'�Ҏ$6��C�
�����z~">�)X�Ƹ��/�������ﾶ֬"�9�j���<��˰ �����nIŷn�Κ�C��taN0w	Kp���6�\N�H��,�(��Nc��&�������Ȍ�s�Fo&E^C��C�#�|�,�I)�i��6L�!�%D��7#rY�D���^Ύ@ �G�1I��Ͻ���C�7�1=W�S1o���7$A������>���<+�㠣�\/�f���H{�
_��EI3I�Ig��Df�(�U�|5w��٘�Ju$�h�����r�hf@P)��Q��vPQ�ɶl��� ��A(6�����m��+Ǔ��H.�d8n��m���ʫ\ʏ�a		&Zy��Y���!ݖ����1��ʞ�w��8�q'���l}T�s�Lnk�Y���a�ҍm�/t]p���,��u�n�������o��CO>���f��C5�Ϝ����[_<o��C�W����ɳ(F�E�����H����+.n���*+nh�I�U��ָ�Ei�FjT��H}8�N:��[D޴
!8ߙ]�!��L�
l_���3����h����8�X޲'%7��y�!]�9srmT�wc)���R�1��.����O��k���=8|{����#=��R�(Ź��O���$$���]ma�qئ̞�-!��=I�����AF$�u�o����\d:�!G��]�j��.�|�&IzH ������.����S��?��xZ�k$���gs��'O���c�F�)x�Y�.Eަ�����Ԟ:����5w 3�u�P��S�^@�m��bć���6h�jYqX3"'�O��c�yȻ�&{�+�U^фo�������!�ҋO),3�����3%bJ��zP5(*#O#tu��g!����65�lB�D�f���Jt�w'�1X�˨pפ�%Qd�Mr�(����t>E�0��$Y^��x��TV���~Gm��,�y�-�*j�����7�b�h�ː�^�T��,5zI&2��a5�G�V1a'���d��}��~��� c�g_�o ��Zm���b�~1��\?��`jJ	�X����̷�SF��ȿ��1ώ��O�i.9	8O��_x(��؎�F�&3;瓈6An���G�� �9�sו�9�M+�C#�V���& �h�p3:�dF�9�hu�Ϭ���^%�^J�.�v�m��j�~��`�����}��t%��/;�p䟛�+�j��R�-؋�H�8�"Q����EP�Ce2Oj��!9��*�S$ 75���|��v�,�$
ވ5�=C�����[�fU����i>�^����T��ԧ'���H��N�k�DB�gI[Q���1R�D]D
���SY��p��PB���3��o��V���[��.5"xe�	�O��j<i-�R����V��� �n�:��?�a�4݄���8(��M�K��`%�b� ��d��tY�j���Ԧ!�ų�Ww�1r�[y`���K�!v�L̍d�ƴd��6X���`eb����f�t!_�װYC�R�ft�׮�z?�Nl��G
�t�#���O�j��Mj�
n�*�5j�c)��F�I>�jH��~�j�����L����J{���f�ou���{;"���	46���/�j�AaݢS������(�H�����*���9���5�3KA�S	2�Ft����Y��6r�8Ae~�K`��͔�#�����-7��p� �SoB���X"�Y;]8ȯHNo�k؛���������(�7��5P;��
Ұ��Զ�~%���&��tf��=�&eg~+g���SM&�&�w�u3�>Ze98,9ڂ����l�p�����jCH0��
��1'j״�e��4f}"/��ne3?��c~J�����:U����~#Z���F��J΅m�qI��i@o�le#6�v����5Rɫ�5*�DUL枉���Qd�|OS��̅���Z�H*t�b]K�\�Y)�8��X�#�����+��ǲc�d�QvI!ЙNͭŐ��!��5�Z��������z��i*�j�C�.�-wg��~����W���0��K�TOA~"u=�΂M�n�4?;p�����>�*��A�N�絏�Çg�j��H�Q}���.��$Qvx�;p6������`#��,<�z�>u�0�ƨ�x
L�o�R�2�>��n9�������;0��Ӈ�!�6��[�A��䶜*��Dm�r�E�I[bG/jo���P\;�NF���m9I��:i���L��%�NJ�[�<�>�+ΔeJI[�Idk�*^�P�>W�Gj�� ZJD�����k�7g-��]��]��7#���M��*;hЉ�hT�_ۨ�ݐ���):�F���w>��x��|>�#V�W~b���<:��e��m�Ɛ�A횪B8{�=�
�,�+�"���V=����i���?@ň.7O����x8����(L��-�k|w1jSAO9^<�R��In��ج1[��v�T��}q�8Č��E��.0sYC��>���ݪG�8G؃ZF������tq�)�&�p
�v��~�C90�;/�
�&����%����zW/�d�\Ԋg�D۪ІҊh�݋׸]7��~�zPn�9�;/���"0;�u��X*O����P�H9К��/��>f��_�' �{���:�]y�Ur̠��ޒ�1!�[��|D�Zş=m��c͊�)z"�S*t�`0쉬Y�T�U����N$�(�Um$CH�)���GQh� �uF��l5�NA\k��Y�y��Kٱ�V<3�*Q2�JN[�*�#P��P�^�<�**�9�,�DI����Os)�I1�aWq9�� �����R4����a3^ 筢Αh,���z������zB7#�:4�ȶFl?L�?b9��� u
���h�3���V�A�&�36T�$$p��0��ؘ\T���̊��c�Ӌ ,>���$�
���2�I|xc,Ƥk3m���V��r`
�`dT�%4yӏ������#�H�/��+to�2�L�(-���"N`4����b'��nU?�1��}IO	n��c&HzJ@>�f,�!rD��j�]�9�į�����V��Y�$��>CkW�y�c�A���5��[�Z�=k�1Z��ً�_�X�>��G��GW=��pׅwu�Ta�WT�=��4�q6��J�o��_N�1 ���S�=�G��j=�>\�!��?w�C��&VϺR��Ԟ��#�i��&(��DP��YX��4�\��A �`��de���l����K.�UsoQ@��\i�ɰ�A��͆��9�~gmL�p�Q1_�̎��LeLn�nAb~;���>�
i���e��[�e�ҕ�_�!���ۺ���(����`TH82w�ް���~��LrD.��xot�,�H�����@���#���;��^D��6?��V��O
��S[E��4v�m3KIu�X���P͠��a(�n���k���R,�b{��E�кD�>
�_����D�L���f��7��ڦ}k��D;>��J1׿J����id�SՐ��\jL�1R s��:�0#�#��X��Q��.��~�܁�4,ނ����P|�H���1��?!���u�&reEa(m5V��@^O�է�X��l߷=p�OV����$(����vṕ��-���{n��zn��ǱJ����H�Y� ���r������Y�j�L�Z��g�\��� u��$
����L6��y����ĺ�AC�c^��']���B)����	��Q�	r�&is��-�)#�S���Ɵ��Ӿn�[M?�poР��Lo_n�r�}4�}�B���n�,�p�(b�ϹM9Ŀ�p�t�@OMK���'�p%�x�_�M���H[ƣ}R��+���M�ƨa��"�z�T@�}���	�V��Tϼ�xxX����l2��ϩ�~]g�d���.Ej�\J��M> ��脸���4��R+T޽�t���l�vȼ�yFno�Hj�ڥ�d����k�܄�p�go�0��E���7B�!b7����WI^���M⛀<[e\�h<<]rN�^7�"zp��fv�B���0Z����)0�aR6G�̐!0Z����0�3n"�g��v�t�W��hC�,t�V�ݥ�i�fM%��_�f�f��]g���� �7�E�f��$�#
?�(V�� L.��	@{�asj9ɬ����$^��f�ѐ6���l9}�*�g�Q��I�1�"C����7l�K��. �w�z~̡��m����u�n^����j l>M�éQ���)�_T����{�޺�w��-��TƼd6���0�@qTM�[�[+��7�A#��9�Gr��O_�~�؊���̉B"�5E���L_֡	<vB�T��StV�^E,�R}��N�Oi�.����'���2j?�!���^��Yd��٠�+ �#ο��zE�w�H�P�|��%���)���!B��k�T��a�6��p�u�dI����?S[�c��@/�����0j���!/+��z��x(2�6�KW�*���J�`'�ɻ�0�Rzf= �6=��8�gw��Y.��f�RKr']���m�Y���=�h�_/(Y�S+�]��x��8�NK 'D���m7)U�0���"�]Wаc�,�ˬ�<c�lY�e�9��p�u�G6�d�T��((�"���12��8�n�z���O7�� ��Q��n���ff��F�7F�5+�!|k�)�(�4܆��J۟�S�P���YҾc���N�ר@�������d\�257�D�a'�˖��Ju��"sM'�ꡥ��M� �\�9�{Ї\�upew�((w��h7?��	���Z��p���������Q�m�K�S#x	'�ܻ۬_���ÖГc�6��泊�Q\� �B �*O//��2U�+}T�Vd�H8��a[��U�@���O�w�?��4�k�Á�F���nOw7t��J�i	'��� (�6��6�uhM�h�85�XY��@�#kZ�:1R

�
�\(e���?Α�OGAG�Q~k���8K��|�����qT�>�o�x�UH,�	��g��J�U�G�<��,ݿ$�Sğ��/@���8+*�T���7u�Q��&Ζ������c94	E�Q����Ѡזz0�fZ��	�ṁ��#{j��F�д����y���RNx�)]���eF�&��7���M�N��i��s[�Gf��b�X��N{�#>�=b�ޘ����JXP��z�;Gr���a�t\�}�H����ķg�[�0jV,�X^n5��j�H��7�) ��r�1�Z�����bE~8z왏���Ad�L(�P�Nq���j���)�����N9�_K�T����2F���k^%*� pWv�`B�Ty���>_3I��I������l��L��R���~۞�b��"�Λ[b�ݟav����!�^���)�q��V��0�?�~"ļ ��x�գ��Bނ�X�1Ŗ	4�׃ �It���9g4KE��M��\�/z��m2�J���9���e��s44,���O�V*W�z#GO:.��m�X�yK㞧;��3�c�xt]Dw��?�����s�Tt)����ŭhx^��pw�Ч��P���D����0d�Q�-Ij�/�|�߼x�[
N���Cm
�����T���Į�������=�K)�La�¦�Щ&G3�f}���bƫ �G�3�(���	q�o#�5o[Wq�NB+�v_�vg�f�B	��1��B�9{��x��Ӭ{W��pft+�23��y�c���4���p����'����3&����(,��Q���˨��t�%��֧c,�.H��1�2d� ��7�d��%G�%E��ty��vgu�U&�*��9cG{O"F���@���8x'�YʥQ��������^B��&�c�)$څ�Y�o�7�h.Q��ުY�F#	�"��&g����.VL!r�k<�6�6y:�8q�?2~�#��v�r�p�B"��O�6���L��Q�=�_�ő��pey�G�:�[�U H��(�F�^5�5�V&�����mլF��� d��Y&��إo�k����4>J��}��x���^W\��C��Z�f~oȽ��'����q�1�^����x�(ΈQ��kgߺV^�E`�������B�	=�?�\ �6	��&�#� ��T>�����<�±���E2�<��x��mZ��4���F3��eX����n�>�A�a|�c3ag�93F���ß-�6/�Mװ@�G������]���>�˺*~p���nb�NdzJq{US����im�Q9�l���yR��gH��]�M ��8�A^%���&4�/=���0Fl�ұć72��b	S|���PB��J��,D����O�����1���&=<�()��.@P?x'�2�蛯U��M���=\C"C�c�X�V�(V��&���ԏ���0����9m������V�.���%�V�j����&���\��=�M�h�-e(,����6+�aE4*u@�ݒ �ܚ��IP�)��*��?�����G���ߙ�� ��y ���-B��FDQK����#4j�QΚ� �́�|���,]�:�a\}6�-:l''v����]a�;�e���m`y��H�+Xd�B�6���pĶ:;��ᕏ#�V�ݔ�/��,9�R�2ց{��k=j��Y4�s�yK�j��#�������a�G�6�+.?:%��O�Y�JE9x9��G�	�P��N�cTڝ�mir<4�1=r�~��Q.���T�$1���3�Ѯ��d��J�e�`�qW�m�6����)�ʍ�de�)��ۖD� c��߳o0R>W�z���5���WYy��0�Y�.��TR|x�e�hw���^��6ᓤ��(vbZL�*�e8��tJ�k��ܓ�ox��!�'�s:ҙ���3J!�w��7�������vmΦ��N5WoX���u?}M�|�|�0YUs�>�O�syQ��}Y�zw�4S��Y~�XA�s���)�V��25�l�E���$'z���M�2�fH���>ǹ"���I1��O���(AV�3f��D
���π��1�r}U����o��zҤ`��y�gd�*��R,Q1��"B�?Y�@�LmND�%��	=Ռ�7P%Ơ���mpT�xk?�~�0Y�ƴ�&2�G��l��@�/^�
��>��Kn�ʶ�<��\(���d�=������^��(W�͐0k�d��R����mU�o.{O��Ljd���_�xA�������d ��#2�s�?a��4Q�mf���N
����b���M=!�k�sD��o�����?ϸ�/P�յ�;ڀ���(y>% -�6�N9��D�6\!,|b��ZD2��Ou�! �Ӣ꺹T�������n�y1�z��?����KM�1�5�� ��ʺ�K2$>s�R�V{1̔-LL��o��pZd#
H�8G��k�ɻ\�3Y5]TY�W�=�2{��%[�]77�ۢ��{2�[��=���vhM��Ɂ's���:Gn�;_�b�f�ǿ��Af;���7�֏����t�2�F�ӂD�i�'g�!C��s��:�P����&���?f>�K����&�h��\3��e�sܭ��խͧ�Oi�,�1)#�=[�t��0�=l���vyH(<�ɬk:�^T��|s��Y������Ǥ]q����h~�-�.�5������Jڍy*F�p�!ZZ�+We�A��h,������%��2�;*җ�H��Aެ ��7h%�9��q� �'D�L0��v�{��(ة�9"��X��Ht%g��KOm�%ۃ�V@PVn�&��"���e@�R�+�W��3�&@ol���]~S��Q��&W���E�{�R�Ո�cl;"�.pp�=f���t!QM��-��ŪO��$����B�P������L+��H@�<��S>�y�I��/m}?�����
��d�A���i�sV��)�45(H�Ew^��(֒�����l����2�1�ϲ��8k!�M���hr�_��>d��|wQ<���7���Dwi��}اQU�����D|w�b�'��rc������UO-3pj:*;�� xP9�y�[rc]׊M&�J���l�Nݺ�����R
W\��OAQ@�a��ǘ2�,ܵ���E��C̾�K@�m\�㭚X��jC�g�C��zR�� �HBQ�X�(麟�c} ,�Z�'q��fB�iz�p� <�I�ʃ?���t��3��b�^�h+�h=$�M������߲�8- ��N�Y�Χ7��D����nJ��5i��j�+eI��s���R�
��1HKT�4��@:�+J���ǿ�e��sX��0�x_@�$��7!����Lˣ�n�4���z���?u�vnc\$�"�>���ie�'>���_9	!#�D�moW?���۷+�	eU���yD�u��*#^O?I�0+���샟���C�����'µN:�Jzӟ��-�Z'�!�F���o�F�)Vk�����fz�8�a\\RXd7��ńC�wu��z�����,�S�ۻÑ�DT�}ft��pMݠ�����9O j`؟��+]����J݆�4��\xF6`j�c��/AU�n�o��v�Ƿ�5�/*WS/�����bB�P쮀��9<��\���'`Ck�Re"u�a
�W��mN�� ܈�J�.��84�?�?���j�'eSl`U�,wF"�Ef�6��20j��o�Cc3[��j����Q����S�V ���PkD$,��j��!�oJc��I7�)�d ��L�0>�A�3�@���v��(_�kh,��K)ߕڄ�� �e��)յ����N��?�����ꃹ+�Vե�Cc6������I�n�<Ɇyd4ՏR�ʷm{Gb�{��ќ���lG�|���0�_�N��F��%�Px�Jt��G?�gǏ�m�n���֘��%�@��	��in�o���ȡeJ���r���GT���{���{�X���	�埮JQ�����|�y0�Il}<Y>7�o�VX���5�z��e�ʌ�.l�a�m����`�/ 'r�=�l�#� ��}%�����م/�e�_�JY���-�4��1/	"�:g�y�md���I�u���H�K'S�eyۃ}�_���fH�KN)9$��y�͂g���5��3�١˳+p�WG Ǎtn��0ã���_ϟs��,}2`ƕj�#��F��>rH�����JTr��&��F�ͫ�ӗ`��Qq&����D��A���h�*fk
WE��}O7�a��S�����s��+@3lO=��J���_e�ۚ⩢n�S��n͜ �ٔ�H��	ocb?\ �ޜ6"�t1��:����VLjn�H�7hpL����o�Z��K �3���q(S&�֧H;��p�h�ơZQ�P��lvQ�T�<>���1k��7p�6��tw����I��,� �4��fĞ_��z�j�?O�o�t�A�ߺ*���s
��Tw6|0�ٺ�(��iW��u�d�^L�tG�%���vj�� M��| ���-7@�U�I= ��o8�z��\O �����Z��؏�f���j��9P�!wm�b`��!Y}��;;�ޤZS�S�j�-B���;�p�to���ܻ��][C�����Q���C<�c�ɌubbB����p ��BQR��A#|4���������
���Q�`r�;ǯq�w�:��[Z@6T��5��0٥�z���-�č��&j���(��	A����Y��(E�N����Y�w��
Q ^�!H�<9~U�&/�������!|#G���<#B೼$v��0;?�uރ�!b��߮Ѣ		�����٬Ƅ#��EH��]�p�%2Ԝ�QF��M�_R��()���J��Ҥ8�^�TT��y�s���P�'ҫ�޹NF�.ш;��V0�z҃%i�Ge�N�z��"�+�t��Ӂ׿̑®X�ݷ"$UC��U�ɿq*/�(�}R3���:��G��������w��{c��K��YK&7���y�p^Z�2��s�\�z�b7s�تE�o��*vAZ�� ���L��$�6����Z��~���)l��uٰ̫/Y�t=��5�A|c����@��zo���/j�s$D���˲���߮���bs�)��S�8�*��l�{�%GmàR*���a:�s6ɭs�E
G��y�˹,=2@�\�RHհH� T���,��zA�VO���I^�M̉�ދ6kE�Gj�V���3�����z���~��<ڡ��m�}aj����\G7��~_�=��#�~%a�ol��"E��%��[�Wu�P���\BA�������ňv�FD�B
�J�Tqp������ h؊��&��˥@�M����_�!�y(õmv�	�NiR�L�p*�I�_���o,����1~9�q�#�d�)�ӛ��t���d_+kE}�KN��q#��ѼWK+��
�T�Ȉ�ٿ�_��)]k�_<�jwiE�\C=�ײ�l۶$���c�%�#��Z���z����kB���K-�R�K�<���P�؀�t�=uæ嗲��ч�X�ŽP��v� �#�=H<~� J�c�j`�#mZ�]y���j}�#$C��D��2E3"^2c��s��ġ$��/Z�����)�E^p5@c�c9.��;�����"�ʋ�h;��p�ɟ澠c��2L�2�:��`���t|��M��49{��P�s � ���P�r���Xi�~n�z�R1H>�h��wX���QAk�}x-U�����y�*����.�!(�o�;��6ʇ��Ҳ�d�05}������SP��b��kS4������;�y�g�=|щ+}9�oam��t8 
Q6t����ӈ��^�&C�=�B>��h6��48`�I�	��i��+����V�����L7��0�.F.A#�a0��k��-͏�l���?-<K�C�c��<�w��W�Y(����m�'�m�G�Sb�K�vw�[�L`;-�<x��$z��������q������g,ƨz�Ʈ�a�U�LQ�����t �!A�箢$mgz���Z�W�PH�?Y�s*�Z}ҁV*���jGmi�!$G�����υ_g��$g'��u���W�-[4�B����$���D���S 6��.�U �4cAy��Ht ~��P��Js_|���(��B	��G�-�����7�Kj��ܛ�SV(��p8�U��*�:����!��W��zv��h�����������Z�D�`�@�,%�m�
"�VgB�HD4~N�aMv$w��3�{k��ҩ�\�c-h�B�'��^j�J(�W�u�dH�Y�q�ɒ�O,�+Ԍ���k�D:���^���5^������vN�x�w3W`�X�kIeh��Җ� �H7ʘt+M�6�ŶY�nrSP0.��H"��F�5^�U.u���-�Y����C�ʖ�������C.�fb}]�m��xX.��{���4t�l�&�\g��t[������ә.�(O�<��k��ш�v��g������H�Db�iK�+<:��Q:�� �,M�D������c�Q��[$����b��B�<�qM�r����ZY45�/��	w�~4tt�LB�{�Y>�BH�Or��`�$�ÅZ�Q��	S��{������I���3�\���y��gc�I��8�ō�y#i�����S��k�����0G��@�~�;�D$��d�
?t�s���%5Q\�wf�)�����5�l~*��xG<�D�-Nb��v� �~X@�"g�Z�����ZQ���HQY_�oi*f&��KN0 �p�S�9���[�_��+�Dc�ģ���8$,����^�?7���0�C1�X#s��ƣ9gj>L��#2Ք�6��7�f�߇b/k��r-�Q&\��.�ߟ�F���y�f:L<����,4�i¿(�D��F���͊*��7��V;��\�&\@s����T�T{�aDX"���Rp��� �W���5�9����y������h�|@�֚���5pT���$w�og�G�,'�8߾�V�)� iί�ԉTzƈo�54c�Nh���&�$�2U����'g��Qe�@A�^�5��ޜ���Q�0}l���ݦI��z\ �I�/fr��)�@��B��di]4+�����5pZ8�$Ɯ7*����ǃ��.�uL���%�?O62��{���hrў̝�?��9��Z�Ų���R7g��>0��HLQh0V�1��k1��7�r0�\�A�s��0�˼�����x���	��J����D̬��t�����3��䧡�#ES�uT  ��p|\�
>�U�q3(�-YuC�2X�A�{�z"͋���>^9�Į���ka�� �r�����U�c��"�pˮ�1���g:�tJ��,4�ցl���Uw�d�V1d�Ѩ���qa���rF�g��u���s\��F6���i
���bZP���Q̧ G�:��32�mU�E�+�z�NJ�{)�]�{^��w��x1yl�,Y�����ҡ�=D��4*��=M�\�P���%���:ub�P�K��G�HiwY�t M5	�L4���ܾ(�/_����gB��j/�BƄ�-өK{�K�<e���^Q��:��aYz���]��AV ��>Y���o)z ���#�:͠G܍�A��V�Y�=7�O*�:^̕<CBvbى���أ������2�;��z���\q�'��}��d���J�RCq���ڰx,�s_�X��Z{���bfI��/8$]�G.8D-�<JҞ�Q�,��Q���$L���d��y��T�r@�ϙ/x�ԮM�Xd��Ogא������!��R^Ml�R�fd�� ��� �(�a�C��1�?�%^�	8�6��ѹ�gxQp��H�1K�����N'���c�؋/3�{�|���v�|�� �K &Wzj�`�k�%~������&�Mr���?V(Q��&������V���Ƃ����o�U�2�NFd�%��R@�}��G=(��|]�^il�����/=J�X���8Sz�A��v�sP����]g*�{����-ı��������|���E81r���o�)�Չ?zBn�����~p>g�B���F�t�h��4����S�
W3���V$Q5:KS�}ƅ�Lr��KΜՒl�[���T�j�����'����y*R%�\��_L�R���0b���G��	yw_���	�7*�0����M6]�A�T�uq�}�9��cM��BmRl;1�=�L�R��ۧ��G���&��@��NM�ZҀ��.jzA��P�(�ySt�O�H'JF��]"Tսw	���~�+��W�ߺe��y�Po�5�����?/܋�d���O"c4���G��7��F��Ż���"����)�`c�˩��ZxѼQ���^rV Mku2R͍�Y�̲aL'��f�l�-|��v�|[?T�e	��X�� ��=Ͽ�r8��F���
%�r`����1e��,5AT;�ki�VU8�2���bX$�⸟�D�.����R�r�_��P��n-��r��[�\(���}�z�2�-�gͪ�?�fW����肁D(Tؤ�]�(�E�9�s���.�D_V$���UDE�%��Ƶ��Tͱ�#��=7��;���2�h�?�v{��Xt �����.��~@�:��зLcm:Z��0"��r߆�h�X��衲p\�8�?��{FQi��n+8�l�_{��&jYE{��J,���r�]����!��Ү��4��6��#?���tLm�V�z�H�*xFk����G\]Ö0���:LD�=;5�p�=����g�. Ȟz��q%h�Ѫ��{�X;3��S����4��zg���Z+6887�qD�x*�K4-�s$��4�b����e�4ze `_`O4������eN⧢�
��3�y.+�֝$�[>͚���ػJ3�P�f�6����Զ������p������qB�br��ty��T�5���I�+�Z[K���u��MDL� G��x&B�NcO�Q+\��x���wr�~H
�^�>`�k;�|(�����=�U��*6��Th�KyQ�%���S�D�v"櫿��*$�N x����bY� 2K�BZ���P���v�唫j@�˅�wўL%9�P�Ũ$kML=s+��$���_i#Z���� _� ���������l�?^�&���?��5��;�ٚ��h�NtI8U ��~t�����b#�66�
Pq�9!3 k�v9+� ʿ43q�5W��d�R7-�M��qe�w>�ΐ����}��N��.�
W_�o����)Xk�2i���جX�hJ��"�j�Z6������}q���{�3���="pOp������[�B�u�IH�x&F�W�a��w~9o��Ɉg�nL�4`Tu�94+���X٨�t�
zJ}cr@Ɖ^p9�wmF]ި�J�B:�3W�G;=[�Mo!vd�6{�b1c�q��i`>wc�͡>f��_�
 X�Rj̈L:�X��d�u��ln]J�W��V�&����eƈ8я�B��zh���%���v�9���|]����dm-$��8	�У\��n��(�`:&�k<��&Ϳ�9L�9'�}i�*�!uc�5�|j,��L�5U�l�U���V�%vJ��}L6H�*F��r���<���R����*^c��u�'9�B��-A .E�U�>�D�NU[`z�쳮ߐ���_�����'����+>j�/K��̱H��\��l
}t��R5��:V)�:�z<�)�����j	/��(�2���<��Lu� �"�S���w�wB����X�c]%�M�ᐁ�H)Q��[��'�1n*A�������0`��rv6��WmR�o���[���H^�L" D��*/��Ql�4��q�~���/0S�u�\Jǀ���o��03&��M��UޢW�ޒY��jXXF������L_t_���e���g��C��D�]��E�W�,?���`w5l1�[㮮>瘯��W�b�؆�"N�u�\�X^<�b~jq����w���_?q���b*�S�]k:���z�^tf9�&z8�5�.�ǃ�����"1�F��m�1�[����"���D˼��J G���@/ "% 6�����!̒�&G��]c����eU��3y$P9�t�(��6V�#���&^����q�a܏�Mm[u��7�ϣ �i�A�Y���T�D�jב��B��l4�I�O�k2j�h��TTK|̻�Ѿ�|oa��[�s���C�ؽ8j"�-6�M�^i�h�K=cR�#���n#��SB\�̛+"�
�d�l�Q��Pҫ�c=ɞ=i��G_N�#�OK�`�,�;ɰ]K��{.�v�f��H2��p6m���M�/ S��јCN_D5'��	���0�n{7$+�V��(d��K�GuؽC�3a�m��O4�Y��d�$�{���Ŧe�D�� LTfк�\�L����"u�6�OA��#hř%�����x�d ���˖-9;	d�jD�ג!�/~��D��"�����DL�gs &C�)|,Xlz<B�v�u�w���*Ԣ�&�SE�HN���M.�h/B���tUZ��0��i�'#�>>�*�]�В@�`���w ��	)�Hf�	
lz�)vt8yl�@y�DI������+�?�ӛ#�HB|�*��)���༒�΋�IAp�.�&�c+"-K�{ך����嬙�/74�ͷ>��T��+�u���t�L�%�O�͏C��Fn������)x���f�Ev���.+
m� 2K�F���˫1[��3��aSΆS�	A)s��8h�dۈ�*���V���h�"�I�x����)�+�"9�V3-Z�WR�� ���S�d&�J�����p6g�J�߳��lE�j��Sa�S�����?�����(̟���3�Oe�q���Ȳ�I�H�]GK��Zˋdq(�Ҁ&��كљ�u�j��ٰ�q�>:R�ԅxZ�.S���+� ���a�����T��0�[L���Zms�j�<��1�q��^j]�T2� OW��?_)�!B{X� i.5��l��_hdSH���7���(S0a���3���1e���]٘K;2,�x�AT�fi�ؤ�c�o2�#��e�*F���t�w�1��8���d�	��MR;l��]4( ���_/y�e,�Ds}x��I1�Y���}��۩��y�7����	NH�\��Ǥ�_�G��iX7w��`/K8*Ty�&��2	z�P
��lwkr�~�wP��#2h�`�����Δ揚x?��!$Z���vJ�S��!�m�&ȭp���$܋�)�-%�L�A����q����,Xw� ?���mSb��x�D�\{YS���SyONQx�ZG��O'w��œH?S�@�to�3��_�>,��t�����w)m��f	��y�W`�I"�p_�[�1��$��;_1R����m���̆�>����-����^���[�e�=� ���a�e�!��YMap�X6:b��Q-����К��m��ۄ%Vz2{���f���Q=���>�	�eJ���ӕ��10�c��w��
�ފ3 �{(�ؤ��걏�"Xq�b�L�`��h��#y���}{�

	�V�,�K�0W�SY,k�������%��j�pi7p@Z6����A��!H�=q��g�8�>�cJ��D�BDO`'�`�c{G����{��e@�;�}�]^U ����<^~~7=�6�%������/0�)+o�;��Ǹ�!�^Ѝ*�^&��>gQ�VS��IN��`4%�ڹW�a��n��d��,*�����G�T�2�F���7�<3i!dCȰR���A��-�D�@�g쳇㏃���j�����K�v�Re�'~5�+�HLm��F
Ą�h;���|~�ϱQ� c��w��Y�S4TΏ�F�s����u��jڰ�sʕv�&̞��6S����`�/%f�v��-x�;���"��|���[#�Yp��:�B�>��֟�W��^P�S�&vi4��TtX1�{���=�ʳī��a1����.0�#�~)F*[��2��X��lV���D��]Пm�t]���M�;�����[j~8p�^�������cZ�f�m+���SEj,�K��P�������"�co����$��Y;Z\*4p�\� �����ݛ�w�ݳZʻY��h�Yd-b���Dߵ,�>��S1�MÓ�fT����F��<�И�	�KO�7�7��T��f��H^���5g��z]؁IP�b<|�%��4��k�f�ң�����s������/.{�T]����#E��3Ml�O���K�Pd��BC5������s��bu���B�>IM������k�s�>����Dy:��s�$��Y T5�g�x<�?��66�F��ڥS�d����հ$,M=k���]WO"(����Z(8�s���縙�+��uO�]�|�JAg'w=�}������0�i���Ԓ�>�����ϧ_�nǯC7M/5*S�mCW��2������έ���7�1�ɂ����)}���𻴃�&��c�Kv��y���?���#�L$�c�����S(/e)�m����?+�v�>Dha���df�"���2��]��B�"Q��=J P~*v��x$��¸s5ݩ$����8�E�ǧ>��mLʒ�j4�A:u�gF[���z%�W�@v]: ���S��W��t��AE���v]��Nxk#�[j�C|d�T�9�.��r��a�O��,3��W'C��Z��t��4(I0q�����V�L u��M�o����|����ҕHֿ�	į/��(e���;h�ߵ@�LJFAK�ϧţ^?�\�B�B�q4�?���	KEE�'rJ�A���*��y[�|k����D���z���\VCG�$�b�rr�4�*��Xb8�]�e�}s���m�Cw���:e��a8#�u�b&B��l �����U]����i���q�A[����|i6��Rثw�>�n�'�.,���RjD���S���N-�)pv^��?�2��QӚ_(���r�їǐ�[��o�__��˧7u�/0U�(�~:q����
��u����w�҂u�z�t�I��Ŧ���Rg=V����p�?�:��gʚ�4��Oۢ��9��F��?��NQ��/�u\/���q[U����B�B��*�`�S�����<;��V��c�a�%%c�K�'^�g;�;�<����:�`�(��;,]X�f��o�d�Ì��.ۣ�~E'.���=����K;�f����!�ws^��8��i���"*��B9k"���z�DC�q,ٮ�5�~�Ķzj�j0�?�rl�J��g"��i�?<Uϊ5�J$�zX��C�b��Ѽ�C,9�s�a�q�K�r�S�������5�LĀˏ�W(":jа�/�}E|��[����uo�Q�n���?>%�^i���סt��gt��]S���E���	��wJ)ͯ��
V6�t�����֛.[�ώȱ�ڌ�^X���?3�`�Lod�9m�ʌп�<�-���3삵�-ף�"��Y3)��>=��?@���Tt$+�'k�u)$���Gi�Tx#|'Ȃ��P���~"�&�f5�q|�����7��9�,�1�`�
�D�����1�.�+J�[,��g�ا�M�P R�?�G��w�'��#Du�04l�����0�S�TOK�������!)Nx�P��	ְarD�	���E�*;�Ŵ�t�w�@���7�K�6�7�d|��X�/��;�������oHp\�_�j�Rs��Q��FVb�b�f������f��ۢꡱ�LeF��g�5/�/���4���!J���7<Xϔ�K��!�'z�4k��T,n鿼�@�[y'J�����o\�1���x}��}������5ݷq�w-QE�=p�K{\����4����F����0p�1c�a�]�y.y�Jl0�1��������}Uyn!�b��d��c�VY�<A�wo�����"��>Mp ����f�I .@��0 zE�Fk��ȓ���M8G��H5�aQx��(d��Z�9�153��3f2W	��Z� ��%�#ej�����f��*���%������e�inV-���� �K�~��3"�Y!w��y%X5L��[�ݯ�_��R
��>�oHt�D�j�D���B3�*�a�6�&��<�N�
��a�S:�$��I���}��p����y��9F��<�&nB0��rhFSvWB;��4���'��椔&j��)=����1F���e��N���^���U#�F�Dmh���ܽf�-Lh��J�ì�Y�c֕��'�7j}�uX��	 � �W�\�7�vIV�(�_q%'w`�h*J�\�<��;r�x,!���OF(�o��HSp����0-	�:�7�o3-Չ>JS�4���XjTl&f�H;���A��9tL��{k �td����V%��3��hb`�,!4����u���FYI�m{��N[-��N�4��_מ�
�T�R���zE ۂ���k���Л{���s�H��^�3:W�X�W;�2(}}��$OW����wpz��_:�k'ܣ��O#�@NA��۳������º����,���ƫ��`>���.IW=���;��?{�Thq�4�M=�]�h[^
 f�2���9*�?��5��)��0��7(o*rW����T�F�^��G�ٝT�8"Ū��d�ݻb�R���
l�S��.G�a�b�[+�9ߟ�a�\Y��i�-�Ȣ�l̘�v�$ t3y�R�ܧW"��j�:	J��S� �a�Ig��/kR���Cs�^�����F�[����㤣v!z�9��jhh�z��Ƨ����@s��+����q)�9_t�z�΀��{����8%7�r���}`K�F�թ�3:�#��b������<�+8�6�'��wf�B�e���nYa!��6��f��\��Xw�\!�]	�"�A�~�֑��I�6�Ӓ}��<�X�׫��)�q�2�\|_�nBxx�1�ڐ6|w�-Sί^CV�d�{�||���L���9��4��f�D���.9%�ɮ5��?$����<�E��A�Gχ;���Z�������T�}��eM�v��e�3���Q����^^r��U�8&x��X�/%,8/�|��q���G�=�Q	w>w����)�q�0�-ꦰ�S+� ��/�#�҈� и�D����I1���u�}�	�W�a�V^S����j��]�!9�ֆ�\/'C2\��D���jin�y��"�&(��t��z��&H����=O����ba��!O8>`h}G�v�����V���N�=��/y��`�����sy�<����>�n8�	ͽS-*tP�W��t%.8�b���|Mѩ�����"�����|�pV�<�'�}�ɤ��QN�i��xH�6%�$H3v����#EXܒ_�f\�H`R͢�ҍ�n~BL3�6� ��m�䫊�-�I1��.�@����X��s1�ȑ;|T���#��Ș�-9��/�n*;ʛ� �t{�sJm|4�V���.��')VY�B~��w�.@��M�:�k��?�6���_����#H�!ٲl@���%�s�|:�^$��\�3���At��se�d�xhB�hO�ʻ�VB�O�xf���ö.�H�s���� |t�v\�?���{l�k��>����j�|4FXt�3ys?+�����S��(lD&�~����:\,�̘����u�/4�>���ʘ����P!�(2��p
�Ye{8�GI��D�^
y��ۀ{���&[��,�!w<+ȺǨ9R��s9$B��0aA�����=  bQ�h��7r�m�&|"N�E�\#��L�~.\ջFiuL�r%��+m��H�MB�$�x��IΜ�:�g���j��m�J���"�Xcq*S�΀�K�#���.c	��+no�=���k"Бx���T��Z78�e����-�����j�Տl|+��T��F΂iK�����㱑��1A��$����ɕ:�kkՈ7��, 2g����}�;E'���H�M��>a̓Rc*�D���E�^�9_�f2���Oca$�=������{���|M��"iO���aT+�O���ay����ua���S�P�s͵T<f��� H��S�65�Jl�"fLU Ή��bU:i`d��T_���{R N%ʎD�5�{#�R't�ꓜ��ÿ4B�q /�G�5��\�=�K- 'Pc�hOpQ���^���"h���tdK%���;�*����`����������e�����2eO�aP�ܟW|��j�J�bk���4��q�����][)cqU���О;qY.�u��E'���>�T{������p�O���5��T8�s�Y��d&z��=-��p�!1X����b��
�ښ|61�fP)	�)3��[KQ���wM--��o`�/o�:uް�/I�֥���o�w����ի��aէ�`��a�%�z�@踿T��`�Էc��P�[T��uQ�\���fMu�{�*�o}~�q6s���@�vy��;eǺˤP,׎�l���c��x.AЅ�͜�wX�0g���U�;�~���T��3l�����.�+? v���nL�sg$H�O���|`�N>Y�
��>�h<��=�9^}(�!I��q���uލ��� m�����r��&�N#��(�=�Pᣐ]7�x��s��b��"K�D*���ѻ¦}��I
r[�n�Z`��i�erΊ�z)�X�Hl'�I'�5G	��c��q����J�?�O/�5���~�V��"� &�>8w������a�׻��o��[��)g�.5�
�,&W�/��{�f��&7�?��8��X��j����&5}J)xbQ��͒�^���am�u&)�4��?S�rg��]�8qRB�fF��3���e�ݎ&�����非�h9��H�D����ĔRňb>���#(f=֧��pH8ط�&��/�����&�������B�l��M��~�ʁl�� ���!/��.��'���JP�B�pf@Ǌ����!6@��,��*��)�P��3p���@`Y�8oE��S�a������Y?;"C���N�=a�K��K�dk.-{y��J�*���(_3��I��Ϩ� �b�B�%�h�C�uh����+�n�DX!?m:If��)������?�nW�K� �� j����z�Q&�`-�>�-37��e���
n��b��������T]��}`V���r��S��`����q��pq�@R�wI��kB����*|�w���)�[PQm��'?I�Y�	Pqr�*]QJ�fW�z1q�9�дp��5�p�,���2���`�Z��d�^�5�+'jm�@�(�8����|�~aP�ܞ���A^]W1�F���<�X}pB�[8W��@��`	�wrR|�H^,�8���ey�b?4��V�l��1�ÿ<���J0է�kT�k0������=��tǭ����jv�o���������	-�j�����ڛUߚ�Ӻ8�{қr4��
��
�~��$�������#��H�oj�{��jo��GM, X�w�wq]��7�}�v�+�bc����uz��8��$5/���)G�
�6��2�0"T5��ر��N�>PX�5����1_i�/95�d��EpH��t��3�V�����������A�5������tȇ���c�~�F�*79jYo`�W}o	� ��L�?3b�����Q�o���c���^�V�0*�c�3:r�*������v�e���E&X�z�T�]wk�+>K?��)㵁gS�t��Wv2��Uڹ�[D9�F<��ѕq��=a�}p"�8*��A�"u����(<�]^!`�#׬����S��R<��~�m����y����U&�
U�K�W�� �$�{׼8@w%(�9 ���fb�a6�Y`�x����,q1a�\� <��~��#c���X^�(������%��e�5�R��������|*i)�� #��e	�r���G�/g��t�a��.����F��]�:_z���?����T@��Vqࡦd��6�����ȢY�?%�($IV�!��+�qTyzLaN�1�U��A���y�~s����R�`�`ݯ�O��]:ܻjʀ��q�X�/�ݥ�S��?���p�����A�V���k�
�8d�c��n�8.L�ca|��j�-�xgW���p�($�{��8�Oh�%`�ٱI0D�2�B�wd�O\���{N��k9�k~�tZ�/?XL1^.�9d� �s}��-}^,�Ξ#N��Ks�{&�'N��ͮs���?��r����T	��J����D��y����'w�}��H�t\��@hm=3]���ع����>Q ��+g�dt�3�J�^5z���<���4s����&W�Q*o�6�Y�:޷����%��yV���F�χ����,�����
g��U^� 7�B�::��e�s,+��M�lC��tQ[���8�n*�t��g���;M��:�;��(D�J� ��r�7㽳0Oq�j�k=HO%�w��<^�Y�Yx(H-k��)��Z��u?�țΚ�u���NB�[o�W������P')|���8���3IBN��D�0+��U3����Y�:�� jciK����!���k{�k����J%g;����ݾ�7٘�ٚ'�pv��Z:l��[$鈵�^v�s�;�
7��)M���`������cV=�*f-ظ}�ꎮ��5+B:�7�[��Q�|Y�K�p�|"X�Us��\`�C_�'�1��4�3i���~E=�>�|�Y�N�
=K,�E�ql�@��U�<(q�-xh��+-�HP�a!>��bF��ɕ���ū�}0i�O�L�tB����i��i�Z%��&,l�)�I� BS��(�e}D��t��}n�����Z�����̛��~A�!�{G/\t�b)����fk�Z��@��A�6:J�յ�F�"���6�x���Sx��
h?����V]���ܶ�������3�Bd���}ϲM2�XX�U'�Ɯ7��|�����`1_��{��4%�IojN;!�x���Xm��[��D�=��r��9/�ِ����B���s�Y�.�Ň;@�4�Q-��׿�!�!Nt�"��0��mc5|�8�N6��w�LTIB�����Lyh����=�w�w^�}0�4���pnΩ.	`��N� ��k9O ���|�y��SDLN��Iŗ$� -�Ҋ#�%��_���dɘ���;8�o�8IO����Sp���P���4�FZ;QC)R�	5�,l�!�b��ˬ�iO|�,��[���-�@�4��K�"����3�?��B�8a�_~�@U�OL�AϫiUm��%"�r�����	�rϸ� ��rW�~�s���FZ��cMݗ�	�Q�S9���q���;���|R,��/�*gls��� x���o}�u黲U�`WYV�`oj�����2j��Q�-y��I�q��$�U/���8`�+��B>�QӇ?"�c�q��[����!!S}��Sb9�Х2R�i�+(%�M���)E�J�!,����_����i=�;E��P��ʖ�J6D�A�9���S�����RT��8�X<֨�1������O:��g3y`���T����<�I�'�2���C_�bN�Rjr�	�����S$whe�&�А�\A��@ќ�7�	Jwg[9!
"�GGq����|[��eu��oqx?�_p���AO5#��5Y�-�J[��cM��f[�+�#J� =����~f�?IA����cļ�eD���Jܔ�̙G��!�2���3�4�n��HxΊ.�X��ב�A?�/�}Мr͌f��Y�-"	3�wkxdJ�5L��
}��թ�c�K��Y����ݐw�*N����sR'��w�!��L7��u��rT7��g0`�ALu3v�t���7��%���'D�X=�E�� ���nZ�_�� 9�5_�]C�u��YuU{ �u p�F�lC�<O78�!��DU�E�o�D�-�:�g�OxQ�l�]���N�G�j�c`�a�5|Ff�vTFڇ�aBΔ���87����hiC���n"ū��ו}]d�H��G�X׀;�Ɓ@�`��&��̚������{�L�lL��㵇��օ�e_�_y]5w�<�K��&�����b��E5�0�̝P���"8ا��k���
��f,?�Tlg6�A�,�ŉ�ܔol���#I}쯦�H�"/�gx�(i��J�e�ə���P�`�xZL]g_J���>C����8��/۩�zb����zKE�<��fƊ�^�����jF3n5��Iَ���)�Q���lDf�׶�R��0��LȀCy3c+��]h�{X�����"�l2AK�;��5!�!��qۥ28��~���Nz���/G���Q���{��,�����E_��"�F������L��b����YLQ�t�(m�z�7T�<l`���x$��h�J�tq<G�9����p7-�4ˌ.��Û����6�S+ت��(�V�1p�L��9?���M�H����w@-����++/��t~C� u6�X�\ĂV
���V�f=Y�z�~Ҧ֊ 6�s�%�=$��NN��S�ɲB�TO�Qb�N �`�1kuo]K"-ʷ���T��%�y�����q��M,�]�k:Ձ�|� ���&:Yn�ئ�3�2T�|7t���Λ%�qPK-�W���?Q��
4�)�x:&4��꿹0_��y$SK����k)�";_e+�2b���-��h��[�fN�����}��I��C:�7�[�_�3����*<�:	�[�� M�� �u�GQ&��8�P<��P�^-���͉��#�kXu�2O/<��c�&�rt>q���C��H�v9V\�$�?ő\��.� ��� ��ĺ�m���6-L���h)��}�?5�FJ�4tz{fҫ�B.=M�H���}�ڰ)��,F�m5l�\�� ��uJ�)��K���aćNێ�`I P�{id������������R��_�%�9�xi�M��YW�?2boZ�1
�������I�e����ď���˨�B�	o�J�9�D4Av2��&c���D2\�����Q����ð(^���[��!�_b�sn̜1lE���}ޱ4�IO{S�7(��,��?�ذ� �[m�q�>Ldԅ����k�z)Bx"E�&%W*9����Y��U��ɴ�8�Yv����`Zcr��Y�1-,�S�X��{�G�S���L}�J����r%`$=";
@!�6]��-
��s{s��C��[��Z~1���p-��k~X�qi�9��o�T����ѝ�f�k�'��3��|>�C�qR�;��2���t'y�>젏��׈V{��d�~j�g�s����L��D	<��^P��3+i�O�^{0�U��pؽG7�cq�H���$?Wϑ�K�w`.L��R!��W�%�i���IZ;�eZz�ڱ��J�8e�u(�[��(�.]��C5��a�F跍b�5�A(a�L���Ƴ76�~u�3���;Ue-&��(f��k{W���W14��L��*Etı�ɍ�j��И׷\Q�v���!�d7��I�b52��� f���k:��M�A$P 9�{��z�r�#&��Dꉃ4�s����Ǚ
z]�qUXb�,�	x{��}<�c���G���Y���Z�x�4��f�j��ǒ������#3�[I*�Mﷶ��G�c~~� ���C�3APn���j�x��_��Ngʉ9��K6Xx2�S��~�K.�(�7JĲVeU��]� ��~���ᓊ���`ŹkJ�M���'��غ
#E���_M�}�H!�ED[��ռL�����%cX��-0ױg!�B�/�ɭzԭ��OHX� 0���[T��3m��Aa�P���f�����$t��M,��ɇ�$·'�a]��ã��U~}���^!.�`s:���q+R�7���g�q]v�k\��e�chP\,��K���r���(����Zl������ρK�5N���E�:�!��!�!����/�ƌ���Y<	N+�B�.�g!�R��ɿ@�ۉv������|*pD���rl�����OO�s�z{���*v^;:�$|�,֝?Ue�Hm2K�(i���E./O�&�YA���t��Up��[?�%��,GBRʷ�ٷOMr��(��5����Ḃ��9�3����k��v��Y��l���'�@�>#nE�6�Ҕ���[��ڍ���4	��l�
�+M3#'+V���_�C�E��6s��:��[2q����5#�ݶ���{��������9`�'�2x<q��Z �މ�jEj��]�U��<�0;�(��&��r���XRY��H�<,��!��d2X�^��/x���)�ϯE׹{�rT�#9������JWɈ���}#YDE����/����o�66��N؞�ɫrj�f|qKwQh�L�*ˎ���$��/�l����C�|Xm�WJ5�0�۪���AM�� ?���A_��5����gS�*�dY{o�wN˂�9��z��R��S=!���*�~`�x�.s�@���?lۄ��=fP�KB�YY؄f��2�$N�~rZW��$o�2�j_��M���ƒ��؝�Q�I���[^��|�m�<���D�W#H����)�p�Q��k���}��1���\ �$�$�8@gv�|g�u�ُ��H�5�� >� j��<'��c���C� B�h���#�`�*�1˫{�4`�uI��{<��Zp��������O��7e���d�4sU�o8yX���������Gei�@G3�hԳ���+H��pR\�{>�@�P�y2�fj�RD	�tN}I�B��K4�n��ؔ�̸�b��u����|t�w�	@:���s*5�ڈ�� r����7]2�Z0uC�NK�y���ge�+�"��U�e2yS�$י��)M���L%�ASUCܱB�yJoZ��7�g��9p���ت8��,ٕO\�]R3A���<R[J������08�Ð4������~(s��(�򃞸��Z�N!��+ԱJX�`h�	�cҥ��l����c���g����+������6�2�*r��$�B���I�@�R�H��@4���B\�*�gF	��{�L.&ℵ G!m9�q����⁒��FeȠP�J�+ʹ�/`)�`�On��R�S�R輐a����e��]���ա��f7 �R �:ҵA��GN���R
&�Z�O�v:f��w�:�D��.�P*(�bB;Z:��C��ha��W��9C�+O���ȅ�nP֟C�Lr�$߭h�^��F�����t�����Y"�g�5��-m�>�=y`�f㥦|v<�	"�p/��0�E�n���$!�5T_%��p1���UDs���~�F�ya�k�ΐ��,�/K>���J�>���-uC���
��Br��Rէ�M��+�)�H�B��,JG՞^�!�\�[�"�r%C�(�R������	�䱚�a�,/oU�V�~���}�f|��7��H�,�~o	��30\�i���->P-w�߾5�cҧ �D4�԰��#@��\�d��K^]U7����cD,�G,���R�o=.��:'��/���F]NFr�οD��� XG=��:�����v�(M�	Ie��K�g��̵����O�g�L�+苲��&+��7n�q�HMw�ŗbd���dL4���M�daU!�= ±�Y��6�Gˬ��A�T��?ET	���/�.HՖ�Kh�AX�"�M��a�d�k۱�g��T��ć����T�n�1�;�'f�\ �mB�G�%����*�G��`��
��G�7C)F���vT;�.�S�꤆=�|�Ӎ������>�V�hSI'W)�ܡ�Q7��B�Ӂ�%�,���'o�� sܿ��B}�B�N��H�vq�hߧO���b����*������Y�hP���q�R\Kz�����99#%���{�[�`��i�1���~Hj����-�aM"<�XMv~�x"����T:-��ٵ�n��Mt���E�;�%�YPb����G�X�~M ,E֣���rlB���W/�[��3�s��ǉ�R�Jah�xN+�=�w��S�L���Jp���-���ZKҶF�do�q���ã|e��2�6���2��e�{�x�����R�<�%�t^#5���M�Ƥ�5ޖ�
�Ο�A"�ϊ��Hc������=ͱ�<���,m�9��{{鏇���0Vy��Nk�?6��e�y ����ņ�3�O��&+}-Jn� l�~�̸�8�2)F֌�ܬ6��%C�R�>��dE��͈d�o�OdH��������|�L��+�ڧ���|�s����n���+��[�ݏ\�#�p���U���c9��c6̾�����b(GJ�/��)826�d�d�1�a�V�~\��/\�����R*f�� ��V�jJц�T�:>�bӽs��)76�{j1xQ��OrO�V�q��W�(������-�Ȭ�P�3N��ʝ�c�S��ơ�εӖ��H�ir[e8�9 ���;��J8-#
R����cIW�А�&U����Z;��ࠡ~+��j_6$<�i����L��	�6�&u$�	�P�J�`MLje�(��~6��`���ڣ�#�pɧD;\r��ݸZw-�Ml��jH�����,���Y��J��k2�<��1�j�y�ď�z��w5$�7k��]�HA�0��`N�4c!Ws�&���
{�'�婢i�⹄��7ޢw8"{q����[�1�| �����t�t���J"���X�W9 �"'5�.A.���1��/�+6�}ΑHD��zcR�V_���;�( ����_{�њ�S֢H��c���Y�[z����w�j�)�>���*� Ϟ'o�, G��L'�ƩϞ<�Ͻ"��'����t+���<#�K���x�UO�*���z=�#H���ё����dB��C��-�؎��y`4<�:b�/�� f���L=��@hەfYA�W�lc�K��\�|�H1q��S�%�W+,y4Z/�z2t]�Z�έ�(^F�|r��b�b�@ٍ�B��e��3�*G�F�'��������~کd�ċ��c���6E�դ��J�x���*�������fR��Xѓk���m荭H �O�/6�:���lþ�WS�Zm�2���Z��ś�#�+�aF,�!�03��}���0]�'���9�1��ڹ/�&�}t0�']f����eW���N1nm;(��&��M��0 �"��F��8��P�j�[q��Y�ת
���|��P%�t�|#��Ju-� &��as7')�7�#�w���6H��T�17nl"�mFj�Ȅ�0�����Z����c���j0�g}cﶧ/ȫ�8��\'ˆ|B����E�7��\��U����.�U��"��F�M7�^;�F�~��d)�[�˗�L�lW��C>��/� ���Wj9�.ڻ�W	�d$h���Cfl�`�B�-�r��B�{R�6��!8= �^��!b˓]�.�ؒ�s�֊����h��@$�L���x�UF:�7x�oLx�-�-y@���JNx�3B�1zqa�]�s~����z�𺿢2J��O~�><�$q(�@y��338��-~GE�q�1��iH6�rp'��9.V,p�i�V����C�)��OARN~���7�4��wP�u�V����i���^D�6��!w`�v�;�y�� I�i��i
��C�`����� OjY�sp0O��X�r��H�<QF3��y��&R�j5t,f�Re�/c�h�� �I�D��Q-������t[�rzW��}�~�B���JP�{h�&
h��s�Pq�;_���9�Y���ъ��)��5������Y2>)���#q�~U����׆ !
�Ԅ�M���@��_)�ʉuj1OΘ��#JG�!�����8�3�X(�=\�ea1�w�'	�>���ɚui�ɇ%����p�3�/�[[���� �:���􅣤��qy Io��ep�ba�>&y���48X[��#z=˳	�'cn���d��V��՚
��T4�Z�jHQ��ɘ	�v�
 V(v�BB�#w�|�{<��:my���s�	ī�	��Zϑ��':�����P[����~���C�* M��L�4f3;CcO�jR���t7*��r���K纏�^ϖ�)��S�J'1x�2}1�Q{�zo̳��� �dd��Ѕ)3��yP��g�UI�������@tc���.���vŌ��@�g#����H�c.@�Bӗ+V_��S��ӯ��:*?s��Gu�lj�T���IW�R{/�(����� ~Vm�ąw΁���ы}�*��2��NT_��Ot�UX�A`)�.�&V�TEJ|�4��������W��C^��(�;�c��{i�z|����Z['�kϯ��dy�έ	@-�_e9�;�u��M-ߢ�טG�C�{� S5 �<z7�I�E��#§�p��R�����u+�]̌U��9�Y}+4�X.�� dC,,� �[�NHIn�����;(�U;�NG�
��d�2e�G(�vt'ǥ��#Pe��B�5`僫�%�%�P
�X� �tҲ�P�k�R�+t�b"ˍ��D��-�$��2�Z�ee�zW��a�߂[�����q�T�eg�G�X�Y�\��)�H�ЋA�eڬc���E�����2N3!��w�5y�@�)�CQl3��z�
��\X��1ţ�b[���ȍ�]��1Y/1m[�_Tg���3F�}��~���EyW��^�7�w.���S�!nx����V<UZ�a'�޴9��Q]~da4j�YY�o��s$��`��{�����R���D�t���g��9w���<���QXou��c��Bx�zs�����=,sxH�ِy��)U��L�,�ͧ����qpg��y:�����׽��B�9�_�=휗IB���t��REHB�D�R�z'n�(=���+����.�Co��Sӹ�APS����6��U�w�������)�̨֜�Y�d�WڤA�$�nt˂9��*��驝}A�Rř���ȹ����0�w��#~�%'g������^ͧ/����n��ॼEr��O9�=쌗*t4x�i˳8Fi���Z��p�d$+c_�0攐�4�i4M�4����q����Is!�B��bͧ�4�f��|�?��X<nG�{<8zȸ�i�� @X�	�	��V����	;�N'M�GA�*�z%gj�-7z��+ҩ�W���-��O��O������ZBb�O3}��($=�NS��e�9���9k�B0z�/,T��U��޽�Z�ځ�i�}d����#��7u��֢H�b6l<Jr5�����P�W6H<��&؛ˉ��u�mJ5[��>�g�w�_�!�.�ވS�P�����85�-��l�*��I��5ґ%O���?�-�kGJ�&YʽD�R �,���ZT&&gO*�q�)�<oSӝ8��\>@T�0	/U��эc'KYyLi��5�Q�[?<Hp��B�N�*�� 'Ԍ�& �,l������!p> �	1���𯑯O0����)($��=����ïR�hU742��2@o���N��H�,���Y��
=<c���%t?����ۃE��qS��^�taq����;�烨�lX��f��a�cWnI<�Y�I���� Չ�����+��KMs}����Heꠌ��1pg�� ��p
}I�o+u�@�q�HJH�Ƌ+�O��H��P)�E���=�	j���"���<q:�����$d{Ŀx�H����x �O\�X��C�zv�����N�)���Ԋc��?���.I�0���J��7�p���B� ~ ���[?����d�(b������a�b��y�O�a�
��׻�@y�F֡X&Vu��͒��I�5\�;�s~�d#�W�>�,��.d���OJ��ي�+^��c*�p��<��z?f"��$8mi����s*j7�RZSQ�.������N��/�@`�e`�ؑ8�j�����f�.1��u�^
*�Vf�>vJ��Z��Ia���n��)�W��Ҋ7�堌c���|�����o^��T�Y�<I`�G��QD�����6�.�2��?�Z��F �]�6j�Ǫ�f����N�J�Vۘ��S�y�ёxj�+P�υ*u�,~P�i��q�Qlx�"}o�G�dDp+C��;m`3=L�f��Z9n<���"�c��3�%@�ǚu5J���8#6����6^� :ޝ�s���� ���hsA���'_h�?<+~I$��I}�$@���K}��g@���#/��(���7�D����bܒ�s���c�?.&ɇ�5�!>��2��"P�Rsj�6[l�K尧b���5�G�1���Ql�WGe��#��Z�k�r�&�rB��JK7�v٘��_��Q����߿#���\��gw�+h]�ĝ2��t�ȋ��O�� [�!�ְԋ�[���1g4�F&V�ÄS2�����Zs�/��l.$�����G�޵fb'�d�~�yR��^	�pl�yz"��=ɬ=����'$�Da���7����� �Tڛ�I�H�[8���X�X���[�Eà�`2H�*e`s��pz�B>�	s���u�5�����S��o��?�	�;cw�)�<4ڎ��u�8�*���h�0�C-���`	��޻���K�v}����"��4�l����Ơ�I�v�P-@5SN� cc�Zm-6 �
�2^z����׶{�	R�-�B	�;��q��2E�(�xkK�O�_��z���BN/U6�̅KJg`�@^���l�T� ��D�58��}�������W��K���0�E�������-�fen|�
�j�@�>J	N������Ni�;i��k ǁ��4-�,���ލ�(8?w��:U�y>�� �|��>Gc�n�`�=��˧f���q���Y�!We��֤�*�8t�<nB�T$�GH{�.�,y���	Q�_�ʱ��ȓ�|}��X��6�����hu����W�ɖJü$$�9�i���J�(��fP-�W-xDU)���?R�N��Bq2�OXÐ�X^����`����`K���3��9�4��lf�=��i'�m�o"����	�x8���5 � �V���3.���������������53�M�����4���&X>�w �������F���g�N��H {�:�ScɌ*�H���ҁ��މ^���bT�E:<�%�T��Cx�C[=���B��`*��o)�"�5�W<��@�k��"�~w�i�3������uK	��
V�B�li<l�%�@������ƍ��t;Mk��U��)�҉kqH�o����0���Xb��'a��.$fv�&ܣ���0Fe(>V���?��L����J@2W	l�5Ə��]!���0K�%���@)?e���+`�.b	f$�K�k{��=G-��� ��O���U��^�?��##K�I��w/�7eu��A�s�U�\\���$���s�~"��-/�wS��Գ�r&�tl/��/r��.a_�ߧᇒ�9����R(a��;���"�����I�E.��B���P�KeZ���Fc�I�fÖ��H��~N����d��>��e�<�H���. g�-�f�RL������N�{Ȭ<�M|���z�f�����cd��7U���VP�m+Hr=c�G�E��3��N�����ڐ~+�ў���j����v��5a�L�c�!0���b؄�0� ��bs�>2�]� �L��F.4Cu��{_���� �c�d�cƐ�:����_�v��v&�N��re�)!��9Q�V����L(�%eC씢s�E'���+Ք��k�s|��O[g�*����D�v�>8�,�\��7��f�5���M$pv���%�p�����=^N�3��V�02����JP�����X������ۑPUߨ�8�������%#)t���,Q$�%�~�f��̊�֖q�-l+0�K&O�n1���rZ��?nF�L�.��g�4T�J[��b$��"�\z�P�S���{�N�9z] ���K�|�D��LIL������zw�y�}s,d.�2�5��c��8�L}�+E1]���k������Rx�`�D�ۡNUt�uo�+�O��e���.������Ǣ����� ����������$��+��,��&նl��w2+��p[y�2����)cT��y�G�q�M}6�Q�9u��Y�f2_��cV���O-ԏT@�H��jy|���ז��Wv��߬ ��[����	����9���|���_�ء?�����z�9��&Ep���1/��#j�֟���vwlz�ʔL^�S����k�����*K���B~hº)���E�W�I����˯�1��N�E	��V�ߏ��W�Ŝ]*	�E��tR�ܻh���*9mLLgc�In���%i+e0�l\Z�[���ȼ�"���&X�Y��OF�P����d�����[�ORqO��F��������Y��7�Al�����[��=� P�5����\��_�%!3@J�xr�=@�H#EQ����Xv�n�n��� f�ռ�')k�~�L��M�'GA�Q�έK�N_+��g���a*ܟ.�H{ �Mp�5��lu8�Cpe�*�h�l��g�g�2L����f��lP�0�H`�GE��%������&�Z�\�L�r�6�FW`�_�Uջ��X���jd\��`2���Y7�Lv�����᭱?[U�ǂ�\��E��B����:�t�" ��A�|Vl�[e!9r�b��'C�R��Tl�<�F�UÄH�ßFM�3A���$�##��v�q[��m�7��e�N(h�F|�{�K-��+j�5�y��̽$���O�V����u��S(��"�f?;X���E�[�`P���]	75��+a���b��
#����M����8�ДE��ό�Y�(��Q ����A��x�s��� 6��;�8[?��!�v�������6DZhw"<$���X����~A1�󟪄�2����Fh���9�3��}�R��s��r
C~�_$�L0!�y�1D��.�Ɉ#��[[���D����q?� K�VL�RXn)�[��d[��h�
b����D)v1��UZ�75���ƽ靕�|�Ue,���u��6�C�x	Ewz�4�vC����[^Zg���Y�I�x����#�v(v�>��=�hi*�Ï�c�W��4aw�����1����R&a�\���	�k(��1_ZA@�Ew���s;^�R�͵�~��!�؇�eY�Q��s`9m�B��3f�1�[�iLEX��ܮ*4���2ܟ_����V��렻�'Pd�2z6�uě��a8�1ߍ�3�j�4+������LYOfr����5��F��/?-����*΍֧��ly��P�a����GqS� �$���sp�<�iz�hb��ۚK h*,�RI�F�ʔ[�.V	d^S����8���t�5�͗�\:j����,ӝ��40�H1�p渿���j�pW��4~<�?�:����;ǭB8N**��5��x"�(��!OoFW�wRt�a�Ӱ�u����LM�(�rIOD�P�u��JDG��u���Y�v�M�9iڭ���D�U�m���ܸ`�����q����w�m���8Nb,����jsr!�}�p@��l�
U�\�BO�ԩ"�:��iLL���� aY��}C^��l��Ĝ����p+j�AJ��yQ�t��E�L�S[	���F�������2h);lX����9�~�L� ��1�2�Y���9p��zd�����G��B��EE@�.����N
>b��)�'*�V���ͻ���v�?9�h?�($�d�aP�v
7�C]Q��z!�lwLR&��������(�����ΐ�~g�a�3�d�����m��p�'o�Xk�� EFw�(��!�"-1{|,s);�z��F�����ε�%B{/��]������*d��AHw �1�N�P�����ₜdL�5N2��@��\ �����x���CC�#K���,kҝ��::/l�Ә^x���K1��/���Ė`(���� �=�h1=+5%�qڛc- v��C��e4�Xf8��E��E��xf��b,�7�@���=M�!���{o�W���L[FC8C�KnS������jJ�ZvY��Mb���5�6
�I���R���#4�x[�	?�Z%�ɽh�������!����ɑ�=4��N��#M_,����5�<>*a���X@���恿 %{��ySP�fr����9P�0F�j�I�5��Kn0���x2ػ�A/��K�aJ�Y��}x.�l}��]��vWǿ��u������ֈ�U�GUoa�׾6�01n�d=⎳3N+�	���M���8�a�e�дӭ���t���3��p�&��d��-q
s
�wi�Q��!��,��ql�(�|�^'N���Ue�R�V�G���@�G�X�A�8�1�\��4xZ���xte�����������Z��
d�ty���d�(�)��%,S���_�"2�#;�02i�O��%�tTx�aa�M�Ú� Γ�� �Q�i�o�'�
xa�zt �C|C�����h�`���
.����!Wf���u���
����mHj�L\��>��;�}J��J��C�P��H�CWh����%��EOe�ZS�֡�pf�H��@'��/��o�u����=X[~33��=$c}�x�vnQ�;�@��a�K4�$�Ƽ��	b��S�Řk���k��;@��/���;�DC��2>HG�.|�Q��<-w\��G1��8׽G/ۦ��eM??�@��cw���1�&����k�!ʩ$�I���J@��J����o�^9�p|J�\6냯{#����n,���?��(�L3uh�#nЬ�
���1�5�`��V1Qm�7���@(Մ�g@~��&�g�Ao��,�����g�aO�N��=���ʹ�.�w|�w��ֺ5b�<��
�������tLJN.�LLhs�C#��6�X�M�y��7�{�،]��̦�5SS���X3$
O0��M��!�l�̙s,xZ�Ut3��>g���vj4^"�� ��p�%��[�o��\�ձ�7��OJ���=�M��U���*��P���D���(�^�_�gq��zد����.�����v"�.8<�[^��b3� �0T�@X��>���db�1�H=�����n����':ď�Vn�[�b��M@[1�zDz�j��]�5�.^|Uu�f��8���w��`U�|�X}��Z���������_�.����vn���͟�y��eAw|�EZ1ڀ�Ğÿ��;Ch���3�B+�^�S�h�"��h��7{m��#���c��*��4�x�"�7����q�S�,~˻/�z��i�:����OM�|6
6�s�xok��J�bϢ_�L&�y�pΙ�M1 
�b||������0Y�i�k�xOm,�ߚK��d�'�џG�DK�����i['d�?N*�f�Ѹ7�乇��uU~"8ء�0+�	[�����Q8�`��֥L��b(����KH����
���з���!&�!a3#`���K�����8�֤hR��%�WT���~�}9��;��%��Y�:�x��|^���ޥ�v��h��tSD%mY��Rmir���j�+�]UJ[tz#�"�T����H�\Rl;xQ0+�>��J��shV�W��۱�Qs6qe�΂k�I�"�4��P'�x��q'nP�e3:'&G$�!)�fŠ�.)�AX�/���A
���a	 ��E��E��e�W�� ��cD�TE��+9�R�`a���R܂^�(�X�Dlb�����I��:~��rmo�,�q9�P� $��(;z��/��23���6�����Gy�N<̿�Kr�,�����>5���\���F;<:���m��Z��ԧ�Ϸ�>
�$�rx޻�ݧ*��.z�ߠ*>����&�A�U�p{�v��G%\��=1�6����q�-�s�u��a����o���TuSi1�$�gQ�	��&����Y+���اO[� 7g��4oՐ������+Pq��H.�����6@����Q�d���Hާ��������nd,�;��i�:�^��4J*���Oc4��Ҫ��Ao�7�B�bҡ�	��Q ��|�z����V�$uq�䬠�2�	.Ġ���f�GYz+-��h�b�i�Z�w��\�rM��u@G��]3$�蜍����A���&"�!M(�$^����GKp����-*�b��y�����@E}>[|�[k�KQkF��SBG�m�+B�����whܿ���
�;g�ϱ��w^��
�F�����ä�~T���t�����p�f,�k��JFI��u��Xwφ��j������w��:3vU6nj�Cs~D�q{r��Zd�N�dW�ٞ�@����4y�m�"S��u�̺��� ExHv�X�+��H�����.�.�����/� "��0ft�D�&�sQG�`��r� �[b�%��ǃ�^4/�]��d��s��L9=W�?��ӕ��y�Qh��ί�K���>ݦ�����e��OP���0�T����eQ�N��ptG$sa��QYQ��������R�`���*�z�
�"m��Ln4a"�ҡ�%�PV����lE�c�|T�4�_^���_cFg�il���5T>Ya �6E�:�;�.�/ї���{�@!�o�ʞ��A�����j��z�}ݖ'te^�O��W�եO��0�|�R4Y���P%B�{�r��8�����R݁<L<�e�ъ��pq��]I���:2�J�uʆ�%��M]($��� MX��i��0����'ko%�`8��N����)�'d�Binu-�[��2�N���\>�l��HU� ���h5�S�ٷ�8j(�0'�트�.��@\���be��q��ݬ�Si��\J�<�{���6��-�~k��A�_&�I��[����V���Q�*��u���*`����kG��=��e�ϢI�רdCW.�S7.JmnRU���]h�R8���/�FIa��E��|�%���*�Il6(���'�W�0��oy@q��!����G��&;�SC�kgCf��2͵�����W�p=��ho�.װ�2����[�t��3�E�6Z����q�3��K(?,W�ɖ���CfBc2}&�P����}�7||�v'�����H]e�l�
����S�&��"cr�SJ%�,��mO4��J�$��D�2��%��N;c �A{Y��\��8��F���R���9\y<�*�AxO+gl|���9=�d͸.��V�l��6��w��sYM��L(���/��s ٳ�:y;k�$S�	��;6	��� x*���j�4_ z��7C��8^8����\A�42Ņ�k�E��v�E#�neZ$+�"Χl�d���V��xbX�;���^eo�웄b��Ϯ̒�-��#_g,H�D�,"������%thG��C���\����?K�-�ʂ3Yx.ݛc�4B��F��Nxn@
�;yDC�z�5�7���Oi��z��Q	��5����O���O��G�v|ۯ�c��t�eG�h���Gъ*�{��YΨ�1�m3D��%�+N�[�Hw�z���=P�����롒���/�y�����g���r�,'��[dAlc ����k��p��G���F����X��Y�b�\Ќ�^�;Yr~��~l���0A���uiF���N�q�&��WFD2l�� X?@��x���G #͍7Ē[@nXGތ�7�/R4/�bc�Q4?��&�R�x<�s�6���V:� ���Qa
��aAޅg��M�k���f��k: �Q��������?�������:H'V��Q�����?;��c4��,�\l�v��Bwpv6�!x<����W�y�0���\ ��*Q�U߯�=LX��巪�8q�-|
�[˧5I���!�J�m6'�6sL���dK[-Jȏ��O�,���ex}�du[޻�KC�Y@��;Xd��+U��v �����K�������Ծ�
~�N�,߀�Ӷ��nG�s�vO��y`|�1�OB/~��F�F�hʍ��Z�6p�H{ʄwVw�ٸ0��t�9S�|���R
���酟Ǔ�#?No�n���+��O7߷d�1d>O��U׼��=Ӫ�׎ ���	\��H��?�����G2���%�-�������Ưf����?�~�`��%"����|/�~��s��[�-�e�|]+k�j�
��7�W/Z-���'�b�O�9<#����fO��w� ��:a�EoU�h�2]�0�mXSn��ж�s#!���������i�x���ѡv*.��>@CL#u����s�f铙~�["�D�e�B���@6��V}�E��Ҋ����<\p�KU������r�� ��O��K�Mhď�ۗ��V��t͓R����#X�ڦ�Xm����'>wۖbՈ��2���̘)�!S�!���l��'�b��Bz��o<X��
X����
�`�b���]��'�/˼�v�۶)��舉�q����equt4�[B�nCAȹU�pA�����+�'�xǔ��xܝ����//'��*�ڡ'"F�Ѫl/��[�rE�vO��A�/2�Zt�w�{I�%���Jß�S�hQ��(���g�qh�	{�n��[Pی`�z����j�V4�3$ĥ��:�w7��{e�tB�H�*yy��N��d	��v+�<��fO��5k�[[�O�].��s�з�w��������G���"?�z�잏̨�e<�����l��K=���S��P.�ij�@/0�\��V�Y��U	��k� �d��0��ì��37;^�d0U8�OX��<�UK�)<��~�E/Ot(�1\���h<��K��/�늓��뀚��-x.�%��n̸K�÷�\"Z���^«pDbNT`�D&M>��kv]u�EÅ�&/*�W��A�0�OaR^�I�l�[gu���l�5p���D�b�_xUS���R��f���
�C�9Rl��v"���p/������,]`��2^}��:��J7)�E�/Pe�o�8�v�mE��=}=�\����,8S"�`���	�vp��s
����ˏ��'@���B��0�{d��Gi�.9���h\�u�41�,�q"Pd���[n��|�e /O����E�GL�U<sDx����6ǣ��>��@��C�7�o{y)%圦9>^�����٪��=t�� �ܷ���)��ZQ�N��@��uX8����[e�ъ��~���^�wǠ�T�cx�Wl�5�?�'�-m���W�'Ȩ���HP7��8�ڂ�I
���\@������.pV;73]�%봻 V�:8ƭ�f���Qa�^#4���D8xQnDr��HS��}��}<m_3���K�� ��J6��7�E�ĳ�<1�E-zZ�4��b��N���TZ�?%c ���P���XU�WϦ�|�o�'�BQX������8[�٣2?^B�3�
�qgw��/���Oj��Sx:�yf+/n��K���@L(��C�63_sб���iKD�ф�+�k郜
��c(����ɢ�aLm�>Rj)M���@�įќ8Ʃ�W�E"y7�^�2�ÿ���/_emé��r�Է"���z�_�AZ�f>��β�3i0v&�����X�FnBU\� /Iz�..��?�;/�mg���S�I]����(߲�U��#z�==��W&v�����2Vx�F�����8�1�ۼy)(6�A��.)�Z��������p��ʚʤ#o���7V�R�3.�0��U�9��**ᲀ�D�����i�����%��r�ro��9���~�Ñ�b���M?T��B��sn}��X�r�a�<Ia ����h6�-���5��Q�W}'�V��|f(���>���P<�t���	�P=���[���\��)��H�e=�\X�,���e�!d/̼R�x��RƢV�5�T�(��N���Xr�+˸�����mg,����rt9(��o���.�����?9�:����*B"����rf�|�t6�.2�.B[���Mt4o�B�&T7�+IH�p�Ѻ|]�]e�t��`�T�6��=��'�Ui޶P��3M,b�i
t�z�����t����N���A޸o�ʲ��<����ra1�m)ظ�}���i��kG�q�X�oP����t�������q�~$<ʕ�07�g�O|�a�8c��}u=)�c�q(q7͝�D��
9_��m��b��xݵ��3�(y��M7F�w�'Yﰎ�~�ǧ'�h�*�9����;Q�b��Vqr�b�Pȵ�Y/�TZ79{NL�ڣy�̚�������zθ�������Vw���я>Q�S�|���~�Ϙ�)�vk���9��S�����2
f���q��<���M�����5Ֆ�&�S��$4v�!���Tb�1n� PV�*!)��G����W��/���[��r5���e�h�ue��-h��\}��)�ì�����*?����_���s���g�c� �o��?R�#5"Bc�g�S�o2������хC�5�֙?fO��ڞ-�5q�H�X}*��}�v��:������b��X�L'Vf�/YlA���Z:F׃����[�O��Ֆ��_��$lVR��y�wq�4�a��nƬcMg��|�%ȋ��ɕp����Rת���ׄ��9�t)��Y�ڈ2�-��G4a%�Jm�(�8��)RA��u,[^��b�����D��`e�tbpSS�H@a�k� �a�f�U&�Q��[��<nx-5|���#N=t���^�获lw��CҠ:��*(���[L+doz�Yj؍ ]�y����4rR�V���&��#F<��m� V8���sF�|Ĕ��S� '�z�E ��Dv|@�xW԰�K 6�3A�⭁l��|�iB>r��
���s��n�N��h' b����Ñ:�X��֏6�Zl`��ch=LZ�$���9{̯]�F�kۀ$�ԧ��秠8����o{�&�m	F1�d��2�Qh�KI��O�Q*^Ϸ��PYT���]5��6&d��)���Zi�+�,�����⛳ĳ�����xN@khrI����` �ĝR�`S��2Q{	W�P$B=\_��X�����B���Lh�#/��h���1��CsL� �)�zM���2�!q*��]'���NuV:��Tg�����q���B*�1!����q�m ���
��,L*��� "�G?���󴲲b�b,.N��7��*	y%�M@q��x��`�9����h��3�	��ȟM�K��{���� �w��׶�זi�N���K8.ִn�L��$�c�U���[���lbd�~���d���0Qq��5�:!��G�C`��g����W��T����lq��2�Hs�2�6����5@���x��(w_��߯4�`��i3X�t�V0��7������N��k�cQ�庝X��DQo�ǆXu��m��ֽ��0��C�mA�DB~��C����Mc�I��el�e`�T�dY�����"nX�w�{�`N$��7��9�;��{�+����O���4�mӏ� �%�{e�Ɍ<*��{��u^��߮�\y��"����Ow!'�L�|T4xv�W> rl�|�tB�[�b����w�n��nr�T"��b�ɘ�X��F��p�����>e�o1�L�]�OG���?�@[euqu���Z�6��\�V���%&�d�9Op��N�1�A����N��m�?p�J�|���N[��u{�)Lata�ǟ�ie�M�O3�C�"�����y��.J�hQ�iKv���Z�����k�������㿁y�q�)���:��NOaq=��CQ~�0�Pɚ%i{���	�Mm�������k�W>�8�sS*A��d�Lg�܇2]�A�|�h:�#���,�r��i!�GP�B�y�1�xE5�/DU!�9��+��o�lG�'�ݶIm�7)��W����Eq�(�$4˦!#l�+}�&w��#N~�Q�ފ��������`�7�.h�_�a��6�I+����FS8@�U%���\r���	uw*T�G5�{�s�r߶��)�nZ��,��r�c��❒�I}�G�O}���r-�	&���r�`�8DUrT�WB¯/!M���$�ab+��4�v�+�b�3]Z�.3������^Js�h��z� ��E>��]KR���Qʬ��ڜJ�b����b͟OF絀��|��<H=1tK ^�A֐S����Sc�7�٬��.��HTv���y�;����ʐ�y�8n�cD�2�p��Z��Z�)뇔!�chŽ��	��T�<]���{��D��v]_H����h�<8����u$[7s��՞�4o~��CȟYg�hFuf´KA�����(��a��uG��=��P�o�+�[��$��vO+z;����q�D-7Kb�����#J�(Jm�#V���9T�Dw�5n��P�U��<9%��I�3VQ�Z��T3�\C��2VR<)9$�bpS���?��}G�<(:MQL�wRSߠ⿆d�?�����e�U��F���>���5��&%�@�'�#��.?�9��"k:��#EkE�֪W x�Z�q�y�#o�2�����q���!�c��y�U��X7�5&��7Y�~�U������d���Q��O��;��R��.�e�7I�;H����b���5um�!*I5u�4'!��ju����X2��+?�i����)�_w�"dY^`��q��#N$4s�9��N��a�7�4I��P; q��r������܅`n�{�E<^F����w��tˬ���u1�B���>9���v��'.���b��G�޵�0C�X3���Pj8^�Ǩ9	hR��	"�r��{	����Q�:����T��Ū��.��dw-���2UF��,jf��;" �-�o{OW�|��o"���I1�C
�r���c\�.�{��}eؘ���Lڲд�!��R�\6a���6���C��x��T�-�����2&���l�x�j�����<�CC���7�I�?
�&��Ɏ������8����M	��1G�)���]�06��)�^~��LR_0m��b�+F�)����p�Q4��`!g�Vɋ��c�!�͖�hc�n�G�b�9l"d.z6�8���������<�V�z6�w	Gf-���D����M~�V%1"e�������5⃕!������R�90x���9;���ȴ�Y��MwxN��xJd�R���m2^�ᖨsP���M�h�k���< �R�<PB1���)�ϻ�$8Bh�0r��yD]��  �.b9�W�<�v�X�;Q�̉Α�n���	X��k�S�(~��� �y��5�E�	 +�����vn���Q\Ɠ�@��1�� <xm]�?*���}���}aZz+�k!n9�������E܂�U�X_��+�xǘb�l���/G�,3ۋ4|�	Z�E
���������_Pʆթ�VZ����v+��$������Ci$��:�swlGu�Q��$e�l ��z~�:�I6����f��JN�ZP^���i��pU����kz�[��d6�(}$el�/M��!@���5b�Ѻ����e�$5����:}p9��bUA4.���b�k}���F*��f_�D�=�A�W�ǂ/�>�Q����q�o�������[v�g��j���8�M7ޤ�� ��vZ�Z�	��P���@��T�����Ï4�I�U!�X�!ҕ�ޙ�7���ƶqV]֢S�p��!�����>d��el��bX�g|���i�;��ܕ5#��T=��҃�U��*�e��20��XfG=�� ���x?�N�w��-D/��v��!����և��M�`�������a��TH���x[�	��)�DQ�	��0v�/p��&(�N�4Tcu�1[�43�$9y���}�]��Ϋr��&�0yq��c��n��'qYVeb��������O�؞9w�t#W�r��76���X����J`6w� �O�sJ)�7�{q��e��[> ��/O����r�
3�2(\���S5����a(����y���` cf��n��^��c��)����5�I��>��	���~;0z��G�����)��sMr?�i�bU��ܮ��Ó9��f�J�i�Lh͂� �p�I������>�C�#�D�t}�3�1����x��Bc��ZUf��Ť:7��{�H�So_M[���y������_�=ƪDE*L���o�� ޠ�d��Z�V4a$�;?=)հ�<��ڝ�\/������a?�֖~/���'Q����,�b���N0���x��jέ$�O⑂�+��%:��\w翝����eS�^_��rT���0���{� 6M<�5v���L ��4�+f����oƙy��v>�e+���4Mk�K������t�wR�>`,�ן�-��v��;<��:�x2+����"=�>d�o�I3�szd^��:4Jwb�k/A��v�)2����'�����'s����F����z��q��&yO�����tM�y�=]�c64�2���b+�����9���u�����BP��ɦ�ȕ�k��{j��,�P�E�i_gA��b�����D�ז:<�6��9uO�So��;��6V(�ݴL̮�@�/��{�<|B��k"���b��n���N�T}���=r�' E#�4vЍG��q�?c�	:��z����gb����n���0�[�6�W��;� �5�P�E��Acn�b�g���k*y���J��ɲ�2ө%�� Z�)<��lA�������<����}��a[�ec�.ˎ5���n����p�S�����Y�{u%���V��t�	�T1�_l�r�{f;w��(��'46^�������6ʄ�����H^q{Hոp��� ����9ڦ���o�ĺ��f6 {�l:�VU#�!�����:�}a���Wtd�)}�2^���_����=����S.&�p�閔�b����hPrQD����W�Q<�Q��{1ߥ�x��AT�"�8���k���(Q=����m��*�w��kS"��؞�#�U��*���9�6YL�"���eLy�NT�9N��=<-������3�{�XA��ki�\A�1�OL����$ ?�T�� GHb�%��+��{o񗠣�K�,U􌣩��Pr�h������ϼD�Eu��4������DỤh�}*�p�/|s��kKc�R���I�H]T8�~���k��za�^~�_qm�00�%`�����|:N������'�y�8\�=B�� �ңP�¶�@AI��Kp�T3�+ćâ�l�G�\_G� 0��Ch��n�o^��l����F5\^둥�Ą�'%v
���\�r�m�aZ1�4A�R��}�����U��c�����v�����1�+r�ϔ���yÛ,�N��a< ek& ;�
��TOW����?/SWbv�0�>U�@�u��/�>IM�HZ{�"�N�oG�N��y�U�-T	�PU���q�m�� ��M;��]�� wn�	N����]Q�i��]���5��oa��j�Q�F��U	k�^�fa���~�y<�7��ym�@8��:9p �pK%���9c�Fq|�#���׺蔐�qԯ���"|��#Ja-;�+Z!�km��B],���_�$Ju��?#� ��b�W��-��W�D27����'E��>4�G|w�P���4P�Ɖg퐑�X'g�*v�^���r����J?�����W0���0��x�?z'�~�v��/R�ݥ�<����f���RۓgC1���[�G��cK�Y�_n�	+a�L}ȃ ����-LC��,)��D��̠��[`;�#�i�������1,$���m}��q��b�G����~-�qҹ����s�ш/%�9�z+0�Δ��j��h���G��mG��pk���p��wH��'Pj%��,Ȑ����m@o`�Z �ɚ�tb�qH��_L�L��)|���ZI�T>(��3��+ VG׵��Q�(	���|��*Vz���R(�t�Y��lc��I�I��ȡ�$�1I' �H��㞯5�n��[.,���_y�4s^'9�v��pA��,[�
D6�RqbۏY�^5ȧf�_x\�(�§A(�����x-�'�aMe�qi�f�2);dT�����	��H�a����Hd��c��%Y5��N�;c��&j0�^"[�u �F������U�7Ȩ��I���'�S��؁��3p�J������:����i�h�ԩ��;�-�I�E�����~Ra���K�v�'s�p
6�l�M��X�7�����:P)���cC��7����	��E����'����i>���=1�jjB�6�®]yV�(�"�h�!��p*@��7�^��Z�޶
�v(��ovX܀���ΉG����3�`�����Y���O�c���mO�#��+U���2�Em���3��q��n;$}Ir���.�(�_���"w�fpؙ�߀w ��j��voQ�0�L(+E@�OVkkr�����ol�&d�I���誠�BZ�H�AR!UUQ��=p�__���G�bϽ�)��h�r���)�o��$��w�|(��jоa��}H�{��_���m���mT[p��. y1�R.y�"x+�����@��q+ν���q����v6 l�%���/����t��ԝ5��E0B�ZS��\e�����Չ
x'��[����N�߫������-jG%O~Q��r�^��l�r�������G�H��Q+0&J��F������t�'7�KJ�y���Z����e(i=�Hmx�����z�QW���]NV����"�1qKC�2�)c1�^ד��0��&�4R<�B=�U�j�SD�&Cx�D�Ð��
d��	q�w��"kJ���y�Q��=,-#m�i#�ZȨ1�c�jM��8D�0�-�@�����]>���>������RsM�|f��
1��E����hv�����KxM��]�����(�y0�/x��z|�bW�p#B9�Ġ�2�2f�mF����8��-ٵ�\d�_�K��e����1�Щ��R<D׹��4�7�[�����S
��׺�����}0P��F���EI<-��,�J��V�4Hn��Okl�Z�K���zJ&����-u�1։6W���Z�U�nY��9�����$�n��Ml�cM�cQ�l����Rp����iO�L�eL���#C��?2r�9�����C�,�#}�� �S��X|��Ci@3.~�ʭD�C���p��%X&��ѨƎJ���l�ۖ6+�h=���䘉�	N�*T����in" 34Ƿz}��e�ܵ�|t�=Xv�SL9�@�NP%�-M���	&�NcT�v}�|Ū��eM��C��X�*}�շ��  ��.���MAU��$��ÊǸ���P_�E�C�A���(�,k4]��5�@��JL�α-�Ca� �����-��}~���'LV��c�����Z�m�٠@&�����(��Y����4��l9"��c�'ё{F2��w�.A�!���,¦R��1#.SCT��E����<B[��B�6��^l-���`U"����z�$�x�܉6M�!cӭR�B/��Z"'~P�����:�B�aݾ>o���TV	�3�1���.�� 1$�>q�dR���a)u�aK�A�lB���@i�6%j�~븮YAS�|�h�;-��14�ܷvevѝJ̳����^\b�:�a��j�P��ʻ����i	�P!e����
5��D]%���d�����E�TU���7{N�WVCQr�"Ȟ'��(�jKz��/��("VP��R�V��s��^PG��9�+7B���H��n�X�
�ovo
�������l�:
�lBf�a�<��ZK �M� �|i�6N�ӻ��'��gI�Hu��\7�ر�}���B�ްo���xA�sQ�I���,�7g��K��w�W��#ӥ</<�4,+�ϯv�)��X�@��6��ߵ��X�X��
m�3sގ�m��e�O��s*�˹������=UG��5�)�>��y���U?P�j�SOt�K"pT�J�~�v�1�d�����w��#�(�}�.�I�$ܺh��<���'��.+���.cQwRV:'��I5������V�)�N�i��ǡ����Z_���>�ޙ��d�b�|� /z雀0x����Z�x	���1��8hM>}�"����Gg��P<�_���&~~G�gm@�I�D�1�����Y|�}ϴC�	�Y����t��z�tޑ��D3�q����}��Z���x��&����v�z��n/r�֒]$�ʜ^vfR0�mL�n���v�X{dg�#?W<9GlJi�'� �K���O�R��}񗠅ӻ��05�[U�y���<y$S�
ŋes�h%����R��i��H&O��<._��q�	�����SM�N��E*<g=�G�,�xfef	Ǥƴʂ)�=̣��� 2]G�~��9ߵN��(^��/?���0	�o'��Zh�������A�����Ƶ��0@�b���&��՛��gj�GZ�-��f)�f�Z��rXlc�r�]�ͺB��8}	�ٷ�g�t�6BFV���C�cP_#Ul�L�[�>}5��Jɳ
���9G�Ӡ�qcj�LㇶԓQ�a�0(J�y��U��&�GX.���k��]$�����U��q�dQ�da7f:v�+`R�����Ҋc]E����)��4��2���z���թ�E��:�l�)i��kÑH�2g0Q��q�� �5Yy�%B5 �&����.���H��2ݰ3�j��|40�>��Ѹ�������4;�y��� =l��L6[$������}J�>�K-� �c�q�ýd�m~6�^3��ˬ5U�������I_4��)%��LK�i�N���$(�eic���ӄķ�f�&�,��A���1�������� ]D�f�v�bf4|�8lꍆh\�HBg�:���4�n�H�b]96��ܿ�B��AGV��S����C��z�)+�{:հ4ҝ����E�%�L�AR<˂�����U5��������h��7�Z9V�?�[�xW�Yַ�F��nt���mդ�/ޮ����#�˿��Ogk	y5m�>I1��}��:�W;˪a�7��;�4T@�{(�M�?�x���b�X7㕎�`�W�1���ώ[F��:2��	�����N�7;a�|ay2Ǹd�)��m"i�q��`{8}�|6~��]�7�o_���ƿ�v��^f�Q(����#���x��L��/�AQ_k�EA
����@��y���5ic�dH���T�^6�(��9����N�ƥgEd�'@�-�V��"���s�0��8���l28K�+�y�忞ݦ"�w��ԛA	�O�H��L
���#��f��W?�R��6!Zf�6��<%Md1�c�<��,���PJ�PR"�F�����L�Ҕ���3T+0	�gaZ�l�qv����sY�F��p�k��}���M�<5�+�M�b9[�L��d��փ5:��%���j�GF̬&4Ȯ=pgu�@��*��[��w8q^���l�2	ֵ���%C��|]7"Z2d�[wYk8Sv��~m� �sc���w�c|8���2��0�愊)�DN���HU��a;M=�
��n�Q��܊O�ʿ���ߩ��O�.ĮN���ؚVd^�g+����b��C����^d2?���j���[7;t�>��	�lN۔s8ƍ����HBC�̾,[q�Y��h�Z��Bz��9Z��|
���%��*Aӭ�U��fsy��x�����>HU���ܩp1��s���`|	`Ta���R�.�g�����>�E�U���f	QaL"�T3&����\�;��'�l�;�^1�um���9����"�󜲺��4�<E�(��ߧG��P��\�o��MĞ�p��[ĶxC>oǝ��RN�5�@=<'�����u�m�ۑ��[v*�_ɴ}h���׼?p�w��h4EC�1�l�.e��9�����ʴ&�z�8����zd�<�0���ES�TCIr�ޙ/�/�E����UU�F}�}��ĵ�}m�1�V����p�, R�2�b�4w���&]ʗ��!�	Ϟ�N�tw��7S�~�2UQ��U�f���Bo�>�W<IPf�M|S/>8�J`g 0�kH��nI�Tj��KLV}]?D��r�#'A�>6�mLzתr�]�Ƅ	`8.+�>��SA��\j� �,�~bDg���0Gȯ�Û���sC�$vB}�/��H�.�-�����#8}�}2��"^M.o�9���޷�I�6�t�?H�4�tA��V �`�px���{�@N���pX�>'���ALp��W��W�]q6T�6�D� �]�ٜ}4��˷�z�Y�Q�T� �?`�����g�g����@�#qJF�|��g���@��&�q�Z4�h�J8����l��=Ujbᕘ��q1���3"��H�}��*�nEժ�O�,�~�B���)��v0Au!$�Z�V��y�q��+>��%�ɗU�Ra�k���^�f��s�\(�O�aE��8���|,QO�E�q��.���bg���Bg�T�5���+��1X�:�i>�d��͆[��{�������̌�@�%��"!O;Yl.�w���G�5mE� d�����6k:�^m4��d�������m5��`p4�v�v�MEwp�9&�6��3Q�,�m��l��>����m��/���,�ߖ��v�!�������#Etn�.����뜩���
��ʏ!�q��(JC�`����p����|G_e���p���
��{f���of���I�����)9=a���W����)�F2p��˸?>Je�R�z���T �z�$�:�.?.T�"�
4Rb���_�T4�����F�����[��I�5�?��3����:H`H���a8k���}��d�>��Bh�\��pufS:ڰO�uq�ä͗%�10Q�L���C�8��f�Ĺ�qX�8�b�%�8W,	e��#AR%��6��.B�!3� ��n�:E�����V�^���3��r�t�-u�BҌ෽�XZ>�&+����녺��␏���,�;��Y��j��:���9�mֆ��`��ж ���MnPd��
�4���
�/)��$R����śgB�R��Ee������@�Dɥ��㊌�2wkǩt�d��I������ֈi����[�i)+:�bu�t�|���r����4��y���m"�2���+As��l��|q�Vl�&�De �{���u��{Nd�AQT_������K*6��	����h9��v������;�'=���؀G����u�,m�8u$G5(FN�<ݾ. �!,�I�o�hMjS1��,'��H� 5TvGD��N��a�v��K�	�W"�f�����) ��s�j!�� Q"�/@�?�)1��6��O�$e����ɷ$3�'�y���'0�4��K�N�p�����L$q�I���Y���"�T��R��K&-@>Kz}��L?���#m_,�<Z�`�(B1��N����vx#��̱�(a��+,������,��3Wv�� X�)yYRz��C��(��h3�iP�o�	x�d���ʻ	�ǝ�+RFפ�30Q��`�H�(L ���N:JE�H����Qi1b7�V#�b�`A-1�,�A_w7�A���G�/`٘{-R�=&K� #��u׺*6.�����;��x��=�$�A���y����
��û��9[7�K�{&s���V.��5�PH��@`;9�ڍP��+C6Ni�~j�7O�^D���{ �3�]hD�#����c æ��>����\r/��y����B�-�@���������8W�/"�I�hYjX�;h�7�}0 =z��ͯ}�z�,y�c�KrF6��֒]s�c.x,{φ�q�ouv[!�ٿ���"���Fd�TDǯ,!�?�Ƨ��Z�k�ć)f6�OźK��EEfUY0�Nw0�E'W��&
 �"z9�67TJSاC}YцDt����UB��d����Hv-�16W-T�?�vF�s��$�b�(6�xF�$�W����v��D%����'�G�)1�n�d�[S�q�ڍ��ݧ�]�X��c��Blr�_�o��+ak�g��O�1��G]P�j9�x�S�s��x�k�F�gJ_��N�M��ͼv��
#���N���Z~�n;<�1 �w�Y˙��|V�N�A��n��vYp���z�#�Ե"C�sM�@�;#r�eqQ{��&��q<1���#O��eGT��D�����?���� .�?8N]8!���B�=�-�û"�ع�p'{97��=0���i䌗�����v�E��pk�:��%ָ����X�J�\�lRc�b���ۨ�3s��\:�ȗ祅G���1�|:Q�9��9Ws����^vݤ#����>b�.JؔaZL����E�r&)ʱ�po�H/����K�s�e��RV�R|t�le,�i\\MY� �šT�a4劷3������UG쒗@� ���
5�ԥZe-7^"��C�2���_-���$*�I9P�d*���٬A�
5����T����a�z�
�YqRt|׷zR�J�p8��:��5����&J8�_��_'�W�jgg��Fbdu'�j� rSYhW>����o�B�'<qi�#�vM+��49�d���{ڝ�R�%1�w����^����)�\8�}�;��ȳ-@�wK�\�	����!B�a/��Č�R�;�S�t�4�<�5{���ΙӜ}>v���>	��-P���h0X�~��]Z�g>��忥��Ji�I'��/�����h!D�C?�[��S��*�:9=�"�D�j^�����a�R�i����F"Y5v������U����� :ufa����L^F�M"N��F>�I�T�L�BL�E��e�H9������/�?���\��o�ed�6���͠%Y@(xL��9�>;����[^E��A���~a9�:�w�Ė[ ������S��Y2��)Y���}�,��\���Z����).89�r�h��]�1l$��40ОB����G�˃X��#�Y`��8��56ʘq��h�$h�7`v����d<M�gB��b�k��7����v3���
W������ȴ��o�xI�@._!��<nĠW :��\�[��l���T��Ww� �/�g�Rw�#�H_�	�;R�$_������57��$�|וڹO�)�O�2y��s�"�Z
�|w"*���>|=��]�2����{�����TA��y�Gx�ǡ�r�u/ ���w�\略-�/���:+�A�Rh��e�+ ��e��h/��}�t�����o��j_�̳ܜj?��=�'��V?��<�.�tL^���5;U�;R5h��J� ��O���K�����Tw֜�K�	U�ߪv���Kb>G����:�Ę����T#�-�Ԥ4,d�m�!D�L�;�ċ0��-�=��3e���l��A�ڹ7<���KRj�0ͯ�UjL����;��Ʈ��-zx���X�������>���a�7�$���0�� !4�$��g��1�v�Q�v��:��%$ќ5�ma�����((_K��K�؄�޴�����C�m�$��ܗ��*jm�� X,��^�L'(j���7�*.խ!�Z���|c��d�ޞGU�� �t��9��9vEK7�@K�hgMX-�\	�UU�6�*�yRG��ǭ�y��84��p���'��z��ﲘ&r�:��� !mfV�$C�CL;.�ׂ	�n�99OfDrd�m�2-�x��d�����ܴ�<�5DG~M�wH����uZ�Vt��M�� ����A���6�Q�:2�w���M����A�����vE�4�L���!�J�	v�~�����!�T����\f.�^J�_2H���5���ߟ2=��o{En�!ξ� 1��]��\���XQ�!J]A��|�B��@������cL�����%� ʸf����
��oz�wL�S�>R�����d3��s�?z��'=&h?��;A�n�����U����aH5�qe+B��|(����ָ�G@"�=����VHO��^N��I�O�G�O���S��[��� *�1�K����l�Ⱦ�9Ɂs�9����[!��y"�{&1�}{�^~��7�`E�v>E��1��j̉�q`"�����Yp(*���?=��p�,�,���H�ךi�|�	m��#�c���d�k��a�]k)��NA��s�����%�E671�#b)��&�I�$����?|x�1�|��E�!pu����{�Q}�2�`48LZ|�)��(��P�����,��Ԓ��[QhS��wO���#q�G���
nL�;H�

�#y��jN,C|)�0�!��9(2ئ�η����aN���$a�cb��է�$&��KΔ/�^�Ω�'��>����*�2w;��Wa4�,i�Dm=�w�7�S���v0Y�ήP/S���~QQ-���������o�j���H��$9#N�)�u�8�H�>�߂�D���V74,ł���=�������Nl@��de�5�S%�Ă�:h&.���Q:�X��z���i���(�v�J�d%>g���DL�x0���˫9��]oɳ�J[�_MFeͱb��gc�`��{R�L�5��L�hg	*��6�{Jb�֠��8{,T�
r�˒�����<�m�Y���)��\�]�*��mX{ �IԬ���FMi�["��{3Z	�"ڦaf�(ɔrm�=�#Sz������Ec(�C�d������M^� ܂ɗ���_߮��J͛��3h�(J��1���s��=��Y(@[��L솲��v�j#b���og*6��g2�N��O�A����E�LvY¶���@�����
��+�Ǭ|�j2��*�ó4����s�؀�6c�v�84�m6��FD�Y�� ��x(�}�G��̐zE;��,EVT?=�+O��>��Uӫ^��35���9:�Ons��J�JS;�$�979��c�2t�����B@.���6Msg����tH"�XJ�x����,pJl�P�E)LGs�A��:�]j,��%�r�|���ޑ���nz `>�����K��Maa����)G�e�2C�	��"�l6/�����|;:��@ݮ`��<�`�=��Һ���3�V�V��3&����8�ho!�<p4^��z�}4�V26�>V0����hÃD�/����W�>4wT��AQ���}^̒����'i�{D��\�%��j��YD4\��W���ز��`x��'�,����q�����:<�T*%�� e#ё���	dL�O��e���Ox���U;l�`�_	x�T���ׁy�E�b.E��-]��/O~D�h˛����E���>���2�9s���S�E���%V��s�l��m�ם<��X�\>V� v:���ǗEƟ
�r\C�t�#t�q�͵߰��V��m�X�5��>�t+��� "I�w3���4�S�91X���GB�m}f+��v����m�\�޿Q"�e���L^<I�'Mg̝x��L ��wJ���ΰtޓ�P���1���@������G4
�R�j��N���LBg�LFj��il�?b���&�O��4'G���ݵ��:|�A�kv~x;+�����]o�9f7w��M�x�j���F8���ٷ��BH������p��85ڥ�_�%|Q�L����FW�;p��?�����@xM2�{�&�0۷�|����2����[>-�����k ^����T�U��X]c�hl�t�6�B=O5��%ɢ27�����`���#�M.��:�H��L�u�<ᕋ:�͔���|�q�P��w��Y�j���m�MM�\63��%��	���ׯ|\~ׄƓ���G��`�y�5#
�m�Ҫ2�I����N��>���7sE�~�9S�=��*r��s�|�[�9�R�) w1�g����dH)ڑO���.��Hg.iɎ�A����cp�ֽ��g�|N�eSn�p��C��F`(�jS���l�T�OJ��4�o�����,�0l��J�d�V�^�۔�.M��E��xGiF��J,��z.�x���b�Y�R���}�>Cyj�L��`�	oʯp��l�b��'P�_�
�=(H�|��������zc:�
k��}!��B�9q��q~b�X��.4�&�C>�a|���^�����G�QnTI�[���S�l�5?�^'�=F5F�@X�,�#�k��k�?+nxR�[8�.��ѫ�*�i�y�;�����?I.��!#ٯ���\ka���"v�ڤ� Y,{�A׬�y�A2!��~��/a�^Y���NHٴ�D฻ n3/��unK鶑�a(�E���O�#c]2���t�X_}t[����Q�	���qun��X����� �/Y��%�%O��N�Dz�~�'_É� }��A�95���8��kY�s�����fx�^�C�4�BC�=�jl� `��x<@���}�/��S{1JA��p�O��M}�@�X�su�B�G�r)X�`����rq�);~8\��5��'5�}�n�'�ѰR����⯞Ȳ:U�I�b=�q�дp���7Ǧ`�� DQ���	ulR�"k����\�؁P)!�P�g[t\ݠ��m����z8���j0��
Cʦ7�X:9L�u6s�U�T �A_����K�(
�R�
D������ ����������C���y׊����������v!;s�X
�KA��Twr��>�O6�"��m��4���H��s��Jb�lw�y"NH�M��_7l��c��bxKH��?s�U�L�SL�!~�f��o�E5/^��&���;�
����n`5E���x�+s����kT�}3��vd'N��ŏC������aW"�Q�q����VĢ�B�(���l�F��V�e�oV8!|tE�d�S��Ti�5���X=����ˁ�|��N}��� �פ�'w���*���)�D$�E�IAA��u���W񂻒Ђ���cgj�5P�j���Wg�e֠��z������.k�6B?M�o�uc9�s��<�ܾ�F�3��o��[�Y��(�j�gq:����ڃ��?���j�� �Ƒ�������sȊ3$�3҂@�%�dѵ�o>��������œf0�D��<بA���a;��6;��3�H!�]���Fv��{g��i#��u��8e5���\6G�c�4�h�*�c�OK�I�`a Ө�I�<�K��Kʧ9���Ε����IG����^��/,��xU��1�$�Q�+�M��&/{���ylF�8k�v���J����;��AtZ���SϨݽ�{��k�@&�&M$�ϩ1���qͷ�b(`N�MX��/V@��/�ɪ۔@�5�h���mN����Բh�2�}��EI@M�9�Ah3.����k�������|*1�\Ե����5��L6!�W�Yy
@�O�59׬s�P��F�h� ���:��������7iӇY�%��Yܹ�68B�Bj1R��D��z�j�y^��c�/ ��f�D�Ҋ�*���0g�c!t,=G�� �+l���˘z�3��{��p����nY.H�0i��P� ׎�}�ɀ��Op�����Gk��3v�r�t����Zk�Z9 �����쪒�	i%�K�o��g����:,U:���m|���nl�7����+�,M����o��ĭhhw�ֿ (Z�3�b 山�-5��v1�0�4L���2��}=gp�܆�J�:��;'Qͣ�f �0󏉋�aO,�œc��Q軛D.�S����I.�5s�%�p9���1�v�}�+U��:fl��jUl�m�r��L��;4ys(>F���O��sRj�V_bXY�$�6�d7|��Ҍ���������'1*7�À��ػ\�F��k=�mbf�	�zW^�m�[e�Y��g��UҐg����(��D�L��e]o���[Fo��ݪ/��Mر.��N/�7��"��U�Y$�v��������E�_�!�����u�Q�.myB'�V�N�heJ��AQҀ����9��`�������&Zрp?�k
��bբ=촍9�&T�S#�������)�i��O^��i�� [����nt:�:�H8�����
������O�[�Nt���hp��$�8�'jv�to�-�=�D+����*��I3�_��X@ZO"�3�|kfg�ќSO�1�C��j��V��� S�I9}u�h �H��X��?���Ȇ�%����	aH�ؗ�x�T�h%�|��fKon{9���c�~>A�-��f�sa��<�G<Y{�����!/3�	��ѽs8P��п��f���ҭ����3���F�uD�d4)k��Շ��)���KN{U�m��[�v�	)�.�3Rh�BY��_^"D�[!=�^�T�(B�=Fx�=�nI�u���T!���?�� 喤��Z<(Ľ׹(�;fM�)�~��J������
 �+�fz��F��b�05/�ok�A�?1�T�o�ӳ%8�IOߗ���o@,�ֿ��D�q�#��H�Z�	�9QY��#v��Q�uɤ~'����δ7���k��&Q!���b�@�P먢����k,:Q(���Ӭ<�/~^����eOqё��J]�փY�������
7+�Ӕʣ9��o�C��2l��Aτl|_ň'=}��6(���6zbA<_To��1g��T~�=�R+��論D�o���B���}�O�Ջ γ�l0i�=5صv�w�o��9�{�pv��(z9FK=+�D�u
-c[�p)TUQ�M����T�O$����*��TY��4V������F+���=Z�=	�o� �����w��+RQ��O��H���t��@�k���Uf����EH��0"�1e/F��RM'��͟F��r���FE�Xt�3�eRJ��r  Xi(a��'y��zo;����p"�]�/��q��<����*T��PN{�v� c|t��'YՀ�lf����!��V�I嵼C��H���?��nx�����d,nn��p�������+�N��*������ ���̢���l�����̤Ѳu��6�w�Ѧr�b-]���M{.����D�[�9���.�����OH�Z����\��}ʨ2K2F���Z�$����u�7͒�\؇w5�2|�C��=y���?�!K���d�w���ˤk%�e���$W�4�6B������܃	��ն���ڱU��b��3�ߺi�Vk��w��>�����v��.���Q��0�[�d-�v��k!�g'�j�l&�Dތ�a�;}cs4����Y��I�<��	oM��\�粕��7��܊�YX�h8U��04B�8��Y���G!�<o\֪9S�Io<��U.z�����$$��$��B�%�7Y;x�Be�f������ԓXr�8��C���)����ݞ�Xn8����U`��(m��R,�C����I_��ߐɠ�>�(^�Ե��C˝��Q.qD=�V�膰�N��)(�N��ӵ���"W_[ߢ�7iA5K_4:��J��쒗�`�Zx%�r�r����E�%�_H�
��%����u�6d��˯�4��M�W�N>��p�%|G�2xu�ݯ�+m�c��/fR�x2��gM�GW�F�,a�̐�͖NA�ƥ�B-���z�ר*�;����#t=X���0^eG+����G��;fM`�5V1�1����&H��uz	*�ީ�v�ʍ�����#F�a9e�=jˑV��5nw���v����͕@ C� Nε� e֠Ě�}e�wݦ��?��;�n�
�����DG:���� �\�1�����,�#{��a_?bK�o3.6T�gcЩr;\�z��b��+7d�7H	�<�/�@7���Ŕ$\��o�1V&9��y(����G_-Y
��DS�):�"Ԋm}�}�p��}ҕaI��y~Ϫ����q0 j�o<�4{�6ϵ��B�yOy����2.<���v�Yܥ{�z����r��pO��vO.X:�^�Z���WZb/w���#�dە:&;GMGDrnয�؜��"%�5WȒA]Uy6En���SŨ�s�b>e^޺h[_�N|�X�"���j3%�Bj��z�0B�P�G�������|ع����/��Tg�>�~��?]�qMe�
=�w�ڒ6,a�0��Q�幫��}��	��l0tR0�]��� ��N#p�
�tm�u��5���n��W�"���~d�R<I�.���pST�ȳ��F��"�3} ��K�T濱U���P�(�bUp�º��dDTb��)2:r! ��L����4��Tf/�MT��������[��E\F�Yo��ۆ
���Ulپ�+����{{�������M�f�g5 ���R�i�:i�-)���i��=��j�K�y\�ݜN�1l}*���%��>2Y��ex�x8�-w����Gn�1���;j9e�5��G|6��h��w�X-F�����H���4-��e�����C��-��3����?�s�%�C=B�[J&�U���hf��g�s��J��K�;P�v\dQQ���Z�y�w�������P\�_ژ�K�4��F�X�۵4:UD��a�Bd����GPz��^�úG"����v+-����Cș樬��K��+�c[���J���K�NA|�7�+������ܥ���$ƙ	�*А��r�9mxj���a��4�#{jbM�b[/�^�Oj���n��彸�j��3�3��&�=����R"��'h���`&�s��ÚhhE&b,���f�ZW?����+�؀�1�O�j��n�g#
啔�,���T��*�V�x��I k�:�`L�/��G�pRC���v��k��y�B��V)��®w�V֑PEl!y�1r\��I#I���"��T!OwM���	�ĄE�l��5S���B����R�1�^�+M�%�	��sxY� 0tR��o��2�Y��-;�zY��Pw�\�����D�_65 �^@756�C70�mT���7�3�&�K�N��d���1�8��#W���,R'2�{2W|���_��=8�D�½�*���D��1�/�AMYS���x1��5�Y1I&�*̷a��eC�7��R��U��>��60ȭ����(䳸31�_��:Z��Q1g�pf L���܇��(���B�([��L��m��0�׹�R�j)�K(�m�ߥނ�n�N�o����+��h���M�I��m��I�v�`�0��9����e��60+%y޽���8�Qҵ����~[=�=�–����6�I�N��{N�I5NG�;�c�YMD͸e#�P7�hU�tN�Z ;�u�����b�c���Q�N5�J��e����u�j����U�trx���@q�[���]�4��p�+4���~����q;�Z���[�e�pW�DL��3���q��ᜁ$�gT��8M�=�T�^��`CL����C0�K��v�%Ԧ��'��\��Ѝq>��ڲGqN�9(�Z�U�\��-8��GKQ�Y�nFsE�� ��`���[]���;ʶ�]�x�*�.���d8�𥺎S��oq;��Z�w=�Aeny��ؐ�d�.#%u��,�LR-���H�u6u����&A:��<�;7&���K��ŮCƷ�BA#`ƚ��-��V??����-�$����g���]�g�b/����Ȁ9b�"h1�z}7A�m�������Y���6�d�F��˕F�0��Z��CQJ&�u�1����z@[���fCZ�VNBwN02\ ;��f��̸�:�o���l������?�3 �Ć����*n�L���kT6#�
������+s��^l<r��vC꽿���vٳ,nN�I��E7�c�"uN���S�/�t�	C����E�7J.�!rd�PƬV[~/��!�/�{؁����Y�v"h�X ��r�A=7s��])[�Y�+Ũ-��� �M�~�A��^�5���]���ش�I@��-����%ʕ�_pP)��8҈o���Q$�#OʬL�׾V���-ĕ�g:j��R>̎�Rn�}rR�O��Sў��<'X.��h"%֠����LY{g�Qp�*L8�@�0b*��j�4���5B̥=�p/�;� �F�dh�cC-V�{';O� �o�ٲ�����C����H�퉝�d��ؿ����2�E7-o�=�1.��#�\	����vʥcj"[+���k��S��.3�j��ݪ�+S���vH����ju�0	؏e>pu�)ͱPs!2px���cb��ͼ��hW9�悶i���EV�\��Fp��d�N�g�=b�eoWۮ��=�i�s|�&�&[;(�Vl:�I
����l��Fv��'��02�v��@KL,�Ⱦv�\�ddÇ�4��G��r�b�+�c/��	��=��e3�m� ���� 1(-��ؾ����8qk�{P������v7�i{m2Z���]�ʵnG�FWf\�;��6���ܝ�y�Q�	��`�w�(��s��F�Ք�j�ŉ!9���/*�THy�����iy#�Mo�l}5�0���{���+-��g��	��p��������RL�h:�����1~��������X���F�kj!nX�f��ˡg�EiO$Y����,g,��곱 �SR�T��oq?'��-et,<�#_'b���{I���؂r�E�mP�e+�\"���ށL�مH�\�\��Rl�X�A���k$�v4]a@��BYU;�W���˜�)�2R�$M6���㜁π7;&i��T_�H��.I8yk����l� @y|��J]���$�� �|L�V��O ̍�c���E͜5�6��bs�#4�0�G�My�ԣ��TB��
bZE�P�$"!�q��4ɱ�4�\�a紈�� �ךh����������β��� �y�� �	qg�UEe]�u���T��rr�7�cҫ��P,I|9�5Y��1G���y_}�Q���-�1� =�d�"Ɛecd7��yw������*�G�jX�������/|N���3�^�Rݐ�	-i>_�l_�Wl:��\뒳#��Cڿu�b�n���P��ojk8a�5*J�{������h��g����6�tl
|�2�n���ؓ[�H���j^��mdC��m��3����0i.����Q3~��4T/�oN�[����oG�R�O�����8���P�u7Q�j�S7 �A`����zI�6~V�~ �� �I����O�T`������g��Z���I��5�ߋ&�b��-�XQ��!
I�;�(ħd���AP� ?�U�c`�3����Y���Uj����UB���c��4��:.fbE�t׍f�/�z�<�2pJ��R;����>GM��~3߷>E�����vA(�y�V�R
��Z1�c���mv?1cM��/zO�� ��Wr*�d Gc����+קQ�&��v�'�H���Nh�!|��˵$��+4�k^b��M/s���-b`(���B%� ���2�0+�gZTnjȇc��W*D��b\�=��|U��؂����{�l�ǭZ�gs����.$�ߴk|LjJ�xs�`W��oS�9?8��$��b�w��l7`$��Ϝ�A�H�,zbr��%���` �?7�x(�D�2�O��k�Qٖ���<AVu�<��T�]���ѫ�4�qI�g�����5�����_��ۍ�t�®n(�Q_�ִ=73�%h�=]v��ї�x㢉 �k�p�C��H�4y�[M�Vt��G=;G �(��w� �_<�T�d0 ��v�~-�R�I\Z��QZ� ֗�V^��`�E��r6���VSQ���T�̱Š`�4�������b�3�����:R���H�m~�~�}1�?f@D.��,����/@�� ��u0�$�����%��܌����X\^F}?���9OCs�J�ŐlP� �l~�ع�G��ƮRw*2+�I	"L�#�r�W���3��P���2&�l��_e� T~�0w�|^��zku��G<�=���.�(�Iv�
3��	.�22r4f�mɡܹ��l�Mat���w����{0\,�C-�L
6�۾}Y�`N ��3���3p�	O����,3�bk�0� �{u!|< K�􊋉�"ZRN%�����qFǘi�����U�߶8F�0Hf'�!Bg<��.�h�꟢a$"�_f.�J���Í��F�f�OH(��6Aú1��bunkك�OJQ��PHg��ְ3��&�洄	�M���FId&��&�Pb��.�q�&����rQ�>ejȴ��)��H���nte��tԦ������+_��q"�R���Bn��gᆸ�R�	��H�ZŗI����.1���1�I$n���{�k��I%3=.QL�SgE>�ԍf��(��T4|�K�.�*${E���POim<}�A��Jf/U�]�Y��RLTm^ELr��clo=l��7�G*��t��;�h��ѐx�{N�^W��6���K�if�6
�ME�Z��V�'<�2U���j��t!{�N�&A��H:��ߦƝᔸ<Kso�<QI��UN"���	F�4���m9a�8�Ht2'�(�7�fF����D�v��!��Jx,�ߣ�e�Aտ�1�{��k;9����o)57k�.ܧM4}�
��^ك�����2CxY�  k�q���E+lx/�+!�
�`Y�p�|��BՎ��1�)< yq�=?��# \H��,p^Ƶ�i��tʄ�5U|��nU�����_<��7�O(���㺲���CM=�h���Y�(�@�s=�xp/���.��L~k�۔���*��7K�9��N�v�6�¼{yUDJ-����qY�Z�����i��YK��r��Vy&�z�yK+��De��Pz��0�'��El�Oa��(���û��P%�;�ا�uX�T{_Fj_R�Fs�n\Ñ��4.��hu�zg!���)�ͨy�;�� �S��8kb��j�z��
t�DR����E��s���]!��H,�]%�����/�Ϥg��.�"��0
��%��ёm���rK�c���bO���u]|N5�x��*ً7�'�Vk�]�I�L�밈N�>l��Q_~b>f�8�<��?
��@q�똓T��K��C�f~�ǚ�VM��
J"�V�A���n���j�w~z[_'k�UÕ^�>_�����b�+�/�`vc�qlHI�Kf�Q����v��V�@��#��I�M�^����ls�wݫ!������զb�U��N�W-���1�?5�)f�-�t����YeJ�[�ɝ>U��!lş[�����뿟���0ې�7&~w�_�ڛhc[ �q�R�ʓa]M�_���q�82g�r�q�R�{�^�4P���폭<�o��_��A_��Oi���9�]Zh���Z�h+?R��e)uVm�u����e?O���3����)(�1�������U:/]�>��ـ���m�(�Kw�0��hJa!U�^K��:t�n����!g=�5-�Kߍk�k�F0����\ew�n��>LL`� �(3�jV�Iм�,��8�j����cq����z�Ru����cG�f^���;JK�H:��Jȇ�WF������J���Uq-����3Z�]�؝3>j�nW9��nG�B�-2����O?�I��mm�th�6R��/R}��s��|`G��݃�9�(` ��Ab�e�G�L��׽Au{s�R.c-Q4���A=���:��x������I�1�2������\67��
�z�C;f�ɂ����-q��E2��bq*L��J��id�)�,"�#G����xI,�^4�dh����i�xr_���Q��%CHqw�/�J��>)2�!�nD���ܢ��X���A��=���}��s�;���P�i7j�}j?�����5u.jZ!y��
��i�?��SS<�0ldXz�,�t�_���_,\��Əh�k�
��}��ܬ��{ǌ�� �s�r��	,j'j���$�AⰤ����I兇s�T���=��e�}�Y�gN��Ȍ|q+�/��gϵH�?f��:�G��i�0o�+��ҥ�V��5��R���w'�=�O`"�ק���p��}~v�|��_���f��D>I��k Q}�k�a�)�Z�Z:Q
�����|h������p��8����^�;���6kR���2k�W%�/t�����V�J}c�P��Q�`�B����Ǿ�.��y;(���8u<ѵ	�^aJ�q"(3C��/�� ��* �<?Tv>2���B��M���l���z��j���ץ<R��k�ʞ"�!�?S��x�-�!�s���p���WN��԰X��2����a��E#|o���*�&���y����|�)�B����B\�����p��k��[�	�-j��,Ft*�H`�^�$��JT�K�h��bHǇ�G����/���ƍDvDwO�\�W�R�����7�����q���;�PH���PNI��:ꥅƁ�S%iJ`jP5�<��%������٩���[���P�Z>hH�X�Z�L@Ɂ� ��G;5�&$��p)�p`2�[(#uOF��Z�'���{B%g7�_?��6��<�776����/��kG~��,�J�}���)�	�w,x������ex���� ��	$|,9M�e�
����[��`9J�r�q���8�2�������;����t&���
/z��G
������J�=�[�B7{	�����\ü��D�-U�_8�>���wu�x��p�^���a
s��zP?�!�m�"ő��"�����0^���B�O�ߕ�(����٬ۨ�y}tI���t�g�Y�N�pQ*=��ӝ�דC N�@��d��T�(�S�cwΨ��HDZ�5���L7]�,�M'�[xɸq]�K�<YG�r� `w�a����$�.�r~�;��V��e���:K��ur�"t�ote�e�Rk*;�-��%Ԥ���c'#��E ��
+ܽ(��]���^����$�S�	&\����JU�b�&��#�tI<9�A�M�9��[�'�z�ޓ����[�xH�R��<Q��-�P���H��x��l��������2�=C������v�;S��a�8�imgaB��NC��ƈ!��8�&Y����5���['���~3�k�0�g'���|�/�ub�"0��翪
�V�>��}u����[W�AC�����О^3t�GN��oi.T��xb�T$�8�Ёq������d�,P���Э��~Z� �0���ϓ� ������ �HI���R�ۀ�x�7�ԅ�b�CPz��e�{xa�\��U���
�_�O���&�6/�Ot-j��=B!oh��dw8;3:W����y���e��TZ4��c2���CD����t��=�'һ�sy!��}��U�M�b6��7���[�U]��H��7|Ӫ���&�������j��<�аr}{ HJq��o6��t��O�C���Ⴇ/��sD��ݓg3��Bb - �R8�n�P���{��I�;�[�e�����
��'�������b�;�Ϋ>��B���h��ti�PqW͑sv�c|��#��S��]�kB�ŽQ!#~ոmJ�
���+{�z����?kA�=�T�z�z8Z��I�;Y�<��FGfx ���;�ێp�K�?����s?��!���0~@��?=D���E|FO\�b�]6��\6�cy���ޚ�EmZ�-�����7��0�����Ɍ?��J3��Y���Y�\��P�U�Ga��b�"�y���r����ǚؕ0f�,�Wbg�$'�ݛ���FZ���S�| �s�ğ���+%�V�'�MZ��ץ���/��BwW���7���I�\��d{o
�z��/GP~s�3Zu����k�J�q���!Br�O�Xu$��pm~��w5�x&�e9��`K4�ɩ]R�9�#H�iJ5�*��y�f�Gi�B0�-w-	�Yd��P���|9�(�F�2*�bBL�N�(���CR����K�߭�_�F�����^�~`|�Ti2M$i�枋4R�����d��{�3�;ͩ+m�S|����tH)��iQ+�L�$����ֳ�-�zcH�αuyG撠�G/E�N�� Jގ�6�+p��ˎ���{��+2$;9�3f2���dg�Hy6�K�YO�pKJ�|�V�]�rjD���c�J�"i8���|\$�yx\<mP!�C�c�&#�Ғf��^�W�B�~9?��F��U�E+���,{hZ�3�Lʕ"p�?�l�qNAɴ�Q��S�.���ŁI�w�z���P�d��ٳ��$���:�1����Y��{VN"��6q���N\
�a��&K�15&��z�؍r�zJ���wof�H�D\+F>l��9�i��$4|	�E�´�I�_.�K�aK!�����CB�'g]�eJ�(��ZL��E@��}�/���.�F��鐙�8qنK`}�K���$��$ߴA�����	�������������+},?M⥋K�� K,�t�tq�%�jx)�@�������~�N�}x㩲�O����F��=�Ŷ�ڴ�_Dͩq����>�Kտ�+�����ݵ�E����A%���܉�
`pK_t��v� a/�o,��m�*���di�|�h��y��_˚��B8P�r��(���,����$�lU�8o!ඃ�Ľ�L��#:C%�S�]\HŅΛ�"ϲ��� ��ۀz��q��Յ8PL��.�pZ���	8��rc�fg��{�-�������[�������\qq���{ԈWV�^��T��^aW���a��i�����Ӡӌ�E3�8��s������Yk��zz�d.�`L`mX����#K��L���é�5e�Y������[c�Q���u�<��*S�;����+ԯ2$E6�R�p���k)AB�l�UU@w]y�����F�R6ң��HE��{�r�4��1[Q �8���b|��(�ǈs���3�zD�m���+S:�!8/���w`y;�~C UH>2%���`9G��#�,��_� �|t{���F�T�Mk E�Z�0:&O}�6���#�L�E)=�&)����V�l^T�V5�Y�>
��;��Y�o�
�jI�#���8u��d��o&�����;�nJ��0��3��꿨���l49��Ew���l�-t�ʣ5�����S�YQ
>)|R����fJ�g�Y�t���~��A�yaY/��ds�*:bF�$A�YhE�T�Q9��W���x9;��g��MԨ3C>:m��ms5�X�p�+ڿ�|:h��g��j��H����H�S�W�����R���l]�QL�,�J�@��k̎y8���XձG
GoUĐ+c,�r��X)mu��y�Y	>��A6>�
z�fpn�����~sv�L[���
|J
��ϵ�C"��z5���>.��={yq�:�zM�I�̾�D|!/]U��)�S���N�7��:f�o�F��v�Y�������di�Y	}o"���R��b~�!��̛�-��`�SJ�rr4��ړ��*��S����y~k��o���g�1����z	2JX=gZn`ms9��QA+��]�6%�X��Ő������f��h>�?�TY�s�B���~L�,[f/;2LDPݶgId��WG��n�O��b͒祖B���-�e�W*vjAd{��f����ĩ�D�Ihˣ��,���z�/D�v���=�!�'��M}������{�����~G,E~�gKw�Iwؽ�_���׷;��k�+?�E�hۚ��y�"�x;�c 	�ѱ�z�>�%�n㻵�1�'<k�,^F�9�p
����Q�.4���T�k�aM3C���]j��2��I&����Zi+�d�O����0(?���@������ĸ,���k�2H�����x�
	�hz�ct��^��*�Ρ�}�CDv���58���P��5j��l:��cY�U*�1M��F���	8	2lz\9�Y~��!7�MՒ���W�k�2�I�� D�Р@(��Z����L浈�=�ɜa'���0A��7}Y� �:��/F����_?���x}۞�)��П?�l=��I��ޤ�6���X�?t5��@	�EټP8�ͺ��O�]�U��ll�����ɕ� ��,�B|���MU��
*��Q�
� MDM��Lj�p9Qp�U�\X�D�-XL��R���8v�{��H����Fɤ��:U &?��h�с<���>�d�j5���6.�����HM�$?��u �+{�1B��X�g!i?Ƣ�S�l��7X|��~Ĝۉ���5L�H��J�ЀlJOг�Ρȁ	�#7��w�{5%n�Zg!�!����@��w�H���:,�2�[�wZ:u&tY�y���&��}a�D��H_��������q��՟o���:mqLE���}!�qb��������ƱG;D#,d%�QW��w*����>���S�ן|��J\[[��a/��T�	��E�^�$�CD9g�e9�uL)�F����˔6��U�v��K�VKH��5ǡ��/l�"�'��Tj��s:�`��/�6��J/z��,d���"I�8*�3j�]�D�o��6�7w�]D_/��
�l�^­���~�mM�9;c�h��Ig���@�a� i&7�5}X� W�;�T(�� Q�!�{{�i�w ��|�,�y(��y��ӣFo:
�`z���E\m�HD�ٯ�;Փ�u1Z
�z�f������N?���,X�����2�Q�K
�>*����Ga	ZЙJF;��4�l�.2��5qҹȯ�u��-�q��j��A*���F��Y?Z i�(�M���cNO9�ܑ�?��<�X��#_�Lu4��P��w+´>�!��*3�]2�H����L'sٔ��"�V#���t�o���Rc'�dG�]��LCF�c���ce +��Hq��_��V"�k�o�`�έ���U���?�k56>-��^g��G�	�}oW)\��:`\׫`{��x'�)s:,;-�M� �P��S��[8��.-�c�A��z,v�N.��>h�.�}H����w���2yL�?����Ӡo:�q���aG��غ�g�#��V�h�"���Cq漕9�ԯN�;5F�YJh�#9��Z��{3�A5Y)��7h���H�=����k��nv:�(X�q�G�<&�'9������! �V ��0
2�n&T��`�4��E�x!]ñ~���-��+=JK���� R��Df�t�[�q��������H���~[�s�``"�x��\��0K=/d��^���[�n�T�R/�G���[aX�����X�a$m�fJô��)����D<���3ծ��`,��:�x��J���1�:;\(�*l���`�A!P��m��ڞ(>�R#�	�3:9��g�&���JnR�����S~"��N[��������R �E㌚?���X�A���ۏ�6ҧ������F�5�)9�Z�2C�!��{�ȵ���d��%-uŠ�Wi*�y��)��m���z�p7"��k@b,{������MU���~]l��jHJ�ˀCk���f9ZZ���_��b>��B<����P�y����ǲ�z���qX?��V[��Mc�U�W�&~���E8�*��2�C#���OZ]��My���I�K�[��f9�8�0�����^V���ko�uW_�j[xQ��7�2�����J!�&��'�	s����+�[���b�wh��ѷ���ΰ��օ���ӹ����8Ik�
�h恖�5E���VOK��|��)�1�֢H�g����r��U 3�C��`�g�����@��2܉�#����G��Dw� �u��c�pYx,��0Q�2�p����p�@�=�#=L��ZX�~��\�~������;Q��RS���sX� ��9��'Y��?�<ODNM�Oz8s��uG���d�4���3��M,:)�}�*���gNj-@���L3$/K�gt��i#��6��C�$���0��Pw�%l_�s�>�����a2�}�lg�G�Q�>���� ����"��]p�1%��z�^
*z{}�#��O���(/�%�|dy��$�9#��3�{�@i��%��E�G]E$۴L$yp聿����:5���먧��:��o+ʌ�"ɀ�w���/�>l�b��p�;�u��4+ZL��X �X��Z��S=�J���ð%�k	��s��9~f�fe�Ɗt��s��
k͹�K�(+"��yU}�i��Du������w�9�0e�Kx�`�G�"uD���:�9E:�5�tE�T�!��`�V-�r%dx�Бq(��ْz�Z�ğ[G���MQ��@.��'��'U�L-vÔ��z���Ȉ�O�\� "tk]+*�rMi�mv�xI�D7[�?����H�L�y�Ƅ���M�pnN���Hp)P�&�m*� qRV�;��x{�)MJk��H�$�w�v�X'c2X��.>muXn� z8"�����yq@=�ś��t��Qf�:|�i�7E	!m?��@d:6�za�����X��gĄ�kO@��Iv�@�a=,cO�pK��Fb�����!�,��v|�l\;�>޶ڙe���w�2�����K
��S�M�����	�+ȓ��Z���EatH&�Ɉ�	:��Jb3G�* +�tJ�P'���bcR�m��pp�Qs���/�E�%zi4"G4���v�ֲ �'-����1s-�j	m������8ӅѹM�	y�z�p��"!姢q9h";
��K7�ѽ�ţVY<�X�\"��z9[��V*n��I���{�x�����ɜZ��ɼ�ڌ��B��-o�57��=�3zAw���,���\�~�'d�t���,5p��{ 8���������>��<�!���пo�cTC�"�����1��_�)Z��B�h6���b��[荍�N��(t}$�������!=�K���\�� B�'��9Q�;;,�j�v�xC������p��F����^|�ȡ�ɤ���K����OZ[�Λ
� �sD�/���1_���ЪW �ݼP���H�g�R�:�:�����
O@O�/���K�!4�}<;{B����ǢE�A���],��(<�<r�%ҍV���yb�m	á����Ы,��� ��Cn�3J�A��B����FF�^���%�
Q$<S'�� �č宾F$�\e�$��b��k�ae�	�eSƊHD$���0����T;p�X�&��['FX�Tm��屢���bX��N�����_"d��jLU�݄�߽����!��Y�S�Cn5����z�,���oƕ��(E]A��Z����jJ���ĸ@ھz�r�5�����N�7�Y��x�7��\��K��ǩ�*� �r�Jy�F��o�Q�tk��t��3.[��$
t�E�P�F��5T�EHS�{W�~5�.����3	���٭~oY<N$`X;�)L�L���?��QJa%���qH�O�4r�O{�ڳ�Ż��������9��::�0�LSÞ�
�~0�J��fLX�M���a���|�-({�(~!k�ݕk����̝�6���������[5r�w��/����8��é�&$u��?���fd -X��L�J���q�5�Ơ,��b{!u_�u��f&�UݮC���,Xj?�1�row�M�n�,�W	E�c�_���F�o����jI�facIi���x��/�c�>=�a�c�
�P�LFv�W��R�gr����<b&� A�\+�Ƭ,��U��"�93ƣ�RE<��<�9�n����i�:�ۧr%H��'C�
�PB+���[��-D�K����Ϸ��dI��B�RЗ���U��m�x��s^`R~�T��7�P1VAn}g�"����x�=WlFG�����k�,S�~�oD�8�Bʅ-BF��5UC|%o<t�b���P{V?�ܿ���=�zN!/I�A��Y����΅&�������\�7�J�w��1�9t�9�#�������%<$7�[k_���Қ������p6[�Z��9�[R�|2���Y�xOD/�J"h���;�����0Q�Dd��}�7�������VŜM��Y��?wLK=�)N�cMA,q7/��)����4�#T�Jw0��Bw�:�xe���l�[!y�-�Sz�y�O#�����������z��:�K�H�u��Y r��,�N7�]�
�Gp��D��$z_R<u�e�D�H`[��X�a~q�����D{�f�֭�禙��T�P7b��hX��k�}��������̴35	M_08�v��P�mYI�i�8�A7�SƳ|Ɣ�_�R��-������U>Y��97]����f0	�L�s���x����"(�-�m��ZT[���F2�M��@«�+�lm��/���g[���u�;m��Cf�z3Bғ�!�p���K+~���I�0µ:P�^$��M�-����r����Q+�kp�5�NQ��̼���"�+���#����|�����T��%NS{�o�/P/7�x?!�P��׉y��${R�=$��		��u��~�H#�?�����ڰa��*�#ɡ��u`M�L�E(��,��B�����a�4�-Af�FȒ#���:k�٣�%Ȅ�[��h,ٷ�{�R�u�������y/�%H��Y���55Z�[�}@|3�I�3��F=�Ҫo½zЧ���~M	���]� #�nn���h�*���X�$>%�<(�|؞�I�9VR�̳�x���E�=U�zY<jw�䥢?M.5[����[Q]��T����� ؽ	���a�Q�x&��[�?`�s��Қ�I��ӫy��Zx��BPT�gT~�jL��v���e��0�:�Q�晀g��kWw_���|&E�%�%{n�$�ֹ=��KG�����p֚r��f��-9�_5`PA�t�} �%��!��P�Կ��$4�����I��ޱ(���Ć'���@���5��F(��D;xi[4�SD䢳�< �77Y;�Ud���imz@��b�a�|�5:��-���a"3!�ókC���9�dsLZ����k�A<v6fZVQ$�8�;?���j&i�[t�������W���-�����+��d� s�,�ќ���'�o����$q�#�J_T���R���C��ִ6M�� j<O�bg�u)�.9P��L�>�� ��H �g�6�,/}�P�kZ���{j&'C&�(�r��u1���֐��s��@���B��Dq�R��F:�s�9�#��/��qO�
0
��`����� ���I��4������b`Wq�k(�x)lf��8���k�"��e��hD5��� �y%؄���w8X�f��(}��@D�K_-��HiR���.���3������[����������l����C�_��pv<Г��N�ӗ��L,b-����@�mc�v�9Y�+nԍ;��K����?k]�m����J%f�b{�����>V���՜ኈ�4Q���&�r�^9jqt�,���g�~(m8���g���o��R�Y���	�|�3,R��O�W���Q}���W�=�k+�y<#3��AS�}�	��������l����u�G� ���r�,�A�R/�/�	4m����t�vJO�Wa����^�ڂ���]���wo��t�4��6;�����68��T�J'n99����@&����;����Y_o���݇\��?�8F/6��>1����/hK��Er�_}ܜ�

J�"&uSA��C��{�^�`m�q�ɉ�_Ԛ�b8$a����go�ƗY�i��M�ZMu6U�����^iR�KC#�P�h���3�P�Eyf�Z� ځv�,7g��{Ѵ��|&�������{Њ���>�B�y�=�͵eD��h��y-l���5:���l��h����l�ɩ�Vs")�d�X��p>p�������1te?��B�w�5e���W�t���ۘ�T/�#b��uZ4CJ���o=�϶ģC�zyW6^|9ހg;�O�C`}�i�i0f4���2�3.�DGs�X�-��������Uk�hvx�C �����(�dD���_tz�9S>���:G{�Hڻ��X��
# �o�w���Z�W좀���~#���/��� �01�P4C�P�����6Qn3B� k��ueC��W��ht�f-�g�R�+�%'��VVG��d`�^�������]�W�\gm�",����y����J�� �s�F ���/�c��S���q����8S��y���R����F�/�]�9���0~h/썠���`�@�'���Z��=1| ���3��K�����q8�K���4`����P����\�ֲ	�Y�r��=�W�����K�'{�u��=
2���F](�j�(�,���(^q�l7����C��miQ�2r�q�ȍ^��^�]�U�5+�)U �BÑ�&g���t�n�c�#��@�A0���`������b̃�Vޫ�g�k�cF{���K��U-#Cc�5p��M���T�� �Zd�k�n	��Ƞ�Oi1�q����My�R�N������F�E����E��Ap)���yZ�-|A�Ԗj_nȖ�SDށK��tKЈc����n��?���6�١��X��w�|���c;���j��+����u0�f��j4'��q,���e��e�G|	ց��V�|��R��n2��L���ߵ��J��!(��Q�?���-�q������P���߅�Î��ZųI�AҺ@)�=�7�:����Z�ᭅ\"tj �:�����������N}g��ThOy�����$�r�^�˕
��σ[����d�R�������0rS*U��YʍC����J#�d	��:H�?Jr��~ƀ�p�1���4��[� �N���L�U���i�&����}��Z ˾ܔȶ
�~���ޛ D���_�~��8P�n��q�r��ܻ�W��p���ǻ��z�o����w���c|���bX�lŐ�0���q`��V)qT.���Ɇ[���?����PV�,�c�y)���6Ha���:�7��b�@�B��	�`Q����Rᚨ?��@�b��-�v�?!�p���w�h�dR�2:�@���)\�w�N�OfuP��g����/?��M��K �V�eT�H�����d�+R����{��6ȓ�#��"�O�o[�㛼6h�<<T���K'��~AR�����]eZ�I5vY��O]��A�&F���@�Τ�~�B�,��/�AQ�[�����3\@Fz(UR��;3����U��$��U�^נ���1��(A8tRrN�#��p���F==�A�2�؂��!Hƴ�l��f_�Y9+B��O�f�(y����\��>bi���Z��iNtu�-���9h��"R;�4�I(7֜ђg<���@V|�pЕs��tpyB o��0�t���<e�IlPb���Yw)Mz���H`��P�D���)1+�*eԫVN��(2VdK�a��@�����@Dd�l��qu79OťIަ+�My�3�gp��U��hk��T�p&�]���<�X9����9�Kl�* FuZ�;���xR��m��;\mk��w�3�|���oh0R�3<�ڠ�M��.L���S|Bp37��VW8����X��<�h@��
[u]â:������#m?b�;��6�Pط�A�������O���>�PF�@�R�8����9��:U�ku�� ���r��B�y;��*�o���X���ː��;>�B�M��\���'� �%�*��]:�iԏ1��U�P�.|6��EeaP`�ל/�F"�q#k�|��O��Pa�02u*q�n��Yx���8Ūf��R`ӟ�Íכw(��[����r�n�_�7W����O���G)x�x�6*]���ME���7��t;��^9���P�D=5]��{PÎ�� U�~8Ї�����?�y�m k
���8>}��d#E�SΙ9ȼ���pF�M`�fkt¶3�]�ZT�y�E��g�0}M����&p~��|�=��E0�́Sв�>�B�
n:��~���$4�w(��Y�z��w&;�'�|�
3яZf����\�E��Y�(�r3��͎�5�Mg6�E��-�!
.#��Z)�L��/t��f�	�����;;���]�Px�j�tD��:���z�p��f�U��-�n�r��W!�
�fȱq����Q����K��g�k��$m�R�����fІu^��d�&�:�2��T�B(����伇����m2�Dc�=��Է� ����_�嘡3���WK���k��D�z�ysѢo.}���@f����_���n¡wcڈ4�4L�홨fK� �؈бn�BN�_`�����R��:&Ԟp ����&W\7KAÂ���	�q�̖���<p�3t�$ؙM��/]��A�ϢN<d���4h�ls5//�^K�S	�O���>W��P�,B�`�}�0�);ۯM�<-h�Y���2�5�v��0�LX������=��H���w�2���T��=���;?nA�snL���t��ͪ�W��X ��~�w�,���3��/w��ח���mX�\x�"� ����̝B��sݟz�z���SϺ�T�"#i��� ��6J��7��aqP]���AD]��Y�E8��J!�;mN�-w�l�%�^�Z��U���$�R�xL?v�����;0�B�x�S��R�Z�_e5e2�8kJ�
��{G�o|�4׻ e @{]�?�#������ؿ��2���<he����}\Q;'lB��5��{a-d���Y3��J��Mg))"ݍO�U��J�N9�Ж�6V4�
��(܏$)�[�Q/~?�!��-�Y��H�*(d��@0�U���Z4}&T[�ɵ�ד����r����ˤ�S����R�)c�llzj��1R��3��«v�UW���wr��7A*UN%��q��L%���}��$c䇢V��YoEl��K��_��^�D�o؞�Y1����hAk������vA��ܚ�k�zo���>�c�q�S����~��Ӧ'�s�R�~�p�,����à`qh�qíc(�{�F��iDH׿e��D��C���;Z_T�K��o�T�����R�*�7��q�Iΐj����]fFx
��NjY<���w��I2���Io`~�D2Et���B��r���S�E���ICѽڏgp�\4�0��9RÜ|e2ae��qX:��[r�-9�y�0�����Ŋ�wqd�ɹQ�İ��@�[-t�}�楙њ���B���?��`������6fD��j���7�E�m�`�(OU0��8��W�J���F�؊��vn�c%64c�W ̖#�#�}���;Xn���{4��&�r'>��ni���<Ҟ��>�~���)g�%`����d�#��'�3t�Lt�zfr>��OkqΟ���xv"�>�Fb�����O�61���}�'}̃�m=p'?�%�E�q�D���2K��[!�U�?_�+4c�������]�yOقڑd�� mӮ9�MF	�q?E�E	H����`��LeYU�e:�ҡ,�D_h&0�<Fю�I��b�5,51J�H�x�F�o��y�Y턕w�*�2�S���}[������QW��[Yiv�Mb�;3L&պ���~�l��W5�������^�5vo�����)��v�.g��]Չ�Ŭ��}�X���sO�yz%��;�㚾*G0�LI���m���}}�jPƷ ����4$,�D_����m���ւ�{��1����чH��?+K�\D�x�=L��zo�l(��h;2����8�D�'����7Mױ[��z}ց^dk���
�S�J+ ң�p�ļ:����'���cU�8��g�Q1oE!鴌oj����c-mX0���%<����m�*�ԓn�&7o�NR�ճa�	B�݋6V�X&Oe�R�ɴ��W[;���6�&A	ڳR�S�މ���j?:l��X�V��jS�Yj2L�Zۭ`�қ����iF,��"�[C=����~yO!-����ba��-�V�m6r1DR���X}cz�Xi�E2"]����_�k�iB|Y�]��b����]�{=.��|Oۋ�I5P�g*�E2Azb�YOKg��� �� �DIWr�n3����SL/�b�u��*���+x����8*{ �:/��&}sH��f�_��o&��H�}��'�Xq� )?� l��2�~4m�]2LKjejN�un8�D�:XaƐ�+.�N{�����bO�\�Z\�m�T�XsL�V��Qr���/�;"�1 �V� pO����ςW%�w2
��b�M�G�e�詊{1�s@UsGj��~��]�`{Ct��笄%���]$2�w��^��\n�w�%:���{~L"᪡�x�S�j����5����'���~���E�{(�+a��l�Y�`xn����k>J9�9NN��YJ�r��:�-$R 닎�����o��L᪎X��ي���d��J��@*�������3�M�p�S�䢻���V�o��SvU��f�/��f�D�;l�����V�x��gCCW��L�a��ms�9��r�XF���#�FW���h�ؘ!(c��8NÚt�HGg�"&/��[��6�"�Ek�t�Tnwà7UZ+�̜Sԑ���;&����^�q�h�g, �=�%!I��5hhd��V�u��]KA��hx۸k���xX�0���/�.q���.���`�8@S~���fθC,��H�UG��1�~N"��6�]KH�L�m��2龮�� n����xO�ĹL3����
߄�c�s[	T�����������W��T�,;[e� D��Y����Lqk ���&ͧ�P��rB軐\�>�s(3K����*S=�Or�5�
5́)m&��S�z�m�RP�v�4�Dc��7)�Q%�t`f�ɸ��W��F��k��!��h�9j=S�8}��\ i3���j�K�l���yi��鬫Z;�E��uJ�|���䤠YmH��[��Gw��$���.Y��>�|�f澥u����^C��;�]���@��s"SA���cO�C�NM��Ρ~q��`�wpOY����Wx<��N�k��օ�U$̜�mx�k�e�(���i����/X|��]G�Aנ�ڠ��l�����)�#J�� �M�d��=� ˄-ޢ]%��)<��2�}���e����D%�ie����Ü�|8 �跦��4d���נXYJ_�h��DJUX{��N�/��H�u�e���?p��ok�.XF2Z����xU�)I� �DH�r���bF$I-x���)�41��C߼�e�F�ϦrpKMYe~�BF�_._��I��9+O{#W��9\�S*1�U��,q�I�����-�uR���{�����Sc�p��>i��'�}Y[�FR>j���/8�`j9���D�y�@�@���6C�E��96�|*����Fo�րH�����L��'�-m�����)��� W6�C�x��1�lS��ґ�e�B��F�r�����۟xGn�8;W��w�����V.`���� ��S
���1**�ޖH�Z�t��C3&7�</�3�q��/�p�='�������`GN�f�%{�]�Rs��8"SӴsHO����&������AYR��8q4U�W��|���!��
�ڈ��Á��+7�kX-qB"%�1@��<����-8z�����č�ź�m�{R���g����E:�g������5q3�#��J|6��j3�)�pRaG��2v	=rx;�5�rǺ���b���};��j����9��ŗ��/,�E��>�rz)�_�*4� A2�&��S�ܿ�U�a}��b��Xl�%@q�Aw�_:ET�+�+'�[��8�i�;C\��4CW��	��`L�G��$5򼤐<�Zokro[f�zͨfT��s]HWqį�'1�h�읝��Ӑ�u�º��4]�QK�3��Qs���qT�x!PT8M41�@�����ӿ����r	�v�>�������ǵ�g��%+�|YH,z	P5���N���c�q�S�C=�^Tf鈝G�,-��>�v<��
-i)�ނy�"|�psT[����I8��`oܖ#�!I犗�����5���6kP��&�u&X���O���x�z������j&WpO�nH����� ����O\P���r�5�;U`i�v%�c�'�8�h��jˉV�=��F��U�e/��}������xL�_���צ��G���5&Ũcj�7D\,Hf��i���k���Z%�W%�қ��I"���h\8ٌ׌g�I�j�0p���V��5<�kD�p�y�SR�i�ߙqhf	�>�!g~��ʞ>��b����6 _�5����zU�&V7S�/]4q�mG��)�x��C�l8��7%#Z�e��-��`����R����%.r�x�R:DL�7u�.0Ds촣.��q$p�S�h����.[H�� o��Mx�A�K#�j��G=��E����ݹ�����?;� Z��³AC�T~��9�~�/��}\NSt{�r���A&;�
����qCf��S�"���0=I��)��@�Y�m�ȋ@��
�%�(/�-�lK�^��`��=��#��0k�Z������&�L�q�_���
=ļU��J�>!$}�,�x3�������Y�;��w��3�3���g�8a�� m?T�}uڔ��L�vs1ԡǛ����Usw>�"�q%���ng��B�qnw�`iW���Q�����o Q�frM9�4;��lg�x�luq��G��S�Y���E?˩�DyO����7�G��&,L'p�u�S`Pi\e������K�ث���-G�5����2���m��F�z�����F��KѲ��H��Z�A�Oi������@�rKrhcn�� �Ӗ���"$�G
��u��˃�*6�E_OYgC����JPX>�$M�<�r�ZZ4��;��Y��Φ��/�/�꾴�6���(�/��0�*r�u���2���%ǒj���i+G�%:�j�+��,�b�j��!��Ig3V�	�t�o����:��o`�.�'�ZrI�cX�6s4�8l�T�9��|y�_Ε����2�P�]��G�z�}�d�c���6g
�_��<��u�N~�~��F�q�#��Q���E�I���`GVy߫�	�ty�,S�� ���y��|n4���g�)�����NO�&e��W�.������/Hj#�KӮ�Ŝ�Z6�|�����Z��(̶�[Ƙ���6e��+fٮ���&�I��*>L�J���2��;<O�)��e��P��z�+o8�����Q��O���Ŕז���X��k�q��}N;��WZ�k⸌P�0������$�<0ND|�����5����	T��<>�n1㒻��������%NSМ<�̖����U�?]�sd�*� ������ݼ���U\ҷm�wUxSm~��!OǑ�t��M����!*��a��nH�n�=%~���(, �Ho��Pg��t�؈�M���i�e�%�&D��	i�<� ���C8�}��d)�OTɇ����A�n��Wg�T>���׋�^ZH�{7�M|�2��=�h��{뿊��zg�+~���d�'+9>-���Z���ͪ��ƴ�	���]�`���+p2s��1Q-y� ]}�n�Y���m���H��Ac[�s��$�8W�}�e̾�S��d��Ҵ�-�pN�Y-���%������������=E��_�vq5�t��ӭ�w61z4q'U�L{ŉ����5�as��KP!|���Ö��3zq�n�uo�Mf�pl@l��v����-oƌ�L�y�獌���@s�(���!-��f��Y!��O�}=�L���ǡ `�����2��'���x/��{k��wYu@���4�9ϊ�PHG�L�x��[S��P>737�һ��>�7s���Rn�[��if��z���P�]&����A���������X�"�}�����T'y�Z9P�2N3H�����JF�}/�a�;"T���g8�g��r�~Xy�	�ߠl����l�f�d��ؿ��v���4V(B�!b����mZ�՛����Շ��	�\Vk���Z*9�Lz$z��?�N�5��b��d�t�X|L����	�>��� ����k�"��Z�a&]`��J剡�y�Isyk���Y�I��Cs��u4}�FeJ�]c;"KT��0���,A�X����	��Q�7�ua��N��.k	��D/�e8�?�f�o��3g���J��
�E&�-1�J��U~����������S��U�F��5`fgY�`	��#z�(�|�C6t��2����3��p�H"q���W"��1>N�%T�\"��y���X���L]��P\�θ<��׺Ԥ�g��b�ձ�_��:�S��ң��w������O)J�D���
m�W��$]Q���ހ�Gz�&�w�BFĀ۱�5ᒓ�b+CJ"H��[8�P�ra<�6�)��\�ɸ��x�`1Qa`�M�8S�
��_���W:�|��y���0�Q#B>�)��Vr��+�B߀nDý��}��f�U!h��_�YS��z8�KF�z�n9Sr�����l��5��hyu��z����� 8���݄'J�K}�b�W	ΰ����mٞ�kd���K}Fe�� [��,����(�4
�>siةp:Ђ��a�9�90�L�/O	��~
�w���& e9���Q��5�6���/���|�zZ�g����4�}��O�S�X� >�򡭆�J���(�<[�d�#{�y,�ىZpЖ�/��\�6�X���_��'�d���#�u����	����'h�񎻗���$t�r���o�p"FY��i�I�+����מ��U�1���۽7b\׀��) �~`�54Ԯ����ر�]�v"�����~
�t��Y��=�`�'GU����|a5��F')\� [������b�j��40�C)&BQ�X����+�8��ƕW7��q=�CE$ȵ���yS���a
�W�Q`P�Ih��6���1+!wH� �F���3p:Xu��k���a�)�ӥ�>�ԁ�+&��n �s�	��$�h��#ު��������¸��l5��|�4J�m\,�@+�{h]臭��#�?��F�F.�:^���q�
��ȍ<��j�3�9��R������������ZB��ԁ��HH ;�j��3�; +`ɀ���$�ۘJL	A���~x��|��)4G�]�;�2C�R0Xa;a!��M�-M�8�5~7bQ2]>�b���)�L�����Y8k7en�G��<�|}SU �/I?H�uk��uN���0��5�໼IL���nC���%أ٠�l�ȗr8��f�>
���"@qn?Q��u*�d��K���}hU� ����2{.+���?�S
+��&kve��]�\ғ�	�9@J�A��#5X�DMe��8��{
��BO.�5׌8Tϐ��g�3�����>(S�N�~ɥom�h�γ� '�{�V��R�p���Ls�rr�&�`��(�En� >Q�Bw�̠Xl����oގ��$�GQ�p����l�7��b~s9�����f�@�Ў�7ƥ�&��[v��8y1'0��4S���9e�ӫ�Ɠ���l�o��]�$+�Y-����]�w���B.B�?M��n��>%��(�L�a0r�hn�w��>`���K����(�Nڙ���)�f~Wlå��P�-�E�kf�+~�H����r�2���@k0Q�f~=�i�:���ⰣL���U y��ǲi��؂�)�2㹬F�,l�=��-�� ����h������C����.�.�/^��b�;d�U��.?ks��;��ϲ_��^r�TCZ>��*Qo�\��zK1�#�w��[Q$V����*���ݳ׼F`B�axf�u��q��Cv��Ւ�o���{SwQ2��J�)���+Y�y�et	!RB�"gD�ĩ�	D?|�b�ݶ��w}�
�%�l������J�cK7%/
O�y�����st�V T��f��Z!gB1�Pq8i|���v�Ț��Puoӎ#E�cq6����c�m =d�Ծׂ�-4R��{]�?+֡ ��:�}��zT&f(�kz��n"�1���
,��gI'��4�,>
&]�� ��߈6h�v�%I�y8�ӏO���a��;N����g��u�&;?̶�F
�� o�H|rB.c��o�Ø�(��Oq�,�j���ʟP^�X��2$��CK��w7�=�"�٦��Cu�~�2��բ�q��d��6�d���	��Nt�P�G�?X)��1n˫��D�!����D�?���T��]`�)a�,2]�/Գ��a^B�}1 �c>U
v�o</6{��bJ�W��0��`���+�����~��]ʙ�X�D��$ь/�:���.�L�ƪvl� �&�0��lTi�?�?��g�|LH�/$�����h'il
��CŘǖ��~`;G���x!_W����HM������[��
vr���3�U�5����1���'9��Pސ�a�\u�0/]��3�/�������R�,��),��F�Q>��y����w��&Mۉ�������F��sˌ����YĠ�9�w<f���rӐ�nE�pfx(�'ۄ��N׮�԰;_�b���4��w~�yz�3誦���D���\�s��t�~j����	�Y򃜥�<�B�^A�e&T�~��.�B�(a�۵#��j���~L���R~ν1a��c��*�~k3|b���- GZ�,�.�>��a�E��d�9��B�"��� ��н#��x��39�w'lG���?KF�N�~��)<q�s��|Z�b��[@�C-�
�kM��A"��@�׈|dnl�����k�Y�(�a��8��_\.��Ǘ%"��HkLΨ���za��kq����`����J*�)��N��ή�R���Ю.�^����åO�z��n��I�	Y�$Xc~�0W�:q�y�:�'H'�-�����I-�n$�k	a��uo��ox���6i�'�q���h@ו`)Xǥ�^@�� �x(�Rf۞X.��ܿd��a�u5�>���~� b|A]iJ�.�[q8��&������~_�+�
���ؘV;��ʗ��Hq�k�?}�/�:U[����u�
V����%����"V�ܔ����=�h�C������H���tM���z�ɻ� g�ޫ?N�9�EU���O� a�Gq#X<ִ�ns3�;G��H氼L	���|
�Y��de��D�g��t��s�T˒�F�W3��K�7JrκW�OpA.��m�s;�ղ:���{W���Z�$���o	��\Uƴ�ؕ���Ǣ���K���h���0�&f��+��w����-��Q�8}��[1�|.v׵$#;���?���۰�+�+��%��V�W���#�ҧ�;��͸�'H���>GC�$���{z�*"sc��M�/�z]��4�c�1��&FY�\�2u�Q���������u~��н`�tX���4#J�1�f��3��'��㆜��`ܾ�vJ���n(�#G�5E����$�J1ྎ���m& ����}|m�g!�4�Q���nm1���.���Ҡ�!�E��E[@���ko7뛳<�����%��"�h��Yζ:�1�0Śt�7��/l}�'x�x�F��!��2����h���؇֠�j��ȑN$ԉ7�$��BC{���\��b��2c���Ok�-�~����	�l�/d���rJ����{��a'�*�B0��?��Eu%��ӣ�U ��p��-�GƚWc��q���k<����j��-�3z �q:����HOO֨����]��s"+��T`wz�D%M:܇΀�Z�ս�B�X>(�і j�������C��%~/}�ux�n�L��ͳ��%���Tϯ��7ZH<�HJU[�7(�{����,�>˺�XJ��DM`����#t��F�`.P0ĸ�w�8��*2I��d?5]A���:)�9G�z�J���W�0>jT�C�I�'�R��j�f���B/w�$}H q���%NZ�J#Yy���Vo���0�Yk��à��#Vc�yz�5�\���+uX�uk��b->�/�[ܭyo6)� �գǧ�R��ARDM=�1s�^H*2I�|���Ӱ����p�F�6�@e7\�l�0�1�:XE������-q3�}Δ$��#�D*���M�I��D��#Y�wq'<�`���1� ��k [Ì�#�Fx�RЄOO�s�2�����<:�Ҙ��s��C�R<`�!�$
����;Z�e0�-�R�ݹ�裫����h�~(�׿>�qe���-�[6�{m��}�i�K��4�Us��(�f��V����M�������Q�1酪�� (0�P��5@fW�x��d��dE' u�(� }>:��9�y���6J�3\T��LG\�|���ςJ��&�_bj�Q������"-����_����4�7���ʄ5;�OX�)>�JB2��p�V5D��	���O��*��ƞ��83s���9�}�u�9��2Ip�����sy�`ĝ�n��Q��j�Q��Y��
�c &��v5�N�:#Mʎ�#W�zⰎ����i��=���0� �t�����U���0>��7	8��"<Ax��u�� Nn�����
MaZ�)��E=�[��	m�们|��W�ۂ�?Ƨ͌H5�-�y�����5��"-�%72)>�WbR2٧Y/vDw��"��%��	�6�>I04��rpb�&2S�D�D����tR��q�h���W�US�0��zIp��Q%I��9�~����.lk���ܖ�7��[-��`'J��\�O����I��8�����#IzhA�]���j�͙Mي5��*
'�\��Ā���"n�5�>&
�w� )^�(T��ӷ papra!o����������i�I_Ǭ�ݛ=&ɖ�c���K��00�>�2X7��uoߨ�2�����i '�@�&њ6��u-����y�9�Qw6���S
�L|�<�e�g��ȂJ�}?��d��K�j	��Fk��<�
�k�[�w�<��.A]3[%A�(	�NB�kK�n��=���� �.�^�=�s9��2��H&-0Ku�Nk��)�/��L֠0�e���,�7�����>�cr�x'�V�͸5�Q�Yd-����l=�l;7b�C3��6U���/k�ls�-��7`>}��&�R�
�U���w/��rpjc�Y�rJ�g�~&S�د��N�y�?o�=m%�-t���n�T��m?���_D�U[��e���X!K[C�P�j�=.�е=������P��W��"��5U�I*�m3��;M!�DM�7~���#�]R0)�K3��m�vS�2n��4��t�/�"Gwq���U�ga�M?Y�z��?�f�@�@�-�lt��ᓺvw���6�1w�tx:�n�(2Ew������<��8Ԅ��voq�	����o&������'˲)o��U�pb��-��΀YC�ĩ�F޶k��3�7��ɣe3´B��>k`�4�������
 s�F3��	{��6~e�It��!.�f�sZ6��v�T���-RfC��^L�E[h*���iɭ�,n<;?�#@]�.n=5iu��g��ɶQ!Q-:�&Ӌ��M9<�� 
	ːu�"}.�K0�4]V_�)+�B��T�"l�
�<?.D��QS.�v������
>��=Dts��]��=�ʅ�I|̀��<�V���0D�.��n_�������T�Q�I@��@0���_�E�/�(2���L��]{v0�č`}Q�WY��d��� ���[����Pb
"�v��:/,��S��eaK�D�N���N�LtM�P�
?�g��2��]� J۳���Q.��)��Xs%�3.c��V���!�f���z`��7Qy��^�m�1McXժoU, ���|��� ơ�A�¹K%W���λ�
eF�]{^������}wh��m2���~	||Z�۲1�O���u��r�@�!z�0�P��u`F�nMBV�l��n�_���v]��YV�p"�Qi�3|���Ƶ��� �T���D����a�W��|ή1�W��y�F�j�V���څ����wO	?�f3%���>d���P�H�������=���v����1���[�����w&k�t�K��gË6U�q_�[,���z�7du�s�F������fi`/I���j[m�*&e�U�pҗq�c��o�-��O1�5M�} (8��@:S�t��>j/);K�-W,yV�hc�p1�0��x �
����UۖO2��ѩ������PF��
`�
^�]�鋶3.�3�U��$h@�S;l�p�kS��)���~������_ �f=ePa���v�0M���DT���hP`~���m®)���~���=-��UL�q��9�L�L�t��6��8K�s3T��(��U��a�z����[ѕ�5htvY����!O$�\(VB$-�C�dl��LQ�C�Ns+Q�I�� �g�!|<~�O��d�kd�j�ȭ=���X�a�������xy��q���,K�1/�����Z8�����t��M��3�R0����B*d���������ƔW��[v{7@ƛ-�R�곕���f(2B�		��xPXސC�,`�VtrD8 �c\��<ID��˄[3�k�'ԍ�ڷ!Y�'R���US��� ����jT4��T9/"��c��(�۾���cM�;�nפ�Y�(J ���xG�d�i}���;nz��?��F�k��1qמ�8Jx�Xl��3�qm���|ὯA�O�M_���-��͹���ݤ�`��Y����W��I��I��N���X����[c�*�&:��͞k��b�"^H=`��u����L�*�v��T���ǟ�hC p`�w��yw*�q�p�U-k�S�s��q�o/�B;��
��8r�[�
q*���N�˷窀I�Cްk�s���O����xj�McQ�f�N��)�B��˹*\��T�T�3��.	���X�с.�|�Cw놮�2����8cjk�~�%�~n�LT�!�[/E�]"��4�j })I�Lʟ���|���s�J��ǂ{�|�s*�97���?A�q*���c�/���ű�#s��3��h���?)��& �����(b�Z�2-����8W�.@?F�y=i��N D�`��Q�W�u<���ݩ�-�B=#�X���ͳ����7u�G���]�	�#sך#�<���q-�}���DxOwj���
5S�n����Xi��ɏ#b�wX�n���j�:��n�6��!m'�l�C&�hw��Z�c����~��S'�7No��K�4v�7N���*�}�9x�74���P�	3!�yn�P��lO�jf�,�.���f��f1����8%�QG/�N@e�u1�؇:�H݀K����.�OH��Y����"�n�^7��r{��R\6yO�kU���S&
�GW,�!������!��Q��k���X�!���Cm�f�#�mx���~(|Z���xst�cN�����:�EI��~Ȋv���WgU���m��ɦ��9���2v��m��
������r�"���{�8JtDOҺ�CsZ&�!�����ܽ>��o	�V-�5�!��Z�>�&,�ѹ�b�)B��M!d=7�AxٛbT�kv:3�	x���&����.I�4���&qô�M���~*T�z����!{�[_f�Ѣ��A�k�Fnz;�D�[Q��8$��d{wU-$�
шb���e� ��YP���?����=�b��/�c���B� 4� �66f�O��s��΂42S�N��H˖��K"�`�:����3]C`!�W�2������Z������R΂�-)ma۽Q�oߌ�@T��p�ec�v2�+�����ڀF6�f}��h���A�\6����p	s���U�p��v�1ҔS6�o��'�Q�T`��Q���h��D�s<�g�d��y�!���T�bX������~oQ�x�s,��PВt���K�[��R����cۖ�m���B 6��;��ʎֱ݁�� �+���i���&N���N�:����<s*W����$�|�H���[9��o���ycWa����'	�g�d�5,`���]��[�1̿"�x7"�,��&��x��"NO��s�~�@^��*8�x5�I"��D��mU�zc� [%�'���.�ڍ�8��|"�o!������"U�F���\��'SZ]�$�B����ށQ�Uد8��G��u|�p� Y.:[W��{�Q���5���^֗���B��ϱ3KmX�Q�^R_�����v�d+�D�oWi0��=��7��k�J���rn�tU�W]�Ǝ�|kAD#��(�Y���y�vk���Є�>p{��&����W�S	_�Tz@�%p""�c�|<� ux��ES ��(Aj��#^���ad}�������T"�Q"�����YU��>|�� �߫D�J��c#�Z���{�N�5�$0Xko��Ȇ>�!��{ۏs���E5PE&�{���H�59țp��m�Q/P:)�����3���*���|�J��> S��r��yl�����a�W|�m����(6.�
�Mc٫��RXF�<��s  ��>��z9��Y;&��XN|q���ir�Fk��t�6��U� ��^r�]�3�Z�_�I0n�{�`s�<ݽ���3��?io��)�VH�t�fJ6��
�,����b���N�@{�ڗ���; �Ǿ*�7YA�k���C!Pj_��;I�)�̒�N�iގ�M�
�6YtyZ;�C7?���[��h��&Rk�ǨO�P��S��<�"/Nd%��;�z��McyB��6.uO.�0�
>ȭ�,�2���7mS�Z*��X�J+���^�¡�U�<�OR��:e<�?�+��ܘp��f� ��J����`T�����G��"цh�,�]���>��-�G�s3�B�k]
�C'�kk����CI$�B*����~�!;���i)@�׆h��j�|}O��Q~��5�x�V�a�x��I�;$V�%ɴ��	't
eX�h��8�tOB�V��I0���0LK�۱��o��.	��Yx���ZI�B5�� ڌ���e���V�}�_��c0�WX�*�}9�T���j�:7O��t?B���U_U��c���r�g�Y,�݊���f4��j`�|�kg8���U����J~�p�v�$����uI��;#:�+����-�Z�[���A��]�3�&�~���T���KB�`H�H=�styt��g�ME p��R�s�Y��V�δ��7�-�
񬺬��� �/`�-땃��� � /=���E�	���.�[�c�}���k���T�BY@� .,!��["�D+å�̗񖰪��eGF
���kj1I[�t��J��I꭮��!w�@X_�}i��1ʯ0���Qz���Di7���g'��b�l�i�:7���Y�ǌv~��
�L�Ż? ����������TO3��G&�0aT����R<���@\;�8�4�63dݗ��6�+�E��dM���?����ՇCoPq^[%�1ړKn�`�>�+�����r�Bg
���繒����L��V��'��+ǧ%�u��:R��5�F�����:�|��X�=���F.2�y�&����2_r�{���������	~�<H�&<��G�<AQl���
Y_�+d�)���1U�U�B�m:��g��l��T���͓n7NUL�������R2���g����BI��	��kQ���B�G�xK;�W��[�&"8frE?�a튼�bKw��:��7���֞F�DF�9�|x8.�����U�9�N���\b�"���"��!}�Y���cMNS�r��coVoG�K�U ��R��k<�8��*K����Pt�s��:^��%��E����z�f��!C�.$䲞 �3���L����Յ�|T�������yk�ku�'/�w#�C�t�h�����G�๪����͊[g�)Hb����Z.i}�`�;��{�fa�Loۡ���ܐ�7`d�X7+�7@d����4��.�۾#�fig x�O���{�pJvœd=���{��o0�����D0�O��(�r�o�8Gc���H�`M��5c���OL�k[��ү����M,}��>�GS�r{�{La8R�:�h��oH��q���kpP=��-i?Bb�X���<��oHlb����)���UC���:�K �a/��=Ħ����f�"��Y�0;)̕P=�"/X7qb������� |ڙ�o�bco����3R����.ARWCl�����m�5.qp�;�cO���~�c�;�?Idb0*� +E�3¬�� v�S�0Cg\Z8�ʊ�e��������j7p簤&�"�54w-ڹ=J6��Z��
\K��Y��4��:���O�`�~�R�)i�:O��s�?6<J�!*F�sjҘ�hи��!>Ig�"�\��LR���_\,+�"&�j�@�����c�l?%�+Ħ�?1�r�Ƌُdz�6 g�{}�����Vi��A(vu�Z���`�2�*�d��C�lA�M�c8MFK�i��v8����y[�����,XZ��h��kmn��?�M�@W@���V��c����]����cX'"��[B]G
q4�ҧ�\`N^��|���#+��8e54�Ms��ț��4�꽉.���~�lX�9�������ev�ɒI}6_\������ڡ�N��<#q�3w"4�V�k�g��OJ�:��š#IS�d~��%���T\d�s��D�U����㵠'�
�Ha��Z�宆��6�a�A�;�����`���[D�����N��i�g��K+|�!���<�y�u�(+�@Q����/@*H������W�g��M,��Fn+33c
9��	/�ϰt@
����/
��p�#�e��~מ������>�����\�x@��@�hc�%jo�*yT�@$�����E�k'kOA��Gk��'!��e��H �6ة+V�
;�.�2�$�ȴ��N���W�ãK�
f#��kz�68UZ=�OJK��KW��	z[�tZ�~r�p1������L|(�t�"QqĈ�-d�WlL�߭�C^�Q��H�.H4��w%�1���Ӥ�/t��>]N�-�B��+�<��9�fa��#r����x���JR�2[2��<#��6C5��$�]4ى)*i�o�!Nя��Ju��7Wy��d�`V���`��A��FN����u/j$Z����3ӼF�6j�@]uw �4+(�>Y=6*I){����s]�1��^��j��#z�G)&�'!��Dp�fv]ЛEt����aR$�\�N��&⟄�n�v��y��?�	�����
}/��2�&��6	�׺Q�;TIu��2��Z��b- fs�ݲU~�B��S}G�#`%��9��<=�[E%V�#Z����o�.���I�=b"��,�� ���n���?}����	�&�����T�tbKȋ�l��%�s��n)#7���ۻ�G���)�+k��w�Z�o3���O
0,��
��
�y',�������Fd�� ��bh�)��{O�>�sᬹ�~�w���h��l�t��T�0ߪ�U�6�~�T.��SPd�0�YM�	�~�	%OtC8�"�c�ꄔ���m��� �ڀ�w������q��������g-ԒQN��/�r�n�׭���F�*�:��#;��d��ɵ�3"�)�i�ױ�?#�X��n��e�L�}s�-R�]�%�Tv�~�����di>�������
�>(&�z\d��G;_�_��j�F��6�X��"��'Zr�=?����ĆSy��|�L�^�׀�aVV��Z��Lǆ���^+ϧ��ߞeQ�9��M��?#�-pi��6m]���-a ��C�����_8�6�h.�f��ʣ��&�C��sq��_'Ə,�j�'\�����8���c*d|f�,$�&�L�J�U!���⣃�2�Ҫ�uG�yߨ}�Y�@���� �9Ǝy���qG$G!ik]�>��kRsR��R�Ti�R�1wx�9eܠ���A5��r��DjL��'F��s*h��~����iZ��0̋ʻ�����g���;���/<Z"g5��Fݯ0���\k!��7�K��\Vd_�D�Be�@C3U��.����ĽLjt��o]/�;c�~ ;3c�'cŎ�JÙ�������aj	Km��0.P�~��Q!QK�WP.o_�$^�uw�0Y b�%վ8��L�7E1(-�n8į�UGF.�I��+n��"��+��3��;��ٝQ��aW�ƒӨP"]������ͳ�&��@��Kh�7���w��C����mi
�j�QIq�U*�fbPہ�z�����\���
gh����t�U-U���b{+���@������z��Z�����'���1#8|8� �0���~�BA��>a��(���#�Kb���{�;P��O�Te�D]	G5��y�p+��զKw�8�aQ,{�����A��ſ�@V�`U�U}3��Ζ���c�+����Y�C��A�\Q̻�a�v��� ?�#�uѺ��811H��M
��|��5�}u�⦅�c���_(���IE���_k[��Փ��e�&=	�E@�b���,8�\�����ZN
�h�㟀cq�zx�/F�6`(y4��3K�z1T	������6$��8�7�Q�1���X�9���9��D�j�iBqo@ �-/5Me02�V<!���(��F��\�14����f�4l㉇��g�9���vR"���� 	�(�Z�Ô@�u���	F\�L�!;vq]|����z[C���PbJ���2�O8��J`����j��Q&�U�#�Zx���b�AݟS]v��OyB��1�zgH.��"V�!o)gN��v��Y�9�-�5#�lM&�X1l��״����Kd����d+�Y5�'�Z���
�GC��ȶr@$��90��[�}�[����e؃����y��K��������Y����K���X�@Y�$��_�!��nz9�{9�h���l�Y�7��I��,_�����m��t��$��؍�-��<�p�1�L�+.2�egj���� ����:]�FK���{��	+���zGQ��l�ow�H˷����<r������!��/�9�p8��"�׶�RgCp��HOj;���ә;c�9��GM)��ZY�&�:��[d�5ę���@ط���S^�a<�8t���� 0pq���RL��(۾s󠧂��EI�+�:�c���cĒ��Ea�U؜��a`+�_��q[/w�IpG(�AĲ�u����Y8ocC�LN�}'L�ևi2��ϱ���F _�%_�8)d��nn+5$|�ȱ��oOK�J�(���w���b���}v�<�*)�=TKW>�v3l4�=E�^Zo\.�}�K-:�f�G�����'*AK8�7�I��UC�̦������^wۣS7G��$��U��k��Z�Ve�5���@U1r��e�%R���n�-v�Fz�{����^k�-�����mZH������v�͘iY�<�4h*��%�Q�?�)6��"X�֖���v�]������{@�P�t�]�	��/�Q�0&2�}]j߻h[��]�a��I��4T�%�=[b�����+�����=O*�v�O�YC��i-1]<;�@U����?��(˭�k2��a�G^cti�ĥ�/n؜�6T����U���$�?/����A��iDJa?��-(ԖO\j��1��r�F��_@�g"Sx�Ubt��c�{ �!wsπ_�~��5�~�9-=�2��Ά �.�4�������k�g�v�w�sC��k��3~0���t�-`�6�`��de��K\���]Á��sp�O<#܏v/�i*� `%)��+���~"�H��#K{5�b��:�c���nvW|�Y�����>y�U͔`�v\B�ۃ����""Oxf
�*k/�.�D���btAJ������%��}U����mީ�D~���*�P���Ae��Fį�YHT�E��Z���^9�׶����S|�n�p�xr�~���|�/��� ��ڕHLJ���k�E#�%.ҿM�ds���V.B��T���p�Zh��ݣ����ц*�T�G��CZ���ŭE�0��	��D�'�o�_�6�B;R2�i���� I򕇦z�N\}���^����-�_\Z2������5��
�<�7\xp]�}��;$�=�;x[R��������v#M>��s ��[��c^�W ��ʋ���Y���-� ��"�
A}2�!��T��o�u����X�qQ�1�v��~�\U��}�y�>�_z(>�k8$S��]���7x��=��z..o�vހȨA�5�J��/�sF8^�Wh��}a�}�AV$�}Vo�7nh�-FVÅeOƙ��-�2;0l��s_��e��Jiݑr8���0�����t��O��G�����b���_����.&�̣�ȟ9T������C�
tR�	S�=db��n�v?��*=-[J5�{��XH�`i��W����d�͹����bO!�Z�kb5�l�T��xe\�A^B:���
á�s�F9xH͍�e��]�:��Ǭ ;�'�f�%o��>^���4�1Ȭ'�O4�!�a��͗����"N�+����7�(�j|$~���R'��uz)ć�[�n�7��o���������k���lrEIC�3rw98	�r{��w�R;K�����^���B�=r�iR ������D�a0
>㐨�VL3l�	v���d7w�u���[b��"�Xir�D�T�_
$�u�2΄Fdj�"���3���<���qő1Ɓ�Y0�,e�Y�#��O�Z��m��!k@�K^��юB�z~\���RƏ�)�n��E��Gt�m�FR������ċ��w�k]<A�BX�M�@�Qd9\?�L��F]i�~bwҹde�11R�G'{)8Ǒ݌D=XL�v�g�?�'ۑya�+W?fE�.^�w �ʙ�+���i�s�x+00�=ӓ�4�*�x�iS��cG��Z-�nq�<M0�ϯ���m�
m�%i���M�� �����ƅ����=a=��c\���s0���X��x�1C_IMkO�(eW��xҕ��9��Ƴ�j�]�<���vh�>�ޗ'b�%P�%~�����aA)��W�`h��;����K}��Wq�hm^�`�I�[U�|tt�"�P�:�v�1ŐF�ʠ��&�+��dd뜠f[���>���x�m%Y p6�\��u�}\�eA�~�W��[;oa��!����ےM\p�Z�bW;'��7�?�&A� �,q�S�cwL���kd��2���T�Xg P(c˯����pk,F�)���ɼc�c��]�7���>��)t����q*��̊.�KN�v��
��ϚK'��$f�{���}s2�N�r1�t*ܒ����\1H�Q�M�32��I��lVt�)c1���iN�x�7���~�y;�IKk�|4YQ�0^
)9�`�d5�bP
�~ĵ��A�f��=f^8�wHw
T\���:���$��SU�3��ً�}B��e�	�Nq��ozXo��*�����T>�)	�C3�䒊z�)/�4��[A��dOn�i�;����i�,�b^QL���0���߭�( �&V^���`8["@e���SA��I歗��r�XMU���+)��Q�ڗex-� ��C,8�k�?zU]Ha���2�"�����?��ׇ�U�b� �^T�%s1�֐z�N�?���ߪz�ǖ
p!Nߤ�{8Pߴ:@��'rd�-���zu��V�E
��JQjHR� %$�=W1����������2K�����5�
1�]��<a-�S��Jx���m�-��C�%��p+��Q�M�K%�qH���1"�zQ���K^Uh�Q=ɭ����?(0k)J�Y�j�8k�z��T�I?�\����iA�^ほ��x	<����ҁ��H�)�-��Hx/x�w`��?@n( \��������o)��q�_n����O�_̩�k��%ȭ�D���&b�6�g���ɍW�0H��HQ�:L�_�7��ڔ���Se�8I_�]�|���S����-�b]}xM�*�R�<�C2��8fF꼎��B�A����)k��RJs{5_y����d�<�ݖ��rξ�����]@
:�q 2xC�s�z���+܍�aA�����f���LP�r����z%�[��>֚T�, ��������3�}z��A��MII�bX콂�:W�[�8g�����3�J��ˡu�|�Đ��8��@�L���t.�7.�ƹ9�z�/D �ҸB��n^/���3�N5ڭN�H/�z�?�ؔ2����!��n�>��c�<�(NV��@�zVB�'�HG�@��v�+�E�l�? 0еJ���x�\ �Up5�A:���u��qE{��sao6�8�"����=���O�D{�=���3�#�q�M��9C�C���$�pb����0x��Q{KDҊN��=+�.�eZ�hB�������������\X�TViT���9�u#�fzf��>؄nl=�[��z�]�3�;�Ѐ�n#��.yY�v��g}t�%���ڨI��!GLȊ�ί�Ða�����yH/-���9��*�vh�#�? F_o�#��qK�4�+�o(�K�W�~Ts&��Q��6�N~ ���߀�!4_A���]�彭g�Yg�k��=�"���95��7�ޔ��I8�!Rg��̃�G���"�o��=K /8��o��D��麈���Kk�"t!4�D�n����rhE%���n�jm�C\�SD؃��B&�A�'�\���pGI�����-O�+�F�+Y�m7�7@��@#��!���R��O뜇�;s��MT˿�&qǦyQ�H	�ē����VyhaЭ��I>V�E�7�����\��������_l����1��R��|c���yZg�Ȍ�|����Fj��%��:�Δ#���Mـ�+�|�^�~�o!�yFx�a[0'��!����˨��mEP��*�;��~��ᷴ�j�J3�[d\P�6�L����L86^6BR������xk���P�oy�K�1�� �.f�f��� �Cy���G-�}Wt���/��4�8����X}C^8fT-X��s���M?Gt��By6�ȺzN@�J�����f�N ��'=���3�C����#��u�ŉ���8A*v�O�����ΩyK��I�����F��y�9mH�F��S2M/����u�*�HS����ۮr���UX���k����7Eĩ�JO�-���s<{V-��^r���ZUtw��e��[y��Y���K�Ws��
[u��4� zp܀5w����_r�U���jB���e�����Xg�C�*�1�<�
#)�6���ٽ���R����X��Dr*"����3}w�um�����s�8�� �����Gvxc��N'�#�H��H�੧�M����@�&G|��%�锍ه��$HrO�'��$�[�����*�O|)�4�BH86�x�ihd��l�ֺWx &��PW�SĪ�SaT�qvV*xk��k,B\�~uEs�!}Z`?C�b�C�������M���(��*O��>��n����bo�X�Q)rx)�%?��������lW-�<�2��t�r}�;�_�[L���l��PWD�����L7q��,��*<�A�,D��y���y��+�R��� �����6�3hY��`��)b� 7�}D��/���$$� �&v�#t��sU��~�f��\�EXgwK�}�|��U���@4���V>����`+8ɑ��$�8�4��X�>ojMhW����T�����2'%[W�LR���Y�v�jY��޳��p�	�e�J͕꤇�M�t@�`ƞ�nA�&��m4�''��'Ou�*� BI){����#KQ!g�/ccV�w]�݈v��yǕ�0��L��g��y
BL����(r=5J�|�|����ѨTԮ�B�H�fX�;O�l����ЊbO@��bI�x�.�<~ϊ��]\X�f�ܪ槌��q~��/r��^��?����(��t��.���Beؐ'tQ��L���ĩ��~J�����U�m#)��x�.���q���gR���[F���B׳����q8���S)�ht�c�mb�?���^^$n�'�=�c\���a2�Ik�<&��
eoc",
ݸF8���Q+��ah�I9^�k�A�kڽ��/�h{D��1^�t*��b���R�N/���	4&0���05��.���Ǌ!�6�y�-ISI�v������_�3
�}{�#�o���j[h�%�� 3���$��!{�����NҾ�2��/:P)�p�S$��[.�G��E�:��_L|��]����]�I�o��[�����z�)�慠�փ�^��h�{m���;��,z�RB�σ_m�[�2tUPTrI{�h�rb�ݛq�L%���?�<8�=y@$ۆ�k�c�s��|�l�\uG��Q>�%��gVfp6��՚p����{�+�%����	�g�?�y\XQ_}��ې��	��y�v|�����x��k��@�S:�r�T-�*K���υ-l�gp�&;��,�� �����_��&���ӝveP�_媃��������u�AB���&X��;��=��pYjʗR� =�%�ܞ��:��:�$Cl���q^10���\���߿n��4X���.����T>�/�qͲΆ=����ք�­��U}~ �9�T��\�ɭ�Jw��`���}gYD��A6���ӈ�{wn�xnG�G8.].�������Z9�~&$������M��9�=��@��z� ]M�ʩ(��O�`�3J$6}	��Xd��+��U�	�*� �
B��fT�,�ٻ3cx��1o	]����v@f�"�@��"e���݆�T#��6�'�ըpv:V�*L�U�M���LVvT��嬚�_rE�$�X��Q�Ѹ�	�^�3�?������V��d?�O%cA8��F�U4����Z���hKI�:�6(�d�����;��Z�p8���n|Ϗ���D��ED�N|�Z�)��.,�+|^/~�}AX��@S�D`���+�>��'\4��R�﷖"v}m��y��eĮ�>E���$��8�I{4|��e�uM����M��7�
�E��N������,Y��Z�p�{�ŒN��f�f0U�`���
�b��'�\o��$�W)�4A���F�j����ޣ9?X��Ot��9�� �*��� v��q1m�(�Ӗs��]G�57��HPi�-�� ��_k��ۍnKÇ��tq�"�����		/��GDw�f����s{�'t�ZC0O̧"J<rio�a��PiMz�g���ɳ?��6]�t�6���Me�}�Lh��� nr�)��U`��{���Q����VC=���n2ϯ����e{���%pހe�.�Fd�)�͈f��˜>p�H�}�C����o\�"Ͳ"k���1���],�{=kے�����у
�<��Ze�R��פ6 �4��f� �������]UR��vu�w�d<��kzvx/v�'97�fq8���m@U�Wdl8���S��*�?��%wZ��Q#�n�����!Z��ן��Z�M�<ovi-GCWQCN���6�RϾ)��В<]�lRR��Y'�&�O���� �����Ҳ�Md����=QL6����O�
T;C���*�p�5w�_h	¥���I�� �8�v�,�] 2\�ʋ6��q����2Y�^H�D���6*� 2��	J���)3�(�j�D~Q�'ڔ)��9���G��,E�3�v� ��*�r�N*coL�<�<�)�8�!t��r�~!�)My��X
i�?~L\;@*����!�
����H�75Άb���ه[��"��@��
o]��n�E��7]�$~�ƤF����?���
�<`����z����H���<|a��^��վb�Eٹ1��U�3���/ج����,��k���_����_�
�zD�5K�'"��y٣:�`����46����n5̝�I����V� �j�l��F�g�U*�F4i�Du�l���r��˩�q@�4޻�������̈́�w*.��ڪ�M�ԕ�O���[�{�t�ӹ<x�?�v�<�O�;�EΘOȊ���$�>�L�=�+�BS�z;[��]�%Z���%ؾ�y��ʂk�!m`����ԢS�&��7ҭ�=x�����ꆳ-j��95k��v�G����S=�wQ��ɽ4�;���<B�p�b\|0-�����%�������xZˢ�	m�p�Ŗ�F�C�[��cc�Н�*�%�(t	���Hչh�%I[�	4\㐝|@�Nw�fLJ'���XW>�u4��I^�ʉ&��w��?���M���I���{�&Y̏���qƳ5�i�M)�R3n�z����Y�ߴ�_�N�󆁓��pT-V��D�ah�9�=�J��<����50b0��>�VnBo�&ȡR�Y6�1y#�{�����ʕ�vrq�`�����W�Z�A��-��6vo�?��A���|6����0�����{�@W�&����<2=Z8���pe��/k���?#�\�������y��0I�:�av��?���C��b�
�xhwF�ӄ��~X� �3W�<��2J�6���K����{$-�ˡG-��[U����Ł]�f�\�<��٤K��{�Q�,ȨD4���Ph�?{K�9�&ׁ�e��`l%dh���:J}U2�L���Z���Z�}C��9�c���U�Q-Q�p���,���÷b+|����$HD'I��jG\����h舽v��3���;��:VSwO��Z"]�vR�I�,���8�2��>XC���(��c�;r,��w52��a�tG�0�tɢ����⏏I��k�P�}�����J()�B�n�5W�Qn�o�m�� �{A��ρ��&\�DtNui~$V��si���3�ڗ�r�8!e
p�j�l�X���+�C�R5����:>5��:�yu��g�[^1��w��_�5����s����j��XϬ�=�]�&簖h~��_������7-�<�^@��'0�o1K%���k�t�Ά�����L�E-A��˷�_�9oO�oK���:ot�Ga�fT�'�O�N�bb)J������S���q���&!@���v�W6����v�)F�����)��\a'[Q��R�k�]c����{_&��/:y~��W�ޛ)(���n��ë�+��e�4QS��Y��y%'�id���5(�'ףZ�o��7[����)뙝)�hR^{�_���0UF��N&�60����-�,�}���]> gC��=_I����~ܖC��s۠����|H��^v��a�r_��8?��QlQ3���,����6a��+�����@*�n��+��|����,�X����WB��x����lՇ���������i�,ͪ��Q����5vz,G|'�^��&��SJ���_Ҋ�>,}�R�:�;|B�{e��3��,�G�]��$�0�^�R�q�U���&�l+�a@�R�H�g*���K�K�Vhbj9~�{D�ߙf�葬��d	�5��2K\E;�������� ��>��Ig����_���֡�pn.)-��S!�{��nU�1I�&1����od7zF�%��e7P�D����e��c�K�k3ii��G���Vx�����ۜh����fF�2zۑ�ֆ�hzٝZ:C�9%����ܻ6Dt�/��Y�M������؜����O@7K�1��aX$Wh4��mm�'d�ڔm�N��l	�>u�{C)���b�	 �`<@1ϗKSm;���	g)籜Ԕ�����"�-�����c\��|��(��oC��A�g�/N��fU��֩������ يS���c���oW�Cp�N�� �j��k���]�3��9opFy�o{�cj�n��|fI�8���� �v]]�GV�F��Z���]�l�T5Q0݁|i���[u�}z5��@>��7˞[��0PW�=�'$9_w�Ű��Be�F�r\�1��V[C�l�f	z^1T�چ��&q�	�TF$5{������Jϒ��7�Ii �5��x;kA��1�P�L�B ��j��o�2��lT�$�3�������x�H3�_��B"3���$���0�	�"K���pw�����õ����KhN��3�lGM���X������W�&b�h���Ôr<�Y���d{Jj,�&wmT���B�$MKjR�[D�]�����?����UX��Aa��W ���^�P+@F��`�����j�Ob#c�kC��e i���d�<�wl�
��7���W�/�ĕ�`t�/�9wZ$5��V^XI���5���&I:���Nn�Ѫ|#�H�Ԛ+�B;xC㜋K��Ʀv��v&�#�X���I�v8��_0]!mC�RX�\��K�n�Bǩ�F7��O4�����5��!�!�weC�)�����9�cD:���:���x_�bMm�ğ��� ��問���u��ݹ��)���10�kA����|�3$>���R�9;����	-�&4�ིP��;H�xsTD���8��7�\�Vא�ә��r�:.��z��Zr���Y�Lă�d �^����ܕ���%�4���ٺ���*Iǜc��j�W���ӽ�`k�y_'Z�&��|C˃�{�K~�m��Hȉ&J˱�Q�3łk�+�]��a{��S6GNw@��l0N�28C�\XL���R�5�i%�=��,��,�����Z��'�G��)�dj;jRK^��,��XTl-�����vf�#��kI���4����х���:������%M�b��i��i3W4�����Cd}�pHޗ�|o�`sY��� S�oBu�)�۱�Vy�"3�P씯ؚ��2u����iOT�QS"�@ܱ��Kp�l/�5��J��313���-�J��t�yRZ�xZ�4Kت|f]A[��e��d���L'I��p���>�"�74�O.0��*>��@G?|{)v ��1͂���U
|�ft�Ե��||@�xUؓ$+�Hdr�e]h�2�,~b�]�|�<ź�e��*2�,�Q�5�,�$��w�tz	���E�����g	4gգ��#�#�̷@�|X�i�݈	���������rmZ.urY|�R9-����7�%�Ѓ���L����m�����(��"vp+����_V$UC삸��)]5����RS~��	�P�ye���;g�͞{�jB;�����g/F�IԿ�*Lp{���K4������&�Uy���F����?,S�bQ��.i�Ѡ�-�C�3���T�Ӟ[U�d�����9U�x�[�[9lH�[5^Ʒ���4��toc�ϰ�ai?W^g`؏���I�7ЛB�K�c��:M���zYR�t����4Y���7|T�����Cc�����7#����}��o%lC�OQ��%����1���A�a��C�!Zg�QK��,�%�7�qۜH)@Q
>qL���Q��p���=ZQUf��f.���U�n�m�e̦3�c�A��<�� f�a$6 6��p�ŧ��a��EJtU�+Չ޻/�Ѹo���J��ֻe����ou�$a#��ʠL��GC���qzX~�%[bOe��+�\ hӄbk��K0�s���C�WK:�����	�|'�lg�E���ޛ���O� ޴���i4�"e[�FM�,!�~�*��bT��O��Q��Q�ZQ���֢�/�jq��*MCa��9�")/U)*p��P�W���X����(�Թ�D�b��t�(���Q��kd}�?n�V֛"��'�2��,����98�e{(Ԙ 5o"��h��n��Md	�U.�L������r����
���7Al@�8���P�x"�%/��0�d��p�0���78�T�E��o�,�~N1�Bj���mP�I���#��w�,M�wl۟d_����m���2�R=�Izt�2EcByY>�FZ w��`U `4h �0Y�7�lKST�q��I����AjG��Y,o�Aw� ��k��Rn�GWҞ�7�R��Ї S�'�5�a`!��3U�CWဘ�����_f�GoOԂ���U?v���}�������xvy��`C�ϊ�G517��N�E�M���x�f���2��Oí�L/AH�&��z�n��N�kw�y=���0�ajD�(͹��G]N���ns��/���7���PIHr-_��S��-��G�2߰5JG�2���r�Y�m����Q���Y�0���t�\��5b0Wt%�Ĕ�2�׵Y���d���U�5w�����������+̳�{�V�G�b�Ѷ��a5�l㽩Ki��!��md��/�A/jv	��0
:l�"�l����,�A[��hWx���kY�J��DN���_�y�b��Ϩ0H���W<�ѯ�>V��UF6=�AC�`Ⱥ�r�1���^4�69���E4��C8�P�	�헁��"��)B��A�#>P��!�����Ed�6e�2��6w�>��S��j��t��\5j�4�gX�A���>�dq�qeC3������1�Rj��K[m�C����R��bݪ�U������5ぢ�f��<��]�pn��>H_t�E��?"y5,ı�m\Akk���T^�4c���GU��JLv�w<i�Fv_S�� (�ޥ��s4��^�.Iy���&�A��ݛm�=��_����}�4��R�̠/Elџ�'�)p� �eS�iP˵���A0����R���D�}���!_�A��-�(�R{�V�P+�Bm�&S^D��|���h�B����a�3���$�m�l�7���u�,R���O����n�Әc�Z�6�͓;Q�qۖIT"j�sca��F�<r	B��Y�I&�x�"Grw(�#	��/R�Dm�k�H�x�/ꌗ��'�]��Ue�g��4��fE�3�m�����,�a"·J�0kK�/��1��S\7#�)�}������(�	��b�~l|�Ⱓ�ZyW����WAfr��͖�E�����-B=�h_f��,.3*?)�?S��O�2��Z<b�_E�чy��C��� �I>h1;�pgG+������GrUT��Y�-�>���oFD���gs0T����(<�}��_h��U��S�B(K�5���֐��P��{�����7;l�QL���a�����SL�
��#9N�j||�S�q�y�]lg0$��|��t�8^�X��LJ����H�n����S24���"X$K�Y90�#G�V�ڬ�}��l���~l6�HN@|���&ٻ��v�w��L��ٙ�۠Y"�����q�H ���1p?��о����<�Ϣ>P1?X�uԇ��Z-�W{֮?Y1m+u���R�j�w�����H&�^;�XP�����g+�V��Y�7О�s���(J��Gʏ< ~%���ѳ�y�Sv`(|��dJCy9+��c���;�S��QfC��M��c�%�	q6U��ǉXZIR�`zf��C����63b~�٩� ���p���1�՗��}jE&r��3��,���*�m��oX����z�lm#q���ߐ������ ��m���$��Jb�\����|�#T8�iYz���Z�nޱ�O��������F�5�;�o�W�W�t���[Ԑi[X+�n�N�J��t��fH�����Tx8�Q�W�"C���(�� �<߼+�w���V�NCLx H�r]7�E�p̗N8���O	�P����#��顖�A�v̧��x�626�!��d:LH��j���7������"�����@/�4L�/<��h�( 2mI�����#�~�
����T���<�'bN��`Q�6�\r~��H%r
��4~����<Nwlb���c����^�w��<Ή����G�>��T�#l���&��Y�)M�W��PЛ�"�sH ����#1�~O�3���M�cWc�@��lKZ�ס��G凃c@l^^+�Q����m4�[���b�=g򘞱�nWk"�EVĶu
N���w�1?�]����`:v���k�U�&�-�x��kKW�tZ����Z�X�z�Va+��g1 ؿ� q�r��ci�X1�M�
TZ��׻�B�ψ�K�Yt��A�l��@VB��P�A�(���*���0d���c���ϰ�*�(9�\�2��U�M�	���Y���4�
@4	�΃�Z ���q�W�a�(�m�?�ˣM�#�|�=�t�^�c�3���7��v@��D��xA�8��e��h�'Є��ߠ0ػq]3���p�=+�|����n��#������̠������ӷ ��J��E�6���L����B�ֳ�xeE��������W�q`RV�f �]*V,I�ᵓ��^[ZE2�R�?�!J��ֻ<��e%���SB)����ܖ�@��p���z	R��)�Ktm��yyL_G�����*}��V~h��y�NA�;F�f�
�j�ߧ������{��r�\Mǹ�s��)@���P�˔Y������+���x�~��~З�p�@Af�
�E���E-%N��:��^�i�CyX>�R�d�q�WQ�$8L���20lf����b�.$ӁY>�e *�T�)���iM�F�\�{�DR�?���)˟��wX-��ы	�3�`�x��v���=�!�B4�?u�n����[�^C�h��L��7�zh�4,�F��nR���ݬ?r��>�֠I��y.�v_מ}�n�o�wt����J�ˇ\c����;ZЬ'�ܶjy�hl$Yk�/�f*�nM1!Z�Q�8�/EYdA޽�A�H��`)���b	�so`ƾH7<yY8���R�!#��
u��<rΕ��=(�O�Y�_�"b���d���Ϳ��y �bx#�+��`%��r-.��(��V���p<^w��C�R7J���y��8��}@
�p�шh]X;Z	�k�v<���	~r��U_�����B'L������IdpJ�����i�XCt���s�V��Ф(p��H��V�(*�
��%^!��Q�L�!Qc��%:���:8��uu͘X�c�P�؎_M[2i\����*��(� �P,`#��H��D��w�Q��O?�J3��6R4ܞ|�+��t����M���r�PM<D��̉�e;~g��Hd� ,�\��\댽��'��9��7�i�<5z����؆ʬN��>�Cq�KA�����̓���Fq�A��"3[���*	�����H�u�a�%MM�x%�C�F���
}YI1�S]$�`�w]?$�|fB�QU��+�/^Ap=��=H�6ܗc>��`�۵�<1#%�^�sEx�-x�pfG�ck0�}�������)��Kfv����r����[�*۬%d]�~�=j�}*B����$���m�n�L���ө~)ڎG��^E�Z��A�E�P憧X�����2��d�?�9L�b�r(��l�GŢ��9�ކ5��W�I7K{�
<L<�]L�[�`�n�{�Z�zk �G��j#Q,�M��y�]o~�#�7���t�L� 5	kd�&g�\�� ��u37pՖ��E�^�fq,e���zŴS�u9wȹQ&�>IE�Y�i���H���dr�ޔ*�ýb���3�}.G%޾l�%�k�b4S��<���g�CF|o�?%�� �یS����c܆�ip�Kv'�q�I��M�`%��ĦYM*lD�'���9ic�q��g�xĉ�g��.ͺ�%QR�����χ�C�"�ٛD.(!�?���X;j+�9��%@���\]N+�:�˰��̦���j�Y��x���y�F���l��)Gֵ'NeR墻	g��*�&��	���(�X�����Wq����kX�!�sR.e����ஹ�;�w����D���D�
��.~�Nn�V�k
?H�j�hM,���b�����2�0��Phi�,3�����.�L�A��b\��wg����&Uu;�c#^*BX\NJ1��ș��fP!�? $&Y�	Y�� uuN9Cv;{wv-�bc��6Z�g���JU�J<��I�Dҳ}B�3�p�a% xRW�>�w	��T� �����e7�4������̏)��ZvT��r��@<}2�W�j��W����)B]�8qF�=�Z��4��������H=�F�� �<ޏC�S��
�|�D�D���q9�r{�iZ�f���-��,�f�e350��I;"7����F��4M$O����%1  �g��&[���ދ�����-��O��tt?@G(Ŏ$9�M��og̚��D�9�q�-z�L�q
5֢��I�D�|��N���mz�$#�E��/nP��x�S�=������"����]�u��DB_��Ð�@ǘ����^CM����ߜ�j'�n�X��t�����r��~��6䐘�tDV'M�.v4��+oIಚɥv�.�)�n'[����������n3oP��m2�j�3��~w3&$��+ٹ�����n	�E�G�a�}vd��aNS�$�V��o���SG��0B��4�����^3���w"�O�f�dK>HrC:v,8�e�o�(�`@[�|��y�02p~�ʥG����5{�6���E�)��Hg_^o+n{���ce�K����4KIe�N�������*���2O�sۣ�HEj�o��J�/��dw�]m�ι�u�k�l/+h�i|�j��j�2��7֩���~�d|�P+��)c�c�Bm*�͓��%�
X�aD��Z@X�6��r �sh�EQ�	%2�)��3��,�M;a�E�6���%��4]��&�%�ζ^>�/u�k��#�,�YO;ۛ9���I���/��>\��dgՔyʬL@��IJ%�
 D����O��]�����q�]�h=Hʼr�R����r"�P��߰`��<_�D��y�H"��Ӿli�/h��t��t���Q��o�I"\2O�$��g�G4��Y�p��9�M1�������`6ZF>ϝ������@�
F�q��<별,�׮�Ni0L	��L3J�@&�my��-�kS����q};ҙ32�@�>�i��=��a�|�l�V�,�I��3����I��3(m��m���IJ�-G���&i����b�o��!KI�����IZ�u��.Hv#���ʓ�c~�[-���n�.E�ќ����+��¿㘍6|o�N��3Y_DS��x�@�������%�ױ�i{�\z�:��)��T?���]�"RM�e�A��]��v]�{���޼�q{�4�J��1�{%6��ҝ!��w�a�\�ы�����+��T҈��Q������AqU��n"�RH�d���������k�b����g��Pv^���`��O{��z����E00ck��#��̏�Gt�y��hJ�%9*]�.5M�pEam�\�q����[=�(��D��r�u�Hu�̓��9G����-�<��0���>�����tHZ��p�_�ﱪ7��%����p�o���X�aG-.�x#BSb`|�k9������3�#+w!�f�����߷�P���WqJ���ɀ�y+�P>�.��e�
Ui5b��o�0M���2?��d��l�b�ߺ�=�U,g(���L"æD�d0:e%r*	��['���~ܕc%���1�Fn��4�$�4��ά�SY��5.�c�X��K�Z�ߍ�9+u��r�!9��.��^�`T��'����u��
��PdN �^6��e���8�R\{OgYq`�=��w#�7Io^1��ly���V����\1��Й���*Z@L���9�4`c&_�uݢ�*M$h��[|��j�0�[`�$獮N?p��'����F�vT�E��琢�������9wQf+�RͧV�o�:�4(�?R=��T��k>Am��]7E�% ��\�*���c�-.L\E<�֜D�կ&�'�C�s���|D�40+��5�(�ʼ/��l�Š��]ٍ�E=y�ig���TǴ)��X%\O��n��_�~�e��<����GMq��6rz��oUM�Ab���8�4�b�0Kn;�FX����v�1p�!� �p��'�9���NȜc��^����w��J��N#eǗGlh�^9����6�t���ٽ�
�a�j�WE)��I�{8��N��Va�[(%��|E�J��U�e�vŰ�T����>��Fݤ�I��fO�*�������g�y�H�F���ݳyЉߓ[Ly�3hF�ԣ��شN�xQ�6����7��֍�3jL�l�}7�Cm���k�D8c�(�
0���5����Q����̘�O���f5l� �n���0+?R�I����0l_\���`hk�����w���8�6k
a�u���z�..�D�8D��D4�0)��D��-�k|�����#֏?�W�L��kâSh��A��Q�ǔ�K���`*D���h/�]�
gƤ��Ő�Rx)0��!{%�9%T��M�"'[�ă��(���]�D�i:���Q�^�}#mJ����©�Z����`m^�v�,%�3�B�N�JM�==*�v��ם�� @�vc�3UT���
ͦ�O��A6�&�>IK�:�PPG���y=��_��Dv�����@�<?�S<��?v2�X��c��ND��h<$�F�tuL'�R���\S�\xB��[n�Z+�������mM�l,p�4XXL��-XRO�N޹���hJpC�W��'�Ѐ�m�h�c�_��^H-��ئ=ZW ��s۵���|n� �.ū�l:L��=z����z)�� �D��N"�d��T$d���AP���@W�e�
_3-
�������e;��8. ͟�$;vm�ps�p<e`��]��yCagӓO~�y�݄��3}-C�_� ���h�;G�����
�i��:D�ػ�IP�H �7%U�9M[����6;��pI�|pu��L�H>sǓ��<T�]C�3蚮�S҃A�E��������Ǉ�غ���s����T�e�� nB��%����Q�7 ��6������c�1�д�}��S���.�+ݬ�����`�VP��'˃�0��C"�`l8��>�������
�@>��7�؟T�.��Ǯ���ҲL$е��l�4�0R�[.)����'��-A�{K{s�;�hm�Ym�G���4�~����9T�%N�!7�D���$�Cu���0_�ܮ�:�հĨuN*VH�	Hz"��ȴЊ�)H-ן�ͱ�h�[K9�\[��cV�v��;�A�4�siC������fgk��ew
!Pw�8Ry�/�����8#.6�+��'��Ȳ��\)Â6��(� �NA0��=�����U�!	N�l)b��X%��
͛�&�tPP٬}��v�NO!�~A4ye�/�r ~����w�>8��ř;xH�@+--�x���r��� Z�oψ�+�E��V����v$+9%[�1�������/�XK�"Uc�?�6�
�~.���R�^c���T�����`?�l�z�DH��۱�y��c���ᐴW��'1Au��ӺQ�~�'b��RKε�ry0���_!�W���bHpC�
.w�K��oR��UQiD|g1n����+�E�~<� �a3�	�L��������6;��l�њ���4����2%[�.]�4<V�ɱ4����]>2���*i�Kq�j����Ȋ��d1W��2GD���Z8�fc��7�Ђ`btG�d�9��yOX�ȝ�,�t���t����ie�C����� ��/,|@`�<Y�U�Q�v�LL��ީE�w��>�����:�o�'�w6'��'�@�no
N��*�5E�?���:
Jϫ�.�آ#I�P��_��}T���.jd�l��)�W���I\"a�"���"���x�O1�; ��-�*W�Adñq�l�K�2E[�<��6W���ďX���CQ%dw4a�8*��` �'���@l<�����A�T$|J���4���X_���+'BNg!]RT�m9K�h�S�A�Y�&�/
�8X�ts�<ԯ쐹���y��ƓՏ��v�^S{#>��]� j�F��AM�jh�3ӱ�?܄=�.Ӗ����}y����q��"K�s�1](��Z���A@:�D ��u�/�9��}:~����_D�5��wZe��5D���n����b�"�5�:k��sF����/��UZ%�Y���8���ΧV5�%�oGp��_�m.��=o9��.�c_( T���Xdf�����+|3������ac��B1qԔ�A&�U����lEtDN����������XD����T�����lz:]�']��tJ$��D�d��� �bB[�3\��$7��Â�z�_Ω�
���x@��V�d���?�	c�ߗq�s��4KI��t�O8�����^�a^����_xQ�ݩ\q�I�cZ�v�U��#v�cqէN�Xj|!*C�rz7h�P?\��EU~7u��>̰�	z4�X����f���Lz�lW-��U�����_��îEΘ)����;1��v��)G��s�`�[�.�cjJJ��Jo���3m�}lsР���
�d\�U�9���C��U1��aI�:1/��d>�CV�$?�j��8�6?�r�d}�:`�W���C�L8���aM>/�ܰ�
��Ə��GJ�	#L�lR��q�?��C�y�w.�PW��5���Ɨ�7X�����"�g������5�E ��;����b�!�e�V���$�TO�PUgC�P�X�U��l�����nX�ϵ8��g1�}@ڕX)T��xLscAa�.���H���������ʣ09��@EM�?�^�_�U)�­��Ɋ���qsʗ�L�M�t�����U���~!�ͅ��]/x#�i�����ˉ�����d]g��GH��B&n�-�g�s����D.�\_4�A�{St��ݮ�䯍	���G�Wyw�m�ϯ�o��%�Ku� �渃�cD���	��A�$��N�����jst���W��Cs��Iy����>���j�Ȯ|��N:�À��o;�m�%�r�J�	m(�m�T�9 3#�w��&D�6eуJ��Vn��'3�j�':
�O-+��!�F]�d���g�DNtG�G�$�1|��(�l�1F��,,�W!<�<�/�"��y�Ѣ5����P�8ĺ-l�nܛ�8a��Q�7��Jxrs!u8�7�E�f���&r�|"I9t�j�ޗ�&Y��P�_����E��w�a���4\�8$�u��򉢘��_{�t��c�ţ����\6�V&~[�$E�᎖2?z'�1��ejQ����3I.q�ܠ���ؘ ���x\�J�zpP��`t�D��UD�a7|��P`��z�V�ԕ�Ȯa';;�!�oی���V$�Ҵ�X����u���ty�A��1J�ɠ%���O��q��w�������_4�ܜ&���i��[�!4wٟm�p�W]�~����i�m׏0&�1�n[����~5�mYf؛�TFJ��2n35hg��ꇐ갶�:��&�Ec��;��r��L#�@连��Ӱ�n>��5�(_�n.�L��M�Xr���P�q� ��s�zH������=s��:#������ ����:=���Q@A]#��=6~m��kn(⽽KDdScd���\�>쇃A=w����'��� z�Ƽ�����������f��;K���?����|��p5�o��>^�ޭ�+!�ԭf��(�o�bYX��ς���e��<�1���r5�{1y
U��,1�~;�V�	�٣/�����.@0ߠƎc��H�3��r@\w�}��^�A��ho�m��gl�!d���%�W�N�E��3��#��
�;1��f^E��_�]Q�C ��Y�J�Ǚ���ZӃ!��#c��e*�LI�g�u�.F]ۂ;f9���4z��@��3;�PJ��Y>��N��cu�E(�Zu�����n��}�G�?����"���y�6�Sz*X/����CUE��y�L��_�����}c��IˎAt�*/�)���}�ԭ���m��B ,`���BM��*���w� �!�Ai�㏙[=��^���Y7&t'O�%�1�Dl?�]DH��K�y�o�|[�e��~|*3US��������]�m��+�֚t����$���T�ր����5���فGz��,�&S"%><�/F���&oԌ�q>���������9�]�&TV}�&�V҉aQH�8h�[3��2<��_�w�Q�"z��p�s9�hPN��!4Q���v���á��uS��]��ȼc� �- '��0z����e�H?q�_��F��허ϴS� ��^H�c�=�����[׃'���f��ކ|���H��=�3`�����z)L��t�*/=D;�<ָ�W�{�IX�c���5T�Qnzq��\9��V�@�xO@����a�ip��Nδ��Iv��\����D-��0X��Y ��}�
�5�]1r�|tB9,�B)��+a�>�5��<f���}V�0�]�C�+��x#S����tN�GDdj�r�u&���_�I�؍���Wf�h}7!5�~w�A"��~��ᑡf�9�@��7T�&���^z���RJL��_KÎv8����+�#]�-�/�k�x+Yg�\�W�}��Tf�����:��m%���Q��zZ��?gEc3wa`qP��ɍP&�/��(lq����Y�Z9w|� ww��֜�ֳ/!B ~�$n%��a��Yꂸ��]fk�x{��$?�F�m
]�Y�����4�Q�<n�I�x��F�����F>ku��d���/�u�8�)�B4��5
��УW�2����⫤}�*��wuX& ��vH����`�|e����ك죔te��|#���rU��1*fO���^�����W'���>F��m����R����$�*7kC��wS�.I`t�I���a�,}�x���k6��K�	��V�>U�\kγ*���s�$T��sI��-d��v�I�3���8{�*�]R'�S̗��^�KB�!��6�]ڬ��	3�fzؙ$�W�!�z��q�M�����QT{�}tv��J俏տ�ˍ�=4�;�t����lՎ���}�BZ�&Xp�r�=��L��<w,�TZ�^CI���.���  ѯd���'�=oX>����
�-R6���Z����gR�2�ǳ��Ц��m�)%J(nq�2�l�� Z2r)�L�3���bD�'��+`�8O�� �IV�=C��V���Oyno��g%�E��b-t�X2�}LT�PL������k��W)�#ƍ�!������E5�؏pV^�<�=ڼmG�l���͊S�aTzJSb�YCa�f�t�Mc����^�x[I�0�hz�^�� 
,e�텏��Q���
蜉V�$\��P��7h�K�D��>62з]tK�)R�Z��^x'�����>ٽ>���u�-���������T1�F��'e҈{d��9���M����D�zTdv8���R�;�vnd��Y�H{d�r�C�j�x���S�lD޷Kb��r��!��*8��N�����P_k��=�+r��_�ߤ���(�i%��Ϩi��s�`� �K��C!��{C�����{���!_�ܙ��\��7W�Htr_�����!�"o�6x�!j��(��K)�o��)�)~������L3�04�qw������beO
�^u{L.}�Β�d��S9Lfۻ-���SHD�~Y�Z��M��O	,Ű�8-���= �����_w�Z�J(>?����G�Q�_],���4�R��T�JJ�������ɪb7��ؤ�c;�ם5S6�l=g����t�H�������bY��}kB^�'�jT!)�3����o��=�W:�M��e_-S?��e�>�vd�� �il��u7�F���K����l��Ia��JuL���x���������>�qo�/�> �{��Pֽ`2��(�mJ��iq� �LFBi����?��O&�~'-����;�բ���TƖ3�-cS��\�`�C��|w��1��
�~Q|�,*���.���NL����'IV��L����5�Z98���}{%b�p�	p����c*�=^ȇ�J�t"�7֊đ�O�8�!l
������*?�$����X�|�!=;��J�H�t��A��%oCE�h���}��n�-�k�љ ت`���� Y�X�xY�D�)��@�n�Zn���I���Z���)�x[B�ǝ5:�m�ɴ%�mε;�Zę�U.�E�b��XxѺi�,�"`�K�/��w���M���r�o"� �Z�Z+^���A
������C�Q@Qz񌔛����t7��]�	��x�f���B$�08����3&�ɤׇ�Q	1���j��<j8[K����]Q��F�d6k�2�f��[�>m=F��8cQ¥R)�<;�7��ɐBd���Z�K��ZI�'�ٔ$�;�j5�����F-⢽#�Ϥ�F��4>�ДfH����O�.�j����ժk3�r*f���ko`n������3U�'/Z�-,����!ܞ�G�a���v���W ����PP��45. �M�>^�\#c���S|�x����/�tR0IRL_U��!�7�-F�i�C)��/˸q��'���43��誢;(*0���a��]�*L��M� �;>s�Ϳv�?�!Ɗ�l9�[%�q*ۨ��g{�@������8-T��$N`Ki��䀯nz&pD��	Em�K�j�"}WD�l����sڙ���P���.<B�a;<)EL�l��j����:�?�<�f6�8}ꮩ1�GF���Lƫ�*}^U&�O���K�D�y�P�Ɏ{��	��q؟]5y�2����<+X��Jں��%0��K��)��)��ĐC��S>R�q�t�݇la�ӻY�u�Ͳ:�bu5}�w��IX�{�<��ɡI���l�����
��K#z#y���̹a�,e�M� �ч�7eTXw,=rW�=�mt�	�7�e	��!`$:̿�U��_F	�Q$�Gd�-��C���r�#�4<��} �f�W�Y{�s�����K�z��W�/�B�*��-�({'��Z��>�]@ލ�!D?qaS�jwe5���D�R��sѱL#C
���!���Pz��ƽ8�_䢦�L��H`�oDG�t��")�8��-����\�;)�)������2�>Ҩ}z$C,z��j�:��vr:���o�/�4ڮp��ݑ\fP�_��$�9�e����D��y���5lr�N���@#������jL,�W�CA|�=�=7_%�J�#f�UcT�!#��HyJ��n�${~�={��F����q< Øv,H/�*.�ג�.Pwq^6���SS���f�~���Rcr��:�(�x��#��z�`M������˗:g�D�ş�_��h��69d�h�b��f�<��yVp���u����ˏSU]У�<�j��(wo����&�\�,�M"��4T�$��6Г�q��s���!	i�`���5�E���m����^�ňpM��b�X��
qm�8�H�t�'|�?@�^`�9">B��z>z
R7��k��l&�4-�	L"�,ʆ�]n������F�.�_��m��c�g�O���ԏ���\aHz7vFF ���v��fh��qn>��Qr���cԨ'u������d��{���W��X�"f��X���&�����cĠ��
	��۫>���YC�a�(wV,����7Re8B�� �&����'m�4�/���M�n�8�O�s�",_�L� ﴀ+}V��OÒ�dG�ID������N�Ԏ�;;��FIz��Vd�`Xy2�(�N���,:jE�5>)�Q���X��*i��'A��4~�Xn;2>)I+"A��?����9_=N�ih���i��D�1��X��Ȼ4���2��W���Y�s���������� �&S���[^O�
����5'�x�k��OX�~�m;N��V�)2S���t���_e��^�*�(��r�>"�dS-�6��:`ϙP���{J���Fp��'΀׮�Qj$W�}gQ,�.L�`��,�!�n&t94�68+�����g!
ۼ�M�\:�&U�����{۸c������&p1��I�P�eHϦ�m6�X������7�jt���T�>����~��d}a�U�w�8��я��m</�r4�n�����z�$�r=�fG�;F������J@�T'U7]�(���,0+��/�j}8`�g�
aΕ\��h�/��ńXw�)]>��$�$	�v�	PF�-/<?�G��^�މ��g�K=��h.ϫLt�� Q��|+�O扣�q��#�x��5���D�-	U}��f�5H�����:�i&~�MOn��a�@���Wn��x��l��BAM��]�k-�W\0�NJ�W��Zm�f�J	8˺�{����xdm=��}�I٩��VMJ�*�N	�0����&�K8u��[ysO�*���3��`�Zq�/v04D4\��x��GҡV�g8T�{�u? �Co?Zޏ{X�d��g!�^J���z�3`&z}&+�%��s�]����BD���eNsL�s���:�pǮNÁiUA7s���%�5�!!9 ���R�O��f�9�A2N0I�Q�&��o�P���K��'��|�(&P��-��cozT�kf��@��?詎�ke�f�G�ԑE�d/���XM��$	��Y���X�8�yg��>����������F��
~�Hނ��<��|v��|�o��^p��	X���A�H�M� 
oa��t��@hs���d	�\'Lc�{����L��0���p�,'1"3n���G�C��f��,3a 
hޗ����l�ͯ��\x�G����[��@o\ޔ�}��q���e8ͥ~M\����Y~�4i'���:����.ECc��-`��B�i?����̓(���ݾ���)�̿�h穩z��~q��7>
�P�è�e-z!��9�T�]��D�9 dZ��RN�{�ҋ�����H	�q����8a�.<H���A�v9��^շ��~�K6��9�G�E��S�\�{�������~1����H��S��v7U�� ��"L���i�N/讽�c��<B�z�y����:�n�>�*����2�?� L@��_�Y�.���ǆ3ʘ� �UD�Ӡ�����㑖���p�&�1d��if�x�3��̜���\L6����BjWV�YV�M���2D:�˧����0gF�%@[�4Z��T�#
����r�x��,��0R�<E"�"H�� Ol���V�![1$��޲�}i;�$7�/VlK�ܵ9��
@M�U�l�����k$x
���c�?�G4��٪[��4Q5{!|���m���8��(�A���(�dVU^Ă������j��cȇ�SQ��J��}���� ��C�*,�A������-h��/�d��ʍ\����C��f'������F�7!����`.�aG`�0�[����-[�	���O�4���d{}h��m���^�E?x}��e��2��o�#�e���DED�5*�љ��M@���zk:�
���\�����?zU!���ǋ �m,�a#`z�w*�\�/�d�x�S���AY��#�=}A徲m<�jW4b�Q-k�@�`��~Ԃ+=�%Z�<i�])&@��ub'���q9��=���/e#���fS�%Z
��AM�IR����ao(�7"���6��s	,�'m}dhq6�)�g���[vVa�"��/�Xt�?RFtX4�hV�0:#(�SQ�����W0k��q�L[b� ~���@g$�p���<!�s�XѶ�TWr�-��S6�.[��Q��ƌ�nEh�}1"�1�5�P����_*�������ox��*L��-����Gx�zq,���e.�^0 ٍrL�����1�/�vx[�nk��J�ã�FQ�$�g�w������f���ޠrh����v m.�3����-��я)NA�@/��p�wP���|f��}�GwV��e��O9ա�I$�{�S�H�*�ٚ.�S�('2���w5���% x���:Q���|P
$��~�}����6�\T�o�y��wzIH�Q^�D?�@Ǣϛ0c�P8D��>_J�U$��%~S7sH����,�C���.tV�ƌv�]�4G�̌b
P�9��2�,�O�A��B\�U���h	jsܗ��1g�@�?H�Y�R����BQ��x�C_ehi����od�*C,�!ݮe�⻊��.����c�X֋'��s��gy�s̻}C�.\�On��,LL�]veN��PhQ�����#�H|�{��0?w�T���`�!?�`�07xU`�F��L��طcw��ST]@�*.���D�)�u=�ϕ6���/&D���R��0����A� �,�]Xsb�6G�G%��.��6'��u��uA6:#�?��?�k>*0&�!�,tO	M�3��6 3V܆�4�IAg���`�n4^��a�7$�m�+>�!b��4��݅~H�Z��9Š��/�
��
��a�U��3�]�F��vē�1�aVŊ2we�Ƌ�2?�p?��͞Us���B\
���q{�N�w��B1/Gc2Ӥ�ꄜJ��~�Z͇�v��e�i$"Â4�h����F�^�L�p�q�Gz���9��m��& X�{�~7��:�>�ʞ�cΫ>t��$x��69)����,�^�v�^��@m
𓿀�k"$����D^8�l<�ʽ�>�^@\�"��Q9`��J��o].��%j���n>G����P�Ӹ�i��C�R��o-��	mRr�Ѣ�̈��vxrޚo�O�q�Q�7�c��֗�ppҽ��@*�J���Ҹ�_�ֱ�t�1�vI���&0�?ʡ{�c��4I��ʞ0����~�(̏T��Ц�[X�ݱ��f��M-�������riVsTx�77QJƼE�\����f��f��>� $g�ϰ���:�?�A9ɻi[/�0���Qy(q**9��C���g����<����=b��i{oy�emj�b�D��Η!�U�����=7z4i���P�|dFP;�%I�U�[�<T'k7Н*N2�t�6�d�\@��/�j��/��&��^�⸰�؂�w:M��[�j3�q�%U����v���6�Qḗ(��)���1�S&�6����r\�m���)�^�7�Lca�Cat�;���qb�"�?�ce��Y&w�,���\3o=&�AD1Tέ�~ˌ���r��Q96���O5I�FDCSֹ*,�~'͢�U�0n��� E�Mg\;�KU������E�ݤM,w�U�0>D���"�Ń��{a'i������)�zB��uPbb��b&�S~�R!Ic������b1ވ�`�B][˦���=�!����2,t�}Xf�����!J��7�lu9����+�@s�$ov=RD���.�Mj�x����Bv�B&�l:�sy�V��O.��8Jhw&bF���~��B;�����{v��O�IԘ=��!���@NJ�eZH�?�����{M}<�%��2��s���#U�$ձ��^+���ן��3�8�,$�m�D!�z�ij����8[4"0h���|G��> �$s��2h�� W·cy��"�(��r&d�;�Қ�Ѝ8�F�p��8o�Nh��Yq�b93Y@�~�1���@g[ei7�
�WMf�o,|�S�����8�@ �%µ�붘�m��&A^��P ����_�/�s���j��\n��f+̐�oL i&��灟*Y<X�����imA�ȔdF�'�c�޻�Tp��F& ��|#0�>���|�|%�� ��&G��5̊�.C�wT�B ��^�Eb�~�L��d�a��X��7�qQR���(�o�/�n�)/<�h���N�J�R���<����3��?��"S����g��Ps[�Ch+��H��ӞV���=W�4�[����{�����S8kUGQ��vꉾ����6�%�1O�&+���Wë"��F,r����Xd��=���k�2�!���N
��A�k��ڀ�9�6!k�=�p�*�����wO�Tv��&҈I���v��7��Q~>Ӿ����j�R�.�B��ٮ���H4�_L���BbGD:}ZW~���I�eJ[�����<F��f+��v��@�u"? �G)�������0x���U�N�*D� T��w��][_5��v�Q�d`��$�B���N�N!��)���G�<Ӹgr�#H(��T�8��Z���|l�P�H���^!��ʋ���9�]��
<�^� ��a�Бz��-Rn$���x�5"��ӯ�ĸ�u!�f���"JY>����JԻ���5���_��ZN�X�7/���j5�ҕLoW�E֍��8@�#X�����
����p�Љ��(v�d2$Wk�N�-�e��A�*�e�5ڕ�
�0`�	D��.$��|�����O� ;:���ɈT 6��Zx�+H�B/��g�\	�k\)�:N�Z����=P0�;�
I��H�;d� [=L(*eǙP���N�Q�L����otK�{��y=��D�pu���~�����Zǫ�Qz-!�:�jz����\/��D)r��)g��3g��E��7�Jp8��Ǉ!i����b�=��S�l�X·�����5�+Ԥ��jN�Ҳ<�O����"��q�%3�����G�;]�J.5ԃ� _�iW�_�o���n���<ۤ��ѫ��n���ތY��Y����D_�����;��.�xv�,���7��|���ZT�-d7Y��hv�m�����]���C5G ���ԙ̰w�BJƨV��a��`w�B:口�a�Z�����w784#4�a�����3�ίq�fڢ��٤HA��f�qMR�R-��8�uq���z�6���[m-;��g��A"4L�˂]x_��s�U�(��3�8M�8L���jxt85~��QƤ��^f�>��_vY,��b��*Х8ev��D��튊�!dګ�A�^��+�Xl�$l�_�zB!�)k�d$E��)����N�DE�[� d�?~��+�v��5pT����y=с��	��zxca����+����$�2��63���n��� ���9�GƗ��_�C[���P͐�#�E�X_"b�t2�@��
�m��i[�rS8�5/��wH`T[��jB��ri�������-�\s�;�jimQ�N^?\�!����`G2<�� ���Y舑P�W��fz؜ �x�3���u��k�����_�Y0:,�egy�G��^�4a#$<����PV&{3F����X���r���JY�ƣ5i�������[qY�M���Z&V��)�bMc�}�<��};���n� �*a�FJ�kD�z���`���QM�	�����=�{���V��m��}c����UtO5��	�����(�LpJ�KRQ����dp#<j
͙����M	��Р�6���6�e�D���8B2�+m�|�������o~"�i�U��6G.4�!M";1�fgD�.�eLp셆��ƛ0Z',,�'_?�C>)�<��G�pJ8�"W�|FE�S-{k��cu�򋉽	��T"1�i�������fc�1�G�~V��`"���}{����rq#�HN��>�6�ٖ1��W��d "l�tG.�k�O,��,�6 δ;�jO��~s�Zf�x��f�R�4{�cQ/�Au�� ,](c<�l{$|�Ҫ�����1<�����L��sD��>�?����U	��"�# ��F��F]G��I���U�f:��+���y��܍9˱lHS{�x�G&�HTDWy����Ж�c��w�/O/��E��H�k lhB�>����E�<�6	�C��@��YXJ��	;4�k_!��B���ܑ�u)-�ζ�\����BO�M䙣=^�����/�EC�F�R���\��y��Y"5O4���S
f0R�Q,� �d;�J��-�O����Y5�b4#=�TZ�@76�:9NisPs����3�&ƿvA?��^�Q���?&]�� ���p�� �S�u{�K��[O��B4�w&��:�C�W:��o����`��+�ZW���)V#����r~�n�A���6q˺����#@!B)��4�'��{�n�����s2+�*��ԿR�m~���~̒�%',�)9�J�R1��u<UM��$>Gы�b���L�=97���Z�.b��]zf��+Q��o���(!7����2�I�f:�mab6�7?��L㼥
bk�[U݄+����G���7i�Xtz��dA-l��(=b*��8��0Ɂ���x���?��^1����zF��	&�����W;�T]���
��C��	������or����
�%1V�����[Dv�%�B�Q�	��.�=�N�¥C���-��
mǟN����+�j"/�כ'bEθk|{?'M獸���ۏ���+�+�����n3�-��~�p�Q+7@ί�甂���Ag��wh #i��T��ʀ�5߱4�-����Qɻ�ܓ�)��s�� v�,�<��˟��f`Q��򖛒����	��a�CG�YԺes�x��掏i��۠�k,��q�*gX:����G��ƿg�~e��)$�1ќ�gOA�Յ�4���I��8�9����H�-P�â���8
���Y�s�O��̵�nŬ-������R�hǖ�}u��#��t���P�� �id̢��-H�h��H<��"4fm{���
��s��dU���	�	W\|�
7��1���3�I ��fW	�{לiM("c�(�2[�S�d��S�uA�F������rnX翢=]{����������p.k^4v�=1M�kk}����n����<X�3�Ь9(���L��>B�\�jV�1Rk�|C�O�ѐ�u��H���>�ې��U�RR_cc$.�$`;��-\�d|
Aϼ�M|sG�DC�;������������N���5|@�M�d��J����يʎ��. ����^�����u.��B�ܟ 0���f�S$䷤Ⱦ�9��,��)��Z�L�G�nj�7b	����(fip!A��3Z�7��\��]��,�-̖�Ko9���Wd���BG�r�Y9A���O�B���lf��G�d�od�����KBW�@�?��U@�d�������D��5W���ޜo�yL!`�b�����E��w�1:�f���_����#��P�Rdo�)P����r>oٱ��C�X~��wQ�����և��7�8��iĠK�e���
�4��r��e���ohRG݀�3G_
�o.7��]��9�����l��U�\z�XiE~�8p��������+7���1Wp�*h�^�\���^�f&�A�Y�m�Q����ʁ����H��s[]wy�'���8�s��|�ҷ�$/�����GC��	�#�W�'-� v��PE|q|^HX\®�:���������=v�N�T� ��ݬ����9Iі;�:�E�(��mPc�LY���!�d{�Q�>[���桠A�8���G�(�g�O�h���q���Q�G�f��R���G�<^���RFhq Ws"u��8��㻥��_%;<����������|l�U�!X=�Wc�K�{���Gt1�8LKo�|x�U#�}ug�cނ�_�۽ �ޤ��Ư	�v�a��%�<�XZ�������j9�����,�������fC\A�K��K�R�I�0G��Y�Iț~��Ha�'�Y���/g^���7�	6��\9��)�TLW��h���$��0���U������5ք�I~��m�?��FK1ּ��[F��[��������O�Aҍ!�����!�	��,n��Q�}������<|Y$K}-z�c)�����Ȁ<����n�F�?>��0��_��\��2o�Yx��?�q���^����O����ρm��	���R2-��Ua��������ü_�c�9}٘��zL��?�F����Ǽ}60E�n��~��-�	;l�R��i����!0�gWW RC�%���U�ջ�^ct���8�T��u���?E���|\o̖�+�&�*��~$�"�m����ux1�U,��f�����wr��b�1��A�NL��L�b�'��9���Ȧ�d5���6��5ޔ����#Y5�<�Db@s�ӛW����Ey� ��F�j��<Dy<�R'ɷC� p(��ӁvX�
��Y�ǹ2@|�c!!?ן[2��&�Q˘�w�;�O�PFqH�W�fl?oV���F�$���q��ہ=@�Ig�	��g�3�l/�H��������k��P�Iƀ:�!��7H����o˨ ?��#��rlh���
��t#�I6>T��Q=���w��%�3���j�`HU��g�he���:��\�y�.���:Fk2��Rua��:�PΣ8��pM5="V�Q�q�|6m�ӭ��o�$1������!�EI�	#1@-��ϋ��w��X�*q����mY�M�c.��	�]j�{��6���aL�H�k�
Q���m".� �+y&�ij�y,8��I���\ �fj��+o�DiTU7+�iG��4!������l�������#����^L�������e~���IǶ����@'�O���^�et�<����[�Ԝ[`���.��7hMa��w�}/{4ihd�O����&�jOQ�=z@�e�)����ˣNw���
ۅT$|���7��ҍ�T��G��?v�'t<谺}�2�<��ҩN��@*�-�u;��n�0���R��jW�&�e�D'��V�Br��2�n�6���a��9��vI�ƌ?��P%����'�8D��>�m���'wV��R�F���bVކ� �g�@DW���'}{@�)�y~zϋM�[vp��I`H��cq*D��b�&L�kX����1)�������v����X��3��~������C2h�M���]����Y-Si���I����]}�9�3�Kܣw}�.�Y��v��eK'M%�R�{���3u��R�"&f���C��'J��A9�5l�t�?�|��������Ig�9���� z�{S�?��K\T�����æ��9�q��?�Q:�.Z�����4'G,��K��b���NUlQ�N��S���T�_�B�X�Q�PqD���s jp�Q�N|���f����NO%_}>�ۆO�fF܍@�DsI��akv0�j�M��D3.P�,z�͓�𜷢�1"f;�X�r�Ȣ���xgW=�֛D�I�\ &���;]4�!^��Y0|�%n�抒�I� :GE>�U)f� ��5�"&������ �����@�<�v���r����L�2+�>����+��O��D�tvT���Gqǽi�F{�,����'��E��o�D�
+W��ў�WG'�j��~�A!Jh�U6�#�e�Gt���Lڙ��gJ�j�D\�C��%W�A�*C����u���g�b��'H�r"����q����i/�.��!�}�+R"�*�O��������ࡿ[^��W�H��:V�k����@��I�e�k��\��N���Q��J��r�~��kC)yj#tk�g>�S�-ȭzoy{�b��`4
�?�#Q�N�
Zw��%�o �w���C���f
BCb��H<� �
�%-?�qRz�k=q�z.'qe_�2����|�a�Ԋ&�tI1��*m}��@����O���M�Bu;�A�J��I�������+�	h��x}����P�Q�X���7o�F��\>9�#��&��R�=%;����8����2�NV� �HC�o�B��g5���9;��V!(w�����t���3�6��͎tØ�[�d)v�9�;�oe(��s%ܾ3����p�X	�Cj�|A�i���7��FU��^�[�k當�DuC���M"�jC���#�Z��<k{��ȆO��9f���Ի�����z�7x��|�o��|b��J*t?ƛ�c�fi�%3�%d�.�^�gk�7Di��^��s���I%���D��[�+����N'[$��%!O	�=N�f�Zʺ=��%��S�v���h#�ڊ�v3k�꯼��w���e��2��t�j����ל+K��[2=����}g��>.m�,ڴ���*�F~>�y۸��m����'δ��`��U�x1�h%���|K:�)��T��u��'�_j���ؽer;O�;���U�;��3���!A���A:&��M������gE
{�VG�������ܷ<.��a1c�'��c2��XŢY�C�,-��b7�f�Y,Aǳg2����%V�߶�er�ڟk���bhXK#ML��m�%/U�� o�9N��*cra�Qˏ�ix�m
�s��ћ`��԰�\�B)�)��$�5I��*�E=��5�S����/U�e�5&��<����M"BEZ��v����~��UeL���}��r~)�DBT�W�vb�I<!QKS���"N�L-!=$T���9�/k���lnt���V$A}��]K���S��}Q�y��<8��g���.�߷�[��++�#E�Ԛ��+ʰ�K�K�Q�w��X)���w
s�{�&Pd�-�}��s��#Z�5�A��v�۝VN_��P�Ͱ y�m,?a뾲q��'�k��A=J�y��SJ��t&�W?r��E:�K��E�n��/��3-:)���|z�wU�/�Q8tN�4g��?L�mE���h���k�R=�\w��g�N���z;q���f*we6���M��-�xHt/o�T��9�aX9���C����C��c7�ZM�n+��3�Ľ�bB���U�;��8Q>=��)�y��䡍o��}��i �[4l��-��ѣ�f����I_*E� *�l��	K^2g%Rdg�\a>`tD��ܨPw�B<�stc��`�����<H�ox���qr+��G�?�1,KH�e�K����P�
�(���g�l��h�� ���'Fx�8I*	�EC�hnAd�ʺ�s-��~�Mz��W�FV���k��M0��V�E���w8����^�qf%����!E�P[&<9a!L̼�85�5K�N(���n��Q�����O �̔1q�����m�lS�}�؊�N}�C����0��tb�ѿై��b����pö'�E�����q%�k ���B����EdŸAq�.;p<?��W>��Q��W��ް=<�2���2b�_iWM�ЗL����hٔ�E�9�A[�!%��S�/�x�J���n*Z��*�ˢ�}�NK2g���0#��<�e72����H��
�ɨ:k� X�f<��6�e��u'��y�?X�|O�g}8*�{�08�f���o{XIg�⡁y��ϩ�&�RpVG�Mm����*����s�e�A>�#`L����k�8�ƳF�c���<3�^�CPdS|� �QV6����PP׆�<h��U�3��G�g؎Dy�K��ކI�c���)l�zI �S[}���uL�W����^4(�8�"M"�,b^B�!5��&+t�1fb��J��h����$�?�S��6
X�̦·�y�w�EӺBt�˶V�[��/���'%���^/9S���T�I"%Q�o�U �ɡ��
<����d{)ז��%��͓F�q�|�i������|��|&� ���_:��
� M&� �����@�����Dm^)�/[}Rڌ�7��YL�%�I��6�^�ٿV�JS�Uϧ;�i�Ui,�{SJ4g�%�9��F[m~Qc`�t`�������Y�ɏ}dWCc��T�T
�Y�>�z\�2��L@��~n�ʾئ���_္��nE�5���������e�=��*�Ns�K��8窟pJ�A~��JTu��~��:t�V�_!�J�i��DΛ���}8}0�@j��gt���׹��3 ķ���ە�䢺6x�~j��,���Rk_?��l��-�� ���Xg��Ja	�������N��+Z)�q���<�)�3��Q�	��J�������K��c�W>�_�G���5:���d��g��1�E�!=���h� 3z��$8ڡ�M'����v)'2k��~Ճ��cT�����P��ڄ�6Jf-r@�5	���(����qX�z�W������FP��./�L���l�W�$�9�����Od6��^�Z��[q�tD��1�,�#�b>p;cyz*C�xU���j
�;iL�?u��B�ǣ0=��28�:5Ō�ڗ �G�^ǋC5p��CC��=!���Fw���/M�oz�6p���4��*��x��Rn��-���k�%Ϲ6 w&�sD��U�ܾ��2t�;>,1ݳ�BiЖ#�^��ɲ~2��O]zJ�Ld=�eJ��ս���r�R�nn�Kq�YN.�G���RT+.%�T�F��o�9u/�k<����c�0̿a��D;�2¨��d�D��?|���=���=�`!Ψ�jW�Eq>U�>��/e�R��Z�!E�I��F�8�#�h����L[���(��8�̥���������Q�2��x��
R��n>�sNTޡ7��ٮ)���y�~[J7�RxDTܺk��\Kݺ=rC�i��:�/6ed2h��$W�!_(���U�xGG�+O	���+jMJ�n��N+KaL�ʷ@C'���#�
�YE�(L��OqẼ5��&s�*�x˾V�5��	(��J͇�p�f�&���d�s3z}a_��zLr�����I0 �
V���P��x�[�5���%��^���ZO-�>*e��R?[?���h��(�0iMme-Y:5�0�N����&�lt`d C7A�u!����57/�a�ho���n.���!�(5��'q�f|�J���Я�!�����{�[������Urny��sc�
6[_�:�m�qV`x ����]��rA���\�"{�c�omsY`$��uǶ�)�k7�{2ۻ�J��=�� �2M��l�420T�t����ط���40�/m���ɂa�
T���Aa���8L���p����ό
@w��j�eQ��`�\F�$s��E�����5�8��3�."�!����a���3U��O�iSi�j,Do�Z*P���Z��2�J\3j���5Vl��ŮT��5=�٤-.!����l�X�_'tlc1��8q�����I����A���a.b�-~�j~j* ʬC\n+~���!�B;#[���L�Pfi.OS�)�y�Mv����o0 -l�'X%�A��g��u?�2U
̌���3	��KOf���4��~b�	�H��y7Fl!t$��ԕ�� �\:��Pa�����c��X����i�y޻}�3���~b���w�uF.7� ������;�vt��y�Gr�z��N�H:B C�5�Ҡ��v����m��.�Oy�
l�z�n�:#��)�#�d�Re����=<��_X4��t�j5���xJE'�z��v�t���Α���'�'M&#%�*wj���<[�o�34h��E�5��rYP�P�o�9Ru[H��a���Z��;��`ҷ"����j��SG�H��R�����4S ��ee�c1a�{��1<�:QgQk����`w��-{��EF���T��l�!gɻ�Q�8'�u�x����,C�zf+" ���Rù.	�J�zJC���@�Co�U�"Ӥ�°l�d�J��ĥ�UD0.�g�q�c/X�g�Nx�9F���'�¬�Z�$;eq FV�T�o����X��tmn�����U��¨�%���5���~�-m`3䇣������ ��A�دM�u�<�j��N��g���?��?I��}�j~��x��" B�IQ���%�q�`�l��a�N�|у����0K�x��_!C�S2.>��k�?���bj�?4�{o�f;<F���t�i]��T�"A�v��,�0}�[���GM�3>a��B�q���j,��XK��p��FBi�{����t�rY<�]p����\�z!�O�5){[P�c��}l׬�!���(�_ c2�"8�^!�s�)�/��g��f�y��W�p�ς��7aU��QDw1 �q/u��h<o�����J@�����a`o��g8iCf���A'RC��>dL2�r#3�dY�m�����%#���'&�A?�x���J��\]���-��|���3PlAz��MN���}�J�%$���1n���q�����3��@Yt��:��
�${�4��Ӝ�(f��$��6�հ���t�FZZ�qMlOGG|O�T ?N�?9��H�ѡ0M�W�@5U��o�!��'����=Y�n���u���K��{ X�����:W�P{؝tL�g�� �,�D��	b]G"#�f�9MG�����{~5X!]�I:�M1$y�n��;��Jy.��A��~h	����	��$���ç�a�8��Llnj�9�f1���7'�O3�� �|�L�ajюgG��[`)Z�9T3�����P1��u�F�#� H������&f8t yE.�^�M�l��g��1�%�؎�j��^�d̶���"o��˶��cV���_���Dg�3]Dl�X=��H��¹1�d��8���f��]CG�?��3��7�2��{�ׯ���!}�v��څ�6����k�KY�6�K�l~
�/f,Y���s�"����`-�3�VW�I�Z"Xm.AW(�W#*���B}�o�������p��6w����/mWo�)w�)(��@�H���M����uƇ�94���h�}�����N���/FkMs�S"ޮ�o��6�,9� �6*�
�_�1�Z
��m�Y���3����&p���F�D��o�p���P�@���Vskp21\�������N�	 �q�{h2&}�1��c���סky/��7�5$��i>�V������Eq)�}p,�d�v�׸�5h�F͊y�.pI�c�N2�7Z�w�l�Fx���U��]b#�	��G�$��Mڰ�J;���ll�����u��:{8�$�N��ۈ~����f!��:Z[z��h�Y%ݰh�'lM�Ĝk��z�9�?��qN�v�5�:���U,.���{�'�p#C�;��<�؏���1��4E�NU��=���ث��|4{,ɾ�Yz�Q� �l�,��97�ض:�>����ٽv����I��H�ī��� l���o^=���D��S���r���Y��6qEZ�S^Er&���hHt;�R6����0vM�=E9�ŏ����� D����b,AXq|fa����{L��e�ީ�Jv�p*I#�GG���'���ʹ\r�t�⳯�j�����m�.�&�'j0D%y4�[�yR�:��`Aǭ�>й0d�jZ�H%�}�*���[�RS��;��xs*^�ߤu(��G9g�e�\t�6p�&_�fv��M�H\u�6�����EP����)��o�@�` <�+#h��]��9���/�OP�`�,�b��^51$�>P�p���B��N�����2�� �K��L��ŜE�i����&��:p~����&3ߣ}���"|z��DJ��Z6�M ��������a7���2f>g�v�ޱuZ��mVl�*���˴��%}\��jz1������=��y�H'��
q\��V�߼��B<3��ϼş��(�J����Q��\'�����qe�ߥ=��eW��(�ʌ��H)JC(>B������Z�R�"2E?`grm���ز���=�;h_�%�����lOf3]�:�&�����s�����������mkR9��dh񙠏EA^ڸlU�~�r0�蔵���t�_�)zӑ�\{�ᙐ(Ə~��|S�j���6ve�" �o�A��3�g�_ppg���ޅ�EY����L��N��_Y�?a�A�$<�}�?ݏS�_�֛|��^I���/<$�G�*#��� �E^��+:���cӬn� �v�i�u.���eVs�#���;G&lMs2��ʗ��Z3���}����-����+�ڞ��L5c�!�+h �胰�����O�2�����4x�,�2�A5O�w:���tO���yj�d��?�����&\�b�2Λ:�
�!=��e6\�Ý^�K�ȵ5��
L�'�P8����Wo�8��w��������Jsb��dP.�O!�b,M8u�p�g��L_f��p��yd'r�/R6N`YŘ��#����DP��ت���,4Ì�T!�e����V���D�A8(���vh�0�9/5Q�܇P���)m��q�W��e�G����c�[��NA�Pb�������ڽ�q�V"��n8�|=v���%p3|�W �����y�!S��K�́T0�5�i��2�G`w_r��������ʠ\�f2�S%����f��shW�~��"w������lێo��i�X`�RR� o�0��|"VD�oS^��'�1+ʘ�W��M�@LF|���xe��^]s�ƶqe�����:�'�\-s�Kx;(	����~!��Oo-� 3R6:�GZ6�n���6��s;�=��j���Ҧ%|�	�gN���]1_C��4{��b/QnCcϷ���,̀"`�� 1�n;�+N,	��j��+�5�����U�[r�0�Y�ʆ�1�uʯB .�V�+��﷨mi�} ^�]o���!tTn'����ɒ��^ۄ���Xd���R��Qx���Mj���%<�zk���~�@�Z��lkx���f�s{�z й�I芲?�w�ɣ�e��a�vt�)<N��z���9��?䝎�!� ����V�.�'F����x��^JvΫ��ـ�@�k�G5'e� �-�왛���c'
VU��F��8�W#�� \mъ���C�幼� '�x/�|,��&���߃�}ؒ,F�̈́,6�_�iw]>�r,���\W[a���$g�#s���Y_����!�Ξ�4�*1�J�W�V����鍧VDr�BȎ�eU޹͏6e� ���n��T��K���4/!c�:Y���U��M|$=�-'9^�	̦u̼�ke�a	3'd�,�[��,H�qл��O��l�dt��?쬋wCO������8�i��ٽ��+=�/��Ȏs`驟𩲔�ˏ�l�fb����iP�C2j�`����]��k��"���,�8^�'+3+EW�����'�-���G�H�q,����s6�{����B�	�+DYCٽ�>�m���*Tv����D����\���Tӫ��	n�3�0���@�9d|s�ͽ׀\��e����p�]�KylľI4�<�ڌ��|���j�z�&Q#u�mu_g�����Q3�X�x����J��g;�����ήQS�,f;"��N>`o�Mm1x�(WL.6�.����t����4h�<C�o��P�.	��*۪`TG����4ԝ���T5$zoK��4���#u��&����û���_2#��.���^�.�X%��(�E��3���~�hו�ʄRõ��a�c���@�Q~o���μ�SUp��4���BJw����[����4d���Y���Y�\���������%+�Y�X6drR��H�ra��|؉m�9i���_p���`���:G�3��ϵ��*�o�%P�ڝ�S�q�E~]�j�_-X���������9/�%n��x�x&�Cd��ꄕ0#3Yj�d�������Z�!E�>�'�F�:T��QM��3���L��^��y��4NJ	�/���f�{��;�z��Nk#�t3��ETM[��c{��>1�.��o�NN��v�Hg��(�;��߭�n紩F�v=k���[�p����	���<��jٹe1�:A����i���=W~����� ����kP���I�tfI��~��T�$�8K�%�L�Bjz`�~�G��x�#^"D�u�J	wcZ�J�\޵���Aw��M`������vcN���i����5\��
�Ξ@�АX���8���Qʃ�{�C���H�9�H�3 � mٗ'�$g�m�J�k��du����T�pj�N�^����p8�A�5I�9��1�z���j�uf�P�r��FO��M��I��Ud�Y�a�#PQ��%]6������Ei�&������2��}x;(�_���0�6Ǐ$0��1��Y����*��џR�C���
��+�C��`�M	�O���8g��6�ٽ�W���r �8�n�93�}�[t��s����"Y����9)s���|8�F������(����Q��l��@;��".���Ô�����A|Ʌ�Iz� s�^H_Qz�m��K��?l#�WN��?f��u��_�/��nL�́,�cd�D`( �2y��iB���-͂�u/�23ك�y�+$�DR���1�J�d;Zj]u|Wz=�k���@��'����~�����Way�*�g�
\&pt�[k�t�<6��q�*�ςB7~�!虓���'nDzg�v߽{�z�ר��̋*���n[��L}x����l�	���p�	k��OJ5e�t`��p'��AY�/�F�����3l�/��/n�_��g��KY�G��7���º�a�BD�[��Ѷ��sK��Z����/	�z;�XJl�^֫E�-��QlM��6�5=����Sx|m6z�|q��s���8�%��`�K��]s(M]ea�Gr7�^Aڮ��RCdȅ�Iܹ�f�	Uܬ��:�b���J:+wW{���o�t]�ތ ��.�1K�/����C�4��_����x� v0�]�4�Xx�# �Y���ȵu*Y��lu3�Bki��@X�ޘ٧��!.��-�pH�U��.����C���&��7�X���*i����V�qW�#��kH{�j�:L�>���Kp���J2�Dt�`/?v�����6n��I�G��q���"���h��H �xd�����U]���
���"+��죾����01�<c��%�%S�<+s��b)ojR�l.���	��{]��Ε���f|v� ؕ�u�˹�����'2fЏ�[�0����;��(	n)Hp_�7��+�"���O�#h��/S�!�&=(Dtڣ/��K���p��\����7I�lz���L(�wJ�SgW�ns���,���q��
��m����o}�amVW�85.yP�ƴ!�i3�lJ�"�ǩ=r��7���?�.�>�f���3��C8Z��d�w���mC!��B�%���Fj������Y	$�v���(P���Ic���cVoaǰ�����Ĉ��y3PE���AN�5�M���_�2�Z��oЎ�-�;!�����턖��>]C��E ��2H߄#d�T%I����C4 Ѭ�}���cݲM>��WT[��e���o[z�$���@ 0�?�12�PA��$/�*[�%���i�,����Eُ�l�Z�����'�|_A�-���������ښsfxU��寺�ᡸB�x�wޱç
���0L��L�	���c�ws��π�*Khx�Yк����K�l����5��1⍱4�I�H��ˬ`SZ�f]�������'�@�6�����Z���UFJ\t
��Xo��4���쀺�|d�Bه���܆m��PS���%���n��S6#RBO����m���[��o��#/͕Y�J�W�C)����ͬC�q�n�$��4tӀ4�H�P�ZfD����S�������P���H�`����]�<�����M��y^�4v��d@�W= �j\�*CE�F�>����y6R򠆯Th���6���'���q;�Ę`Ae����K�J��J�"'a�{d�M[�HwK�M���X.�U:� ��_��mA6�q����Jr�Qа�!�i�u���k�'�� f�ơ0��Sc�}5���m���A��ƽ�W�7&�h2=����`Y�z:�Ó�ǥ�C�T����^%r��۰"�N?�B����n���8m����Ѓ�]��0���i��
�]�QI]GJB�L��L�>2�To3��'�EŚ"_$!h&��ɹ.��v�0��s��4x�7?�o�Ҍ�y�7��<G�Qyj�P&V �@�
W��� ��4��U��<��Ȱfj�i{)T�g|�,���!��sX��l$���ҵ%���m���	�q-Aա�Y(�E|_��Mp�l9HJ�;�k�z�
�S�k��T�E�P"���3Р��/��)��Sd�B_�l�콷�˺�z�*�7Mn��&Ts�=�����\��>����dE�9�O���j��W�PV3�>�"�>�����pp���hu��+��D���8��qc��_�9���.el�՟2(A�Q�xo��f�Vܦo���U.�Mk��ݻ
�,��#|b���d��J�lS�Ճ�{�R�y	tI5�n��9"�D�tr�\��C7zN�$���� ?����B9�<0oX��h������S'o-��D�9n��v�����/)w�����cR��CH�xc[�dZ�^���;XD����r�֜R�d�CX��e6gs��.���U�IZi�aYF�`��&?��dB�\V�GS�-��q2�x���+��,�1����> �2�BB�8�b�C*"��A���ꥯ�En�V|������L[tO�6Hk�)pT�$������e�b{ �~F����m���''w��q@D�S\����ۜ���zm�����mZ�¯C�ho����_f{�'9�| d���#OR?0�E^���>���:����U����j؇�I�«ɴ*/Mj���ZAP���F�ڠ�k�T?"�zw���G@�����j�̥�������l��}E�R��4��K���\�e�B��9V�p��͡og�We��m��/�b��~=���{_n�n�TI_{���:�}�E�}\+�K?h72L=��Q��D{�g)HS^�0UHO'��Rl�2HgT���R@����@�p��5����4TG�L��#/aN���V���E�bʣ���Gu��Z5NJ��Z9���#3��N5�P݀�ŎK�;ۂ�Y��)��"�_�vu)�E�sgM���jе�?Z`��� O{�������"��k�4"���"R�^f�+X�8��3p��a�\�*� �a��_|�X7x���|޴~[��������r���t�߃
�s�L�|�EgD��r��C<٘��%�XV�[�9<���&���<�,Ķ����+ٯ.�Bxd@�b@��PBV&��S�[�����t�׎�"�i�ܔ߶���>���?�:�V#J��u��ŷ�XVXp"�\۝�961�7�h�����5��e���c2�� ��A����|ʁ���<��԰�e�e��M��l}CoS�9_�tpJ�\�t-�h�! �SKxP\�爀i�a���>�d�ĸ�x^nj�xz�Թ�Xt�49-a\�8R�=�+oZ��D���7�����Jx?��a'�#4��p�ʓ&�>˭ZI\W8�������P��%�>�y�t�,�J���H��K@c:S���E���i�:�V�t}K�Y�R�F`�8Q��EyEp�e�����@nB���y�'�z2f|-7���W�qȗ�sl������Sx��� �{��K&9���"�i���
������@��8�}TueHw\:`f���@{3)�mA8��0{����h��ǘ5#Bo�'�Q�հH�4�s��:�%�5q8MM��L���[�>����U>$����p�n�@�9�L�(5qGa�g^��R��$��8?���4ed,.TZ���"3�s�~c���&�Ȉ��w�x(�6n�ֿ���,�� 2=Xk&}d��Jy��g���[?�2�yc�2�B�,�[���v�,'[RrI|��JP`��)j�	�حQSI�I4�:��C,>�
5� 9��z�}/6��3<z�9�y��1��̑��W3�؏��~�bym3��kh��NvX�&O�V�)�C8�$YG� ��N�-���/�����
b&�޶�64��홌b*�x��4�47V'�
h�q=�z� @����O~g�'G3�`��C��?e]f�~��������}J�Knj�M"��t?:�#�K"5,��:��jV��%�V�^�D����;����bk:�����X���9�*����M�O��@YS�]Q�m���gδ���[�'��[�0˒ģ�����S�<$�]}`�k�xl2�D��)τ)���S���	>��d��D�Iʹ��O7����D7����V[K�]��^��@[�S����I���]kj,۱��&K\`��I������n0s:�s�f��W�P��GO?�%;.�h�m�8˵���5�=;J|:�UT�#�7T��&�VO`��$c�sE��R�)\f��=���ؐ�+���݆v�$SP�#C`�L}�L�'��W�IP������`��˝�_-�`�%~/ �m���©�걀�:ط©�V�G�	9�+ދzF�.���G�,e��*��=˩�݃�׹ݩ�!0P����O�D��C]:�'�y
�fDY���({op������M�F����M����z�[ �M�7_ B�	������¥I�ͧ����ca�	0L�1 /5���2&�z�HtxmW�H�n�z����$��x�j�U��3�Z�#��Y���I���m���8��z� %�Q��yG���ړ�� ����7��´$Tl2"�m2�X߰�p-!�o�*�L7j��������*�c�m/$�{���H���8�hcz�!KAD�20M�>����Kr�����V�s���xD�b�U1J�����HLS�&�W�G�)b�z-+pgn�W�1S�\�bvYm0���NH�x�Df�ݯٹeHH�|�5�S���]�DY&/�L��h�\E���� �Tڦ٭� �c�t��O�0j*v
�>:I��d:��&�EWK;�(OtR�l�Y���C�Pe�i7鰩U�.Ɂ�"����n��-��#����K��?��J	��$S��5��@T3�t��'���>]�������|HyL�i�˭hPX���������Z�ݚq�!`(�-�
 S���=Qkjt1T��{�� u��/�m�F��>�j/�.FF9 [�u�,2�le�ߦ��0EF�N��|> �VnP��3�%�y��A�Ȃ����U�$�-s�lw) /Ӝ�����.�)H�]Ji,D�qڴ�t�C�ϱ&/1B5�b�:j�K�p�@�V��*��|�L��鋆 >�!*�x(��	BA�
y(��	��~l��Z�_�������ip�%J`,�(��:
���ᾓT��S+�io���������)�XEN����� k�;�R���p�^u�S_��f��&D�e��W���o
nX�b�����0��u�Y\^* ���y�Ņ�n��g�$�v%2ԗ�W�>D��@G�>Z�JK��@:6#�%�	�À�B�-%rSF̆��`�0�4l�b�O�����~*@�I�e���[�
^m�;ɑ�^:�'��/�d��Y�*�.��-A��=�}��ԝ7
�g�M6��'�c�$��A�(�h�0}:�	�8!�*�p\y��衉K�D��~"щa�uW�$�����"���*�|:7+��'�����ONa�dT�����9.1`�E�KV�w@ 39�IR	塣0���I
{�����M���N��{V����L�������m�hi��vG���5-�LaK+V(�s�/��)A�_�r_ʡPՏ��YW����bF@����_��3<�L�������Q�.�a����'D=Vh������	
�\�u�,=:W籫O7�
�B�^�^����!�s��6���S�?Ť�WY�,[�qvɕ���zHϣ��i`*[�N��V���K�/�\X�Jj�ɄB��R�j]��4V��`�+��4C�+N!qؤ!�vp�Iy|;�E�H-05v�ܛ���,A�B����[�դ�X���W�ᒏRU}Մ�6l��I#+�x��w-�8�u�3�Yp�����-Z�����Dgb-9���!<0��6{��ȽC��D��lYb3?K��=aZ>�$oש�cl�kn�ĳ���Fuf�=�զj�x��s�`���3�)Ƃ�A�.����4�9+�vw���Q����@�t��)0���Gt���ye�t���D({��P�p� A҈�~m�?[���T�\���vFv�XЍ��K�[��3��{��U���9��;�=ږ�����5=|��5��j�	�z���{|�DtE��H�+��N�S+@��Jf���kѭ�t۩��m��C���U���x�)o�c��1&�Bmv0�sBF�x�N�~E�;��&������6=洚c��,��6bp�����m�}*�ؙcbt�a_�����*����&z���+���@7�L����v�<�c%0�c��x���T� :Wa�;��������|$D6��#����Đ�L���C�����H�P��k���&�����z����گ Z�@t=Jhȝ]bt �跗�a�ń-�w��oK���(�R�_t_�Ա#����w�.O#4���:;񨦫����FrCǳ�h��n7��Ma"����@N�:�p�o<(���n�ƾ��S�tD`	���c�]�F���x�B��v��s)�Aٶ�����;� ���,��	/��jD���4y
ڄj����ڂV���E����o��,[�)��y��a�����j�#�}zD���T�o_�|��b�����|��+CQ%��ӄ�'7�K��sq���N!J4��j=�#�$h�ug�'K�G�Ԛ�g�u��K��(���C����������f��q;�\���ON��C�9F��y�iqј4!�]��\j�tX$�h-D��f�H��"#Y̓5�� ��4�ݘ�h`r�P�M#:�U^G+p��ԷR(^j�A���6�ȄQ�3��m���os����<��b:�?�Φ�Qn~�P�Q�,��ق_(�fF��E�oӒq3j&����R�F0��B�]����M��k݄mGU�>c.X�v�Z-|�%H�ZpY���M$ (W�#%�.g�����B���28/��W��Kj^�%�t��D�gM��JΨLS�����W��Ds&[�d���r��J�4��S��x|ܫ����Tuh�F��m�!n��g�хF���{���{R�@qܡvd�W�ȴ��}h�w�:�^e����?8W%Gi��	{Z�,��8g/,�9�:��;�x���A۬b�$�20���"NLHM�R��:9��̲-��Q��G�	^0kͭo�.v��H�P	dRi1?@�|-G`s��xg^\�t�ukޠ����I�/O/I����v�T���@ey�����N�T9�K��b^MFwy�5��F)^�8�4-j���ft�"�ԞH=��t��8ܕ(<S�~�ґ������5�?um�E��'/��q��Q�����x>iP"����l�i�����;�.9݁�Eu�#\� �H���|�V��R�K-�CU�����j�x8�5��(j�C������r5��,��t	w� ��Z��(<Z�A�;3��y�_��˱��� ��_�G�����\����"Z^�7��L��4ie3 R&�c��N����1�W%��CwQ��4e������cq�"+%�]r��(������4S2V��[;}�m��1A���T���"�!�_0`?Q��Mg�_rW��$�Qw�	��۪�7]Z��b*�-sYI�zi�H�:}�L(B|�V#�t�`����ŁO�P�+6]��LU�4�H����������$E)��5�?�]��r�J|ұJ�
�z����� 2��&R�`>X�Sſ:0��Tr�h�xq:&�A��i��C�B":�~��t��<~�q�Sr+p�.����?���bd�����C�F�O�`oͬL�z��֜����-��b�
Q��f��и"�#�+		Џ��Zu�M�,�硿�,r�1��e����%76C�ѧR��C6���
�����ީ,H�r�u��:{R®�l/��.C]�c�)�]X �?��^d�+x6M�(��#!��l��8Q��7�$,Ʌ������T�����B� L��q���!B{%r]p�,�?������`Q�w���yZ0��9��Jۏr���0�I����ū��� *�A_������! Cl�D�h�V�y���\�j[�'��A^lʦqw�p�s���s���U�F���DM���0�}��d9w'2��e�q�?x).�F���rB��.���Q�ܨ���^�c<=�N�ǻ:ރ�"��p�QQ�����Q8F�@1Jd� �G��#���'�lI���p_ �!�leq��:��o!�nUl��nZ�-�m��̾�
�۞�*7��r��ᓫ���zێ��P%�p�yΘRX@Хֹ�at�h�H45Ԯ�[���@H}!��8~c�.���AG!䔧��֗9rE�&o�f�ˆ>Zj1���^�$F�����8��և4 ����Lf�4^� ㎂��<�xV�Z�8,��#@z:a
Ct
K����]-�I7�:F�Oض�"��_1vA�P�)_��K����q&-L}�,�h4/Z�wڣ^�+#J4]���tX����K��:�/�Ҝf���|�y�L��^/BJQ �߽���O�T���X��[��#����ۇDʴ7ԉOpfkS�c]����[�h�Pp�z���-)�(��m7��&q3�@^�~&��_�g�A�b�\���������`�5 -�K��t毧��|��v��5 "��z�����3��ј�ȿj�>�X�_�b2G��a܆�E�{eU�8��8g+����kY��j"�k�2�����	~f8�Yi�P�X+J��տ:��5eXϞ���h��L�R#9���k�q�h��y?s�٢.t�H,��m��F�Ȣ<�1���F�=��)���ۭ��B�H�m�-�X�,&�K�'���B�d �2�ֿF�Ͱ�{̺]iD�u�ƧZO}�I�����N�ۘ�����Aa)�����P-y	Ř�OB��=�Vo��]a������$���Ֆз�,�3�媎w|o����P��V��%�Oο�6����{iߌ��v��C*{h�A��5j1L@�.�J������ɇ����_����k�'m���`�:$#��%�a��1?A��
^���w�9())��Q$Ȝ���(�@���Q�,�#���H\@e!�pR��[�
���*����t(w���*(�g(HD�G���G��Α�w"�;��Ĵ=oY�����(5n�sx�3( �YE��1~Dȥ\����}�
��"���ʋˊ|�=罘2<�6��	Q�s��#��e�0�k�h�	�"|gv1�p��j�����1����tV�/W!N���SbK����fq�Q�|���Q��I��Ķ��
c𖓀��S����Y�2
��{$K!l����06F>����A�����j���tC@M��� � �M{��J�WwtC�^8�A�&6��O�x'O�T>�lt���r��k� ���:B\�����K�Y����P>1g!`��Bq��\��{�סJ5n9�wR����x�mN�ӘQ��
�B�b����:wZu$����.�#T]H�8��q�HS-�z���d�\ZS�~����J���p�(/4�&�rn��9t�FX��e$~�P��#����쁖�]�N��&&Ep����R-S�ټ\�����[�݇ V�x7�� �G ��6�8�6A�-ī��j��ػ�`h��+"R��CW32�
�fr�o]��5�G֨�y�����VO4�2jf�K[_�#��#�~��D�s��CE�%���"���ջu_e��YC$�nL5x��mh��˚��~ϲC9���^��%ފ�a�4���7zO�Y�ؚ������*p�Т.*G��t��h��e3�'I����5/J�$uz��C۪�~�B�棟���Vr����w�R�֔�s^w��`G��A����`�wwr3?�<���_bY"5���������B�s紗��-+�hʠ,Q��ej3[����j�DL�g�����6	��u�+rO���b�l�F쯅HU����6L�o�a���Rxj��%��0����(w���$��z. e�<���I�>�D�P�_�||�g��Oa��3������p����N�X.*��W[����6�LB�QU�d�6�^/`;�b6�I�����j�)Q�[�Cf Ĺ��ذ�թ�����1�?���>��m!B�ͯ�1O�o�M��a{�;+C96}�;���!���n�x}�Dc:dDwz�)�p�wK��
�i�Hao\��a��pI}>5~�JP�{A����Ȓ
ɱ����mn�PlɁ{*�`5��ِ�{'n�M����g���W;_?S�crЏL���bF�1r�.�/�/m)�U|Rxֽ�KdX{�ř���쒰�n;.f0e�4�5H��V&l�9�r��i�3�ȓ�S�P`v��ڸ^��lE��:��F ��.kZJ��Q~�`� �
��'��ٽa��]��P�^~yѵ$V/T��n�Ё�A��	�~w#|�j_��Rȶ�'�V4��cY/���_G��x�
h��`�dFyp����X��W�&�}l��` u�I@����w�Ŗ����X���-
��AJ�{%e�S��(�Jg^C���$���g�X0��@��g�|8[�r���)w�(ǵP�\!{	kN�D��}�4��]�	�wb �2�X2B��f�O���"@؂5��Z�۩t�.s�xj#�=pD�K�K\�@����F8�#S�?IzT��UmX 篔 �С���S�R�GÞ3��ґ�.�N����{,ǥrޙ6��E�U��GN����	�����/j�*��w�sާ;�"����S�_�o�M̳e&MYn�:s�_Ͻ����8:X���&X,_^*��I��̤	0�Ad)y�}�w R˞��!�_P��K�*�{}�2�;|;�l��>lKm|m��q��(��w?g�'ej��p�'C�sbu����Hc�i����Lť���e&���Y�R=kE��f�k9`s}�����w<�YyG�8��|IG���x5\��&�R^pC{*-�����#Q�J����|�Pκ�zZ����Jdl�=/$�#ɛ�ˤ����ܽ��+D�Ł����E�"(�m�� /��"� �q����?�-�$7�͐���+���U���Z��2D|&:Ph]�-��@Js���*��NJb}�!��	C�<�`�%�����ҩ��׊"��e1���j�AL�l��?�u����o9W�)4��a�
9�T�^5����Fc���f�	Zi�B�7�p�� �:�*�(hֿ��9�x@5�=ͬ��ӎ~PԲ�:�XSK��>W�� 6�׹��_�$���ǁ�V�̋�C��}�C��ؔ��q94����D6�il���Zo'lz�g@��Q �Mh�o��MW4iY7��Q���=!Z=#�V�A���f�#�7��0z�X�C��C/Ⓚ���r�&���.)*�8W�J�,���[	�ς'�������nn�>�S���ќm�g�5c99T�9���CZ$�E�j|���b�jڲkIqRy�
�����ݤ���JN}�"O�'H,�Bz���)T+���dP��ԋ����W�I=<(z/|��@`�s�"�����|��W#f�����uk�A.�������&��zN:�Z>>����=Q�ib�H\{��z���Z�
+xQa��m������z�RSy{-�bB���O�)�P�Jb[]3�)&�l\��١Q���j0?�����P�w$��� z)��/r͌1�-�E��Fc�Z�Q��HQ��J�bM/*�HT�w��V9�G9���5��<����s�`䔀i�`5�8'P��؁��}JZ�%Q��(uTj�@�˱���g`-<��P���� Kϛe�AZI��ɴ�'�ec<��CmE��oK�ߑ�ƌ�"��Z��O����u��?��^(�8�D�_�;qM�\�Vma�n�0nT��L��Lq`�����n�~����Z�D�h����֑KycҞ��䫓S�<��G�8���n��D��_�!��I���,���!'Y���_@kq���t�"܂�jBf��i��|��M�dŒ4=o4Kz((��jJib���Ăd�y�����V,yQ��L��9���˗�X�~�t^��()j�"���\���*j����k�i�P�k%d�Z�uIf8u �? �]�]�s9Ik֔�g �8��1�"L�$i�*Jj����l�P�sⷢ`^+�5B��R���=`4�~*\8-���a6㣲ݞM�eB��*��nFR ^w��l�[L&5�&,�ﱯ����j��jN�iB��}0��E�$HYIi�<�{�	(��hy� hY��>Z�1{U�s$k|5��6Md�s�K|��&���w�&�;�?E�f�(G�"��v�S�,�N]��~����pKJt�sُ�LJ�\�dEE�o��0H�/A�
 �����A9���6�6G�Md	�x�_�t}�.M��
���/��'��F���i#[���,!Ҋ�g:=�0�f�>�̄�7��������1�K�������
�-�6��%�}�0t�Ck�RǕ�(1"��ᯯ9 jE�^Tn��|�z�.S8E��4e0�f�ݽ
��d�X�l��Hb�����m�^��h��z�К`�Pށ��G��TSy�QS�%��{}2�l���-��ϙbN(V� X��*��=9�dO1o����	eQ�gJXe�)P�P��y�5�4C�q�&%C�W��.�I�N���V�
K��FG� ������QH�����#�W�������jP-�dM�y���C�k�S���VGR���������)MJ�Ԓ����2D�8���近���=:7��b�t��P��#��Z�~��b"��g��6�W�r��v�zB~<�_�=����\U,��ҵ�&�[���a~|�ė�:�~��L,� ��l!ڐ�M�&�\��j��E�g4��QHq`P��[	|eЖ�{��XJ�<C����c矲�%e�"��>��Dms�Rl�P�Q�L����Tlѣ>�O(����-8DąB�2��w!����kV��W�����Cb*�i1�(��lG���������0�dXh�]F)#��,e�į��|�<��' ��X,Ho[B������!��eJ;8v�A��LT�\�*Ubs+_��lo��q<�j$@�ةL؁�LX'��_g_u�*�.��SH�Z$L0P�m<B�W�1��T�=��X�'�c���9od�N�B0���g6 x4H3�ߟ�&�W����a������>Co2�乞�c;K�;fs%}%!L�M��Ǜ%���j�#�${����T�$�h�J�I�k<�pE�m^%�G��kHP�s:h	x�`��\����&�;��*��K�`��D�h~���>|�9��\+��X������\�D����%��/��f�ȬNB�m�z\<G�!��mqV�n�B��h��$�Xt��9���?�B�fs'N�!C6�^����*K��N_iS��m��daç|dI��y,�c�b���B5�c}..�:�0�����X�cL�]aL�v+����7w��=�63��X$��K�E�}@�5<�� ����B� #Gt��PO�́��g���<u���߭��}�$���a"�hE%o]�MB��M�3^e�\^��r�s�!���0��u9��y�N�5�����˫��ڮϭO�U?E�V��84׬e�%C��(]%�����r�7�o3�\Az����R۲���j_�.�3A��q�%��⎈�j�ۆ�>�������r�!�IE?s�$lq?�>w�L���Ϟ~��_)60��^���p��.G�c3D��A�v_�>�������W��~�@E������֢rx��b������0�����Ņ�C�+����������Gy��<�J0(7�j�"�.��N(���5dY��}�� tkJN[�������%m^���;���#r�Q��Hx6���ޛg�$toa<<\��bjt0+����&Yik~��KZ��?|���s�"�N%�X� ֣i=-����^��e�͵�3l��d�A�,��\?$�R��I�(Cgݮ+���ѧ�f�=ڴ���5mlRn�Ԭ8?qP�
��,�瑷PU���J���i�D����	ơ��8�\Һ�(?�vH��]c�1�^�^C"[	z��z�k�'����K�c@x��y��(��Q��w2���.X������=�'h�`蹸_�v=P�[cߏy��<���d\�5��4��H -m��kg�\F�}�{��sHg�(�����G�"ǜ�
~5_���JlK��ژM��Ȟ�v��>��?���E>��a������Eu�cؒbZ�``6`����U{��a���4�N��W-�u���zҨʅ� ݞ^��T�]F`�+�W���ʛ�D
�.����]xG�~i�Z>��U���LNZ�>2�D�|S�2�],���qJ	��)���?�✰��7'a1��k������W�8U�Mbн��ju ]�8&�N}P�<I�U��i-�俨�Fz�f�nuH�Z�p;����9�(�Bye�G�F��	��	z�Y��H���t;#����(<��a��^�!D����8] �������hKM
�œ�<r���:�֡�Ɉ��� 6�{�� �a>��_��"��cQ���[����w�S`'2ݎ���Ѭ��4u���;�˨+@o�KF� �R�vC��.�?CeT_+��Y[
�a��H�:���1Fab~�.&��S�&;b�kgq�=�J�Z��i��Pϒ�̉�ͣ�4��`�r�Π>��o��tɜH�1���u��}M�j�ͰH��V.FF@�����9*�ho�Jb����3���\8��S k�I�ah?1����-p"\� �ԴV�XK���E5#w6lH���Ve�۪A���{��j.𫒽�6YX��B�����R�Vp-���"ӳ�,���Ӎ�K�E�^��o�c}���H9q�[(�{g���
�{�J叶��\M�ֺ�x�}��D�?	t=�됔t�K����R�hh )	D3t<��3�0
S�X��ׁ=��d�,�j��+�'�<aP�Ǌ$�ӻ��fCB���$GD�� j���JY_^6��3������m����*ɒ�}*e$��!��
�ze��a�a������^��?\�\��x*���&!��
��(߽�"[�؛�؞��zB���T�k1�M��ʝA�<-�+�����
��ǥ�j���Q#��']����QǧI�bOO�%�Hs�Ǟ:Ka	�����4Y��C�ֶE�j3����:>��߮����1��$�\$/�'��圂�w��*C0�|c���b��0���y�Z�ƭ�/��	QI^���7g��x.�R�U����ŇK�TI>㦐ş�?���m�Y}�P�9ܽ	��t�'����+�\��k:���v�t>����;b? ��T�UؽP�*rU��c{}%�h��O0�U�$��ݶ�t���֚A���ҙ�,Y!�ݷ�GDq}n�����,�C�_�(������9�Hso� E����y�ja�����j*��&s�����C5a�߲7V~zM �|D"�,	�Al�Ę��Y�_>>)�Z�x6�N,N�ɠ�'�*U�M�O]�{soH�$��t~�͛�?���P����P�᰷NG�ef(�b�\8�&���n���'�<���;��}_
�-.��t�*��Hk#V�����
���Q잰��u��i����qd�9����!zmV3���g���~jGa�̋l)몺x� �h���z�DkH�\����`?N�s3�;% 	s6�{�i�C�쓺� �ÖD������/o>�/1� ����Jg}h�lr���&FTvƓ��"2����iw�=��Jl[��"M��/�Ac�H׾j���G�t,Dt{���C�T��H�����	��	Fn�.�z��j�0�7�f�Dn�а:�	�9�y���n����t�(�Q��CD�|�0�oȬ��建���R���W[��T� I�	y�׽�(x���8���<��(,"���W���í���-ofk)�c�!7;�,(^ZJ��4���9)���@�0Tɜڀis��i�ݎ>u��%�7�"�-��"����r^���p�́��s��O��.�d��2RCbn�$<ыi�,�eXOOd�F�V^+�z���͎N5u�����*�|s����᲎��@�0��ƞV�l�0���(`��zl��)S�ՑF,j	���*I 7o��@����p�b�UA��|��a ����6��H�<$
��W[�X�1XB%�I�.�\�x2�a`Z��Uz�f`�:|�r&M�Ú{�UΪ�W�C�A�cCFHӗHVP���3*[s��0�Nd\A�ʹb5����������q ����*W�}��s��A��c7��n��ٹƆ�*.0>Uh��A8+E��:���]Y��#Ś�0a�Ԏ�6�./ym&q$u�2�5��b�QD����	e��;i��g����k$~]U҇	�Zx���,�9v����dW�b�c�.�+Sl�$H�]w�C�X~Yq�	�ъc^����*����C�����
|Ka �5-_�H��:��ZΎf$��CyQ6x(|uo�@ϊG�p�pI)�v�0���1l�[4���(�}�y��!+�CF"0\n�B����M�����S�M�c���d]ʑxuf�k�<�!���K��S`We��:�5
>��Wb���Vr9{F��j(s���S'o��E��	��$�u�����v���/㱿)E��d���iխ#<�6 f�D@�v�y�@�
g9�^(cF
�߂t
�[ל?1��\x�Zy��	��hm�Mbvph-��53f�g�ު��+�
R���n�Нt맇u��O�PcY�+�IZW��Չ���H�0����Z�ޑLT�:h06h٨���o�@�t�[�y±��MR���e��+�~Мo+��Iğ�
K�Qǒ/(��m�Be��(�����8�|�[ʄJԅ2��{<-e�����$��2�S�Ԧ�.�(����1�&��a�U�>�� ��U��h�7�B��E��3�\�0l#��v�U5],Ң'��7�d���4���`��u<��io,X�Ғ[<�Jы��!���~�{�#�	y+�/��rd ��ޘ����ipF��n7HU��r5iĎ���}���*6��z�����8n3+q��j7Ճ�s���vP��GO�Z�|F5��"R�f�vg]YX���3�������
I\ҽ�^�X0C
_[�E��}��[FN����+���--�S�(W�@�4�zU\n�.>k����>[a�|fpGM��|o5���r8�7��Mq-H�S���{�p����.+V��h�Ok�x9N|0���o^x��DQH�D Y�9]5�4���Rx՟O�E�G��HVQ����r��,�f��֛\�o)�\×�1'���y���.��`?߰ѹu���hhK܍cE��C���P��{��%��������L!�[�� M�"
:�BU�\yЏ-Љ&Ȳ������p��Ujq��a��J��
	Lt���M�y�����Z?�o��f���(���|��x߽�J�;mu[�Z��m\��D�&����NN���#^�n��E���6L�����oG7���U���Od����ט�ZA[�xd-��}�G�^	
}ě�.����"8vp>��<g J���(,:EP;�T�8�)W3�a�];��	��ޓKk<�R�=��`�'������)]y��΢?2�x�x��B���c0�jq�6���
{2�A�#�i�s�����`@�Ӂ<n��-�"|!��X+��:t�����	�@��2?ӷj���J����e��5˲��F�po���>�Wc�1G��޲L#&σv�J�?��tia�h�0+��C����W�p���Ȃ��3�P�ae����ӣ��v�H^⭛���kz���d��xA�S��lX�>Ù)�J��x�������nIY��։��Z��ϚY]"��]�.�����_?�Q´��9]����k����]�g!�}�9?� ���j;���1g���Ќ��D�"�nO�71?<fjJ��xr::�y"�2l�V��.Y%�9�ꅼ�˞1٪�v��\|�8��..� ������N��Y�%��,�[�����>�n4���\�	ԿU;,W-�4T;k���/���Yv���SlHe^	�N����ͤ}Ji5Av���#��y���U�&�X�,D�s���;w���'���.�X�����^��(�+����������+�^zN�f�%j����Ϳ�K��u������A' #O��c͌��(�����͠@�lYBX�]�A�<��UR���g37��à�t�e�$Y�������mJ��՛!k��&ߒ_���"t��B
������[\9�����Ǡ��1S��.����K=t�:n$�;�U��1\����;sqw��6y9���-7����lI[����]�m����0x~�G-�����-$�?!I��@�Q�9k�=Xm%.z��٠�έDUMG��ߏ(�7G�9b�vWn
e�r����A�����6%@�n��D���L�|`�>uo�>m	'mQ��P��&s�h�uV����Č�ž���īힷ�3�c�$�5��[M���d�5�.�Kw��V�IՍ,EYy�
��]���ȞsF
{G��s�;x������ۢ�z���'�����^I֡��,OK���ź��FD3d�|��W��i���K��L�I�)�I����pQq�qk0s񖢣9c���zj(C�ACo��>5�W�p׮���t�Z��H�����oo�a�u���W��>hs����)f3���������Y^2�l�K3O�����lOH�7��(N�48�>n��VY��6$����J� �%�������G�}Vx'�Ӗ`#��✨X�_���lN��bC�eI��%/i�*�n���?���E0&��yg����<������;��m���L^�m���?��d��]'	��ǄC-#�r�Sc��0�슬o8�F��d����*��o��D>l6x�&����Ӯ��5~��������EF�9(�!�x4�pc܄�h������X�.J���Ws���q~A�\�(Q��Z�v�ȗ��Op63�,�QM���R���h۰&���nE�H�r܇*AD�6�uf�Fwhʓ�˴��N�ʂ��k.坠�4h�f��~`�e���0Q�����V���qxм+j7nO�M
�vh񶒤����*c9��m�b}�
�⢏���)l���uq����w�XBn�	v٠{���D{�/�+:�ٯ����u�����*�A�����v1�ǫ݀��@e2� ��4` <nξQa�-®c,����x�5+�zWψ ��S� ��v ˚0�%���� �����l>�e3	G0$(&��!J̛Ov�b�
D��#x��Mi��V�2o��^աp���8@'Eu}@2*��K��"\�/3�����=S�������@gN�g�w����z��5ޠ"H|��G�����> �h���3c����Q�q�Ĥ#�ᔞ�q@-��T�o<��ڟу � l�w-g�Wr�aR��F�/�`�[l����O���+ER�N_�:VVL#쏾fJ-����#�M�*�
g޶�x��N:��*v�D�D�'��-��V^/�M�z"�i�b�?�p�Yȃ|����Z�ߪ������� >[ۄХی$|��Q��j�Ah̓��v��e|�2Iy
���#E��k�� ��'n�>/�&�֒�4�a~���3���jq���m�G�'�*�iz٧CW۬����K�O�Ad<&Hq�d���1�^��&�������:�Ǜ�0�η�f��V!�� Y�e�:Z�(`m�^P	-�r��R���W��]�O����5#r�R��Y���Zr����
1��WT��pAf�VU>ѵE=Օɿ�l��T�D7b��=����b�YV��Ɇ��F����Ӎ��9f�A�`����J�� ���r���\���;UQ�_Vkc��юa��"��~�q����m)�y�'[' ɵ�������Y�p���qgjK�c�r�T������0�=w��O�Y�����"���-����C���z,���"5����9�@��FfiNٍ��>���kH>LO[�yLʳ�G����v>�o���q��=�4@��wØ��=
u���zP}Gi��4�گ�ŕ�I�TU���a('�Ԙ�`�L|I�AQ@'�����!7�w���f~4�������%��c��ۙ: )�!y�~B !>�K~UDx��.ȸ��0;ֶ��L|�
��Ԭ�zX;���P<>���@��<���澣� o�K�xW�p/`y!�e:��g��1&� ���\_h�LY&��dq�,��5.��	=�&�hO��Y��ϣqֶ��v�6�0~U��uŞ���Y.�]�9_*	�Y����7�r��A:�5A$J�=hrnZ.��m�� LvUڍr�?���H�L�D�29�Y݈$Ѩt�)�.��5�t�oq����!�X̱��D�Q�4�����"�˗�8�ZSKD�˿��y"8�Qa 0�Y��
�JQI�F޹��k���ߔ?>�\
��_j?C�%BB��a�}���$Q�=MR�u|WeL��[$������D��O8�oB����\B����V�'�ώ�5��aإ'�9�{lb�}� N.1�r��E�'D�H�����j�	� Xp�����	?�����=8�^$�:6@�ĵ@���}��L����U��޻��Z�nb�*��O��
�h��{�r�C�N��9SX�+��Z��2��z�<]�PU v-
4BQ�w£�03����S:��J�hگ �F�\>s\�LC�E�9F&�f�$&X���i�#��.�twv�eYzw�]�M��z�h%�}\��8N0�v���<R����C��h\� ������EL�q'9R�)�!�8��+�s>���t���ԶgNP�=�>��:~Zn8�QV29�&-|��{��+�]�~e��l��S�5;��>@���*"�55ay3�����<�f���'3r��{��Y@�&��l��n$�`~�s�ϗ���B����6�o��׉%��b�u3+�����	q<�H�:��E`�v�1 ����i�ep`M�������T� @pK��t1���L�@<5�46��\*=-_1�����`�~4lI~�Ia��v��G�nhU�� `E����x�&ӱI�@�'��V�h3�$��E���2�a#K#T!^�EXe/&YM�}ij�D�cV�b`��7hί<�x�±��D�2a9��d�̕ح$Y��,�K���L�j|�_��؞-�Bmo��X�㠁i��N8��rf>�?�t��:���J7�ɣ���تB��v6v���$PO�gB�3�{E�qС��ߛar~c�"?�z�֕��Ɖ�K	��b|DK��{���ey@k��p����r
'^�k��K�`+t�bS�5�&S�4`�J6=��e�O��zy������`&[����$H�UZ�A>C2�Y�6�[S�D�2Yf�X����چµ0~d�F�6�N\�KT��GB��!�V��KSb�l����ƿga��զ�&�w�ٝS
f�}�J��Ȧ�܍6��T�-L1VMdA���1�����3�2��2/H���c_k�$��Ia�w���������J��,��qTd>���:��"=m;:�������˴�塴��mO��ȋ:�jF�t�,{���MSH�=�09�cR$��G��D<o�]s�7�y����e#��)X�pˀ���L[���w�O�"���ne����Y�:�K4��Om4�*�"���Ŗ^�������s�;�9�⎡A�҉s��2G}�@��M�O�b��&�����Y�W�E�w�Ex��fw\;���YF3�)�w[&�<�b��&��^zör@�w�RH4�}����=�\9�4ҕEEy軫Xq�L&כ�kʲr�����͢2�kFx��5n�i�4���P��T�5�K�@��#l2�Qߥ���w%b�j=+�	�l��rߊ03J�W��Y��J$��W�5Ԕ�������Dչ_����E�uf� T�m�Y(���o���g�]W�\�g�����]�;p�p��]`e����i��G���p���n�������r?�1/6@��
�L�@��K�� �����x�W=YȎ��4��05�Y�Wb�n�ͅ���b7�7��?Ϛ�.CɉX+�Yx��<:p!�Q�qr	t!6޾�y�Ʉ�eb"�ZU��@3���l��7�c���К�/���ו�o0"?`�W��JcB��
1r :"�Z��`��<���5����~ #Ƨ>���Č$��{ '��S����뾦����ʾ���/¶��Z��̞�U~b�C�gZq\���z�||�$��`�6���S(��u2��sc�n���1�B4����$.��U��)��8�d�߻au�kNo�_�j��Ƣ����4+����r�a�b�CT�(�������kT�>��ר�Ac�߂VkPI�e��!�)7�W�_� 7I����3wxg�׆q�^$O��\�݃�V���D!)k[�� ������I�J`s�Uq�PAM~�,�S��2����%�R���޶a�d��̓��^%ؗ��~�L�l� �ćZ�ا&�����q8'D��\�U��Yp��ʇ�����A�;n�WX�:!`R�5ړd��+-C��1	(̳r�_3�
^�r�F��H�lzp���`"�UJ�F�}{�_�'el������e 0g M/ۮڿ(c�6���
�mE�w|����2��S���V�aE��,�A�SƸ����%���Ϯ6Y0Wd�5MZǊ^���觷�pH��D"�~���|%�4�������mۣ1�PI��_'{��}2
\2�C�u�x$?W�z��U�� �9bjwɬ�����m�NW]�&߲�{G~�`���{�V�$%ft�i����*�W^��	���$�g���|Zw�/w8Þ�޲�S�Ξ qc>n�:.Y�6� )��޷���(Ї�~������'�-��%w�n�%���G"ZQ��X�J'ʉg6 �0n�i���=�"M�%#/��%�hQ��X&CA�6���y�,y��2Bda��e���I��B�ג����ո����;����G�� s&��V��%�e�O=����5��8]��U�SD���E5�a_I�Ί'3�`��"�8��8�U5\H�}�F���P�A��V�bA�8�~��2}��bVC���5I�!Vn�ن�(�grѠ��e�rְ �M��_Zj�`�Ԏ���<UFg�7�V�&���Qg����or0��9z���[w�����0G�#]8�Я��ŧ܂bϜ8��|�͎�UW�R�.�K��� ��]3+=#1ՓD졚�:���$A��秈��8�a
c@|e�մq������M#-V�xSaPߴ\R����( ���i0�ښ4�W������ʲ(Ά))�F�����`	������ࣺK�����'���MI�	��|�ݻe+U��b�Q���qo>51޿ܡ��40�O�>K��k�Vxx̭����|�XN�ܯV�p�� ��ǻ�����T��l�J���)=dܨ�.�8�eD�^��y�D��h������N�N��8tD__�_"jN�Q�SB01����2���t�^�`��BB(��Q-*��T���k^3��8fs�he� �K&����*�98p��@���Hըz[T߄Ư���x��R_B�M�����,�Ӿ`֗*�o�3��(�[�Z�x``@���Qs�Y����UM�KC��P�)������=��In��ڬ9s��c���|�:⠊�[lx�%1b��m~���F)Z*L�ֹ�(+f�
f�a,Y���ڜ�k�ᆡT�Ǔu��%c��T(�J���eO�(� 4ޱ���Շ�DAKn��b֝N���0I�����=K�'>qFu֢G�@-+�F ����H"��\w�s���͵��D2�Z�\�������e_��
�`��3����j�d���?j�;��Q-����ȵl�\j�M�y���_�	s�GA��S7����N$Q���'��)�j��߻��39g"������I���Ƣ=��:�s��A}K~Hu �n��պ��=�K�o|z��=�M��CO��/�C��hȠ}��=ݗ���V /�#ȵ���3�E��ѽқ�T˞�{�����=!A�b��y��=��._�#Z��U��O�s�E�]7s_�ʱ7���N&�Rɬ�s�	�;:c��!pǬQcYB9p�݉.<���������t9��� ��<|VQ?#���	���o,R��5��V���1ʝ��_��E1l�?�q?�)�)|+����~zƉg�JjJ����e�P����<ܴ���&l"�AGܲ�N����biW��+��d4A���Lz-��~y{�&�l�20��H��N"�}�5�s:��*�gن&$=m������w+o:����U�b�ƴ�Npt�Bt������m��V�� [$Ge^��u��(�r����,M�L6�GPn���w�}wE]��}���(��-�?����:I`eq���L��L>)ybtRW�6�SpY��^�/e �S]�hN�Q�^�BlA>1��_uC^���T���%ȁd �"���K�6$ȐO�1.��c,�s�$,b�J�=5\�|�L�`��:��pO2C��i�XV��B��K�d�!W"b���9o���#c໊b����ЏՎ��Zf����m�SO����l0����I:�P ��2��P�bP�������&��N+<t�,����~��U"��]����1>��=Ȍ�yg�l�+�hօdh̲lP�R�J�@��R�Lw9_]��N��,�Ȼ��!��y�O��V�����>��ȉ�_�ċU<��X�kl��|hS�/-��\W�Py�B�F@�;.����X0d���^r?�	RT�'�;+�L� S�����@gC�h��$إ��e��.�
?���9jZ�Kϫ��*�� �.�)Z�����-�4Cс�B���C��A�B�e�_�ƶ�����^E��HF./k0nჍj�:${g���R�[Gw�Λ��C"�n�͡Ҵ$����Q���d6ב������i���.�.�n��Ό��S%?F�XJ�����<�u�X���&�F�ꙕۋKi�Q�nn����]�H�!�ɂ��� +��u�Kޞ��BIa�A���M�v,�Y�Y�;��F�F�sKd��9dZ���Ѻ�`�.�
��S�C���(]�J;��/U�j�BG3P�i,�#x#�jA�uD�d�yK`d�;&K����r�)�z^U��|��ӊ�d�}}��}Y�z�	��Ͳ�s_�j|��e���x��d+�o$᳢������s��V���>*���	3�~w/�R�ߤ`�"�]���\�T�Vwr��o�
 P��M� F��]����'��MA7��*��<J��D�Cuv�wJ�v�!��_�y_��-4g�+Tldt�pewr�z�{�7(�������|F�kQ�e�[8�B_{#����P>��Y>�2ʛR�1��#�Q��ntcy�� 8.�o׉�2����s��Ty˹��Xo��h����8�j��lNV�>�@`����c��ȀB��ok�p��[�v6��r���pH�, ��?۾��߳E��ojأ~)�zKݏ�,���"Gjn\!~f���Y��=xF� ���8�m�JS1 �ĥrL��F����3MNF�#�@�J �yOи�@|
�5A�ZA������;rfeW��p�͐վ]����2m�?K�~7l����D�mL�odY���,�,<Vx E�5w~����+�\W��DT��ĺ�թ�7�#kT��r�<��(hI�E�L�e�l2�JvGg�@Gn� �GȠ
��h|o�[U���js!Nh��Y���5-k".���P�q$ϟ���G�&m��u_����_�V�|��W8���N(F�!��jo\�J�m��fk�Fk+#�1���,�cK����n���F�ɰ1)��I�;X��Tè"��X���T'�(q���i,JK���o�y>��J�~�3� &�ƕJƂ�uZ� D��q��9	0tKPҸs���v�2����3�-���b���#)Ri�����?�2]+�����M�U�*���s��{^RRL���W~��k<j�wB@=Z;�F��+|�So#�\ޓN�����5K�5I�G*��u�xV����)��h�Ibs	��1(v�\s�'�KÃ^q��jcήzT�#2��?��\3(?�^��C3��P���C#�é⧁��ȻK�P
�N�ԩ![��*}��-����:��;jb��M���f�?��Ԟ�&aYzY���/IY����Ӄ�"G�o�4�tr��Qz���+��׳��E��Ə����Xۮ�^;�|�\t�g��I�8��%7)*wi�qQ�*��|�`|#����yJ r-%�z��ߴ��G@�׏�S���
~V�(��r����&�I��I�RܵQre�G��u���~��݉���y�z^��v),�:�yR�o����x" .z��2ؘ�?3�h�Ύ�u�!>йQB�Gf.?kA�%�c�̦�.9D�����!-�u�S�!ꔖ����x�+"�!ӈN��ݡ�]5KY�?=\Q�����w��Z̺�Tj��8��� CB��)�q� ./l \���;_��(r$�݄�My�f?I���4�cE�k`���� ��'I�&.����*�X/���"Z�e����G��{Wu���z�h(9�s:�x�p7*��%�j\nV<y�ɑ��S�n�|�f�5�u��'��Ҙ�[�F���1-0F�����`�E=FY�H9��o�O��٧��Bލ�� ����L���5+�����$��K�%?y�����c ���ףYk2�P�;�3�H���'�谤�t�<�@/g1�4���*�0�&�}&^; ep���菨�>t�)���%E�YKQS��%��S�F/9b�V[B~�2_<m[��4�f��pu�TӾa�V��<���B~�\�<j;�6q��Q�S�h�RaW�����;n�Wѓt��i�\�K�w��s7���֚����|\x��QP��.1�D�=w*���:^y�(�+1
���.�} 		�[���oq��r[���;�8���E�k��ѽ�ᓓ��nIF���I)�`]�|��_����z�zs�C/�"�$�<�~*G���i�1f�,���%�<HU9�/I�`u�r�r;����?��Y^�G�rS��-�����ƭt�ЂC�Xf>W_��o�أ�f�?�)���ا�k�߳��Ƽ�:!c.z*�ܗ�N�X���ե�9Ў'� 颻��K���0M�z�(�Ƙo�sT�����Ƞ�������Qt4���Oƴz�$�[�CnU6k��{��RRv5g��ĖC��<W��3ڛ����?;��!�s���`��+η
G,�����ח.��*�����(~��v�<�n9����ʜ`J�EX3�e����kr�J�\RүkHI��S��w��A��׋5��qk��0^�������aMrU�+(*/笽�ژ�j�� ���/���*�0b)[�]��E�E8]�������zJU���n����A�=>���HT�L;y�6���j�y�z\�ᘿi�9h�B�ҿ����j����K����8I\��nI��"?��&��^��֑
-T���u��ZР��=�bI�����T�����E�:��k�������� ��;(�N5�v�i��4����ɿ ��3o��)�ԗ��Yz�ugN��%{X��H�F����;���bi�	5
VZ��v��yj�;S�._������$��'�S����m4�p�F£ �����ڸ-�LE9�dc�qOi���ҾTlAn��6d�y_��l×�����f}�QB�S�O�?�s�E�K��
]�c=���&c���2��|�q��������
�3����J ��ʝ��D��K�����g���>UC֊��{-�[���biz�h��p:���Ax��t�D�<[�*U���Z���ʒ���J��3��i�3Uy˿�q�;������8O��Uh�wM���9l���w܊���xB���Mi�Vd��ӖA��~�)��	_�
$=J���v����i��΋`�%Î13~N�p�\��)��i�
�3��6]�IK_\���8���؍�Xb����u0C	}?k��67��i�tf���6��|�w��*��CgT#KM@	��נ`;�ܾw�{�^�l����8b���*�H)i���e��˝�:s����UX��:�O��d��d�A��t)ȋ�����%L�fl�&����V�}�
2���18c�*N�Oqwd��Z�������f2�e��^&+Q&��d_N�h��#��nx(�Я�����K�����x�qP`�`��?��H��z.�R�hF����A<�L����)�ӫ������{\k�����{�3&�·���DKiH����yȯ,󓲉;����Λ�n�`k��̭=�Ҝ�wձ�66N��٠��6�$��nle���K�X��2����� ��),A�'2�X���7KHI�eD���2��s#ӑM�jQӜĹ�*#�N�q��Q���[}� ��\^.q���MH�;m͘���Z���
��ª��剒�;9�� �t���R&NSF����&�A��,OQ�U2� ��s�CR4�h�:M��k>þ��g=��4�9�Y7	����l�Ϊ�h��`ϯ�(j�O�,�m�2��J��s�o�]\k�xZ�N�6D:ѧI*���bZ�U��mU�`�#���7�<���]�-d�Ճ!p�^���E�)Ixx^-���90i�ۆ�W��}X;��ژo�����0#�}�7~�������1��؉�cC IT�!ZŅ�%�"í�)�r���L��%U"ˏ��bɡ�i�ط,T�5w����� ��5c�	����Qth-�&��Ꮊ@�a5�#96�R�>��&2Vw�2�Lё~ԫ�C{���/��]�� ��wU
�H\rչ|L�R/��K� J��]��.����DR���T�Ծe~'V�&�[ɧD���#�ǡ�<��i����z]3��>I�m�aX����L�#��z�rW+1]���1�U�kS�bp��9�T�2�q�#�]5"41]�w��\��ɣ7��N���T
6O�A!SY�]�%��]�̖^y�
�8�r��1�1�Kj�){jVi���3u(n4�mU��r��;0vE��s7�?Q�H��i�z�E��/p&V��0�k��p��`i�&�K2܍M�E!p�x��k����2l��Z�*�B2�K�2���a7��ŸN�\WE3*$)��߁uw�e7���k���g��:�|<Ճ��K� -Tc  ���E��qo�R�g�@$q
X�~87^`��+�n"�\�,ˍm��t�0*�eW���Б��Gk���iTx�N(���z*
�=LSDCĖ��A�(���ҏ}��C �"K�5��J�n�̞1�^���[�δ!��b�L��аnLl�=!;G)�gv�s�ґK������ߞ?C7����X�1�1-��7%1�}	�����g�v3uY&��0뗂۶�S��j'�@	5fg�t�*����T�>��?5�]���!���b�K���Y���Z2}�T/՝	�O�_��E)1F_Bu��q�� 5�\�B�L�f�n�O0��5�
�D`[�T��#v��OS���E( �GȾ���O!4LF�г��=Hk�Fg��������ҷ1���[v�O}<�V�� 9牁������a��.a4���Ԫ�M	}zT���a;�QZ���'���Ժx�>R�܀�A�B\�Yʝ"nB����AW�u��)��7��tv�ON�1���`\���}pcPF�R}N'0e�N�����¥\R"�����po��.�<�����
)��?��SYN�1=� ���Ws����q�5���߷�R�P�[�w�A�s{0��
��q�m����k�2{��sB�{�l��Zp���k	�1�9H�R���<W��mC�������jo�?��n$�p���z
�
�B�C���P'��i�b�a�3��Ѓ�S�י�fB^g�f�n�g��r��� �
T��[������T�:���5T建)@��$�ˊ�=��()}i\�<���x�ٽ��5�Z�>S@;�2��*xJ�!;1�6|������`Q�t��$�)a���=�]�v^�CQ��4{�	`��s�m?=�s~�Pl�1��� =/�*��y5���4RG�A����&a�����a2�;��|���J���s�=��e�-"X�s�_r�h��9��F89����ө�w�es��%�����CK��(�E�!S�2	�2)��?�!�*e�W�X4_�t�ԓ=w����M ��7����c:Ʉ��L �^���燯��!�5fu&�x�)�CES���f,0�Y�g����G4�� L�H�&�X��ȸ �*�0�k�3�����9>���C���ֳΌlz,*w�T����^�d�c�s��يv���_���M�_���=�F`��̓��"n}͕������b˽DR}��=�����$`���x�5�3�tX���Я�Rq{!x��`���A��;�K��������q�������J��0uw�h-�����%��!�Mzŋ}!r�|��rh]�A�yK�E^�ҦE�Ζ[��C3��҉�7'�e�-�"����_,���9�ܨ��Ɣ���gP�-.NKΩ�m�'�no˷)O���X{�r�|(���į.+=Cs��KBe�K8���HB�QH>��		�a���8S�'�"sF���}N.�-OgOi��H��%���XD��Ph���5�| I#�����ٲ@]8�4���)�[�V?W,�v'M���R���;�⮰k�Q��F-�j)�>��������z/Ho�f�5�;�GRA����p	�<�˪�m��pC����6�����m���5�������c�1���]���ѭ)�~����^�'�/ZSh����𦦒d�`����ge΄���е0�b�*�IE�6,P�.��$�ʴ����l�i������d��D̵%�N�#�!�W<����!�q�gh3� �Dy�'ڪ��ӏ��@έ-L���>�P��������!K
�c����ޙ4���H�e߾�5�Ξ��X�Ϟ��ko��ޘ|���#ub�>�9�����Z��x%~;��F:i���x!M�Qf�o�ő�+�H��X��	�7����o��Ɫ���`�*2Q��t5����ӪH�D��r�>����v�
oR�a��J$�^���Z&;�,⨭k�8|?4YtO�bq^��)�W�䪷�@��IRt��~����\��L�%�0��@f�<4!D}��0�࠮jhB1�8�;�=���o"��c����s����K�}�$�����dU�B����ü�-�헲��?_��ԓ���Ǵ  Mx�4ݔ�c����$�]
F^T��e�֯To����l:��ϲa�A5�x�ȅU�����ac@���X��j3K*��Ͻ��4\�դ�
�" �B�)��ڱ�?o}���5ϑT՗'��>i���JK�ސ�Z�%ir��*��w���������>UH�k�i����U��bP�������V3fȍ�L'2�19���`^!S���%��}2F�̐i�o�5�0rε�k�P����ECH�����|�1�nl��ig4�G�N��o-�޷�!����\�ɄxY�ĵZ`�!@mUX��6�7}�r�)`�ɸ�2���,�!D��v�ǥ�,�Q�$��2SŪ��NoP�������'�5ַ��1˂y��n�@W{ry�%Ϫ�rh�0z�����6z��r�1��g�1h����j���]�Vzf_O��~˜��|�S�x5ڢ
��}[m'�JE+�����
�mF^׫���@�y�)t0�ŏ>Z�X�����I`�>}�gR���������$�6\^�LgjZ�S�o��ł ��C��Ι��P�����vK�5l>����%�i+����������˔\{^c�����ҕG��g�����n$���N��XޙDCХ����S�:d#K��w�f,0cM�ʳ҈w�-)���9��P3��7Un�aj喡ɨ	J�)�5Z�c��\�������i������N�C�>�b}G?Yy����CzLo�$_��|{�h4�N/�S��N,q�\��׍P��/%/��^F�[/�[�	���᭘Y'����Qq�]���Z���>
���e��Wb�G��4Ģ�nMc7Ώ��_���k`��a�`#u�z��3uL������^�o��w\�_J�g����B��!��׽"o�a*����q���b $oҤ��2*�P !.cp��	~��t�T�
�ݹ��6�5J
����]�j]Ygʥ���\�/�N-��qrTd`48����F�%5O$�_ҥ*��57�����i���¯ ^#��>	.Xl�[�׳�((�%g���ꪛ_2w;-��L���t�:Aiț�B�%�
�g5K$��q�ն��=.l	�$uw�����ң%���ȃ�Qu�B���7B���L����d��Ⱦ��V�RwDDü��)�'z���	q�mK*H��$C
ĩaR�yK%@�`U�FYeW���d��JM�2S6<�d	�T�|�=c �$�̎$������Hdk���?P8q��E^l���'�n�ۡ�m�qfm?�W���s�Vq���D!x{�i^�wb�.��(T��<X݇��a��1lLM����L�!�(���lt0��U����ȩ����c �����덩
йi�vvR߭Y�o���N�k�������?VE������Ϩ�}�uiq�߰x +i�Xd�?v�Ry�N��7�Rit���J�ռ��x�-'8��i����|��G>XZ�=Q/}����t�1|�2��=oO���q$��B]��v5���G�*"��N'��7Θ���ȩl3/;.�B��oۥ� K�OIK��,�m�d���/�޴��;��3M�f��F�	�!<�I�6r��_�pB�.�U���'�%)tR74*G�4`��!9Pi¿�6_X&˫a�s�ܟ��N�x�ie_��ߕ�S�p8��Zޥ�O B�s��c6X5�z�����:q�����ȌV���������Ht=�u���N�Ť!���sXב��L���Ia��XKQ�Өn�̗�{\þT����4�o,,3"�H����EL����"= 9�.��T� ��̯�����W��À�iW��]ɫ|���2��N�4�0�h������f��n0pj?W.�'N���a$�
��#��1�1�ٛ�<�4�!![`��R�Mz�,Ɂ�Sl���3QL=���\dg%�/$P>���K��W�'�x�V�QD�g���A�!Q��	H	ѬE%��\`g:ཁk�6�RK���V:e{?�6d@R��S+xx0��܍��7/��!jtC�<E�t�K�*�l@�R2� 
��_�����dy����>)XI�C*U,8��v� ��[�+�������'<ht����c��P;}�Y㫠��I6&�#�D��X��,���|���$�$��s�G��-w�ȁ�<�_��IM�� �*g-{�C�)�ҍ}����\t\(?��Jl�K)��Hʸ�Myq�Ls�}0���)��p{�q����8�:ڠ��g Wb��F+���xE���/N�]����F#��nk�Uѿ��� l������ 	�f��ZZ禤���o��S�O=eC-ư�^xBQ��,�?�s}��U<[�m�]X7p	����m���Zg3�io��T�^T>�}�서�o���=߁ڲDx�٠��i����[�UQ�G�_����B�J�Qw��y�[�Ʒ8Q���C��������y��	ŧ�I�zՂ/��̮�Q�V��*���z�fM�#��'�)��F�8�����9m�l��i���j�3�3��)x�����c~�2Y�<5`ԩ����}=O�$��'F;V�!�	����Q�TvLQ
���?O�*���!ˀ�}��"��!D�G���2ia���胃�'t:�������71Λ6k:���X/� *��� �Ǒ\j�K���`W��Y������Şo�땛	H,xH���.�9���_?t��a���:�U����w��z ��,�3p`���4[g%t��Ĩ���Q/m��w*8�4��k�n���:Z��v��$h�zs8��n��>�������ԫ94^!��kh����L&�1�x9�ϤJ	��&=�o����ȲS��Hz���S�C�K�2K8~�2�@�t�~�/bSx�K�������WAA')����b��è�<�2�OZH֗Ù����|B+`��b��ޛT�$'EfG�6��{���7M��e�l\�����z�`,m��ie�\�-�և�D&F^t���y{�Q"�gYEM�e�c{ɬ�}v��[�B$P�y~j���� ���ZS�A�ƀ�b���>(���i�}1�P��|�ѧ!��4�� &KU������E֙>�u[a70��W6���Ү�C�����O���4����*O�'����C�hh�����[?� �za��d�"5�g���Gq��J�Sq�	KZo�D!��d���5O�)#� �X��'�y�x\hގ%?9���Is�L��{}wN�3�i�R�1�i�*�j7.n-v���V��K��Y�4N�eڢ2�A -@�d.܉Q����� E�5���!�� AR�<�\�ƲQ��>3*zk�^�UcI�9�#��Ǵݯj�� ��;��u4.N���, 349 ����e�����X���k�����j�6�x��K�ˢW��y�A�D��5�8��0��s(x�&u�t����l�[>�m>�;��GYx��2��Ey�^��"�y�����+�;�t!�;�=:��[��fW��T<��& ��2�-����X���w����9e��܂9���q�pX��h���I��x�J��g�Ϙ��7��v��zvZ.�[%�+����]���}�	�!n���aT�YM��3���K�s7%7x�UI�k�]a������+�������*IYN��|H7�<��'p����[3�='r���MJ��5忟*���<�S�gRR5�e�f�$(��m�
���zK'��`q2������ʆc�Za�!��͠M#��ԸP�{,j�J���TG-�̣�@	gcU=�Q��� ��0P.��|� ��u$S#Y�:ľfL�>�ˈHFI$\��*��.���N��k��N�x﫾����w���MR���Fo�`�%��Eo%OoKf�o�΃�<y暱�-��v��Ғ>�hi(�V2�b��[i�sPZ݀���*�Yg􄲗f[�<њ!%�׾�H��|��!�%�V�>�Sĳ�ZJ^����}��s|2��B��~��T����ͳ�L�+�n0��J��@�eHW�ṱ�]�&lAq��^/Z!i���,�Fon9a�X}�_L�>螩ld��p�M�#�?�9�@��2��R���r���v0]Ueŧ c��K��
6ʅQ����}ُF��͘�q��3��7�T@��b���㵖�d���"6!q*}��v)���Jedœ����66u��6s݉��5�A����˩�(~�Gl��_�`%�IÆ�/���ǠhWb��k{�G*Y<�T���>u�0�T����;ʇ�!n-Q�ux<3yY�[��!�t�Z��A�8k�����1�u�YG�����W�'"�t�m�]C�+�N� c���rt�=�����;�"����^�uCJ��Ʈ��~�]|�٨1Dдt� �q��[L�����Q|?��~��3�������J֊N���N׳=���!o�ѡ,�#��?���&�%�+}����ycpK���_l��,������̀����6��h�ȉ���b�h��"By����X��0Z4iT{��N��Fl�!hC���m��,��7�!O� Җ��ι&�Ҁ�"?N~5J�	=�N��(sc�Kf���l����2 ��9w\�O����D�8}�>��LS�fU�%9L�?��]礽�p`�!$Y�r&�*��w+�C�M�����{[niL�pb�xc�P�ɜ��B9�{����N�j���꙳L@�pDma��	D}X2����G���=;��*�6�6���fP��I�L����SA�}�8���81�'TRY�{�0�W
z
��h��j��N� H���$�bF7����gp�$Xh��j<b݄ӵl��^1�gcz�?;�9��ef'�����@��ͼ��S;�C�ߋV���z�T��X���.d�P���q�ɹ�sQ�+���-���7�oj�5%�?#7ݷm��Y@QK��Yb���ޠ|x�dܕ�[��8��lރ��t^� C<��Y��=��#����t������e!|��BdX�53-��I�m2[�e���F��tAxc�Ji�yu���	����.�r�uG{X�q��mo�x{O����+B��9�lzF�ZR$�#¦���+������I\��4���-����^��]��x�o���/ =Vu5�5��R������;k�T�;��ʽ�M.�ӟL#%�?A"�p��˲L֨��}p�3���w6�b���̷R�Ǜx_!Y�H�H�3t���8�O'�O��Z�`��R+�!��j�T8,{F�pD��Lx�ϩ�n�Vm����ꉧ=����õ)���oP��0ݤ�c�א��)W�D�c�6�������鼡�����v���f�w�23�yL� ,v�,CN0�\T4�zJ�#�]�!�O��4���E�O�"+a�h��`&��!�;��<�ޣJue8��a���b�_�y�I�tO���\�qǦ�N��sA�h,�,�U��7B}�NI��@О���%� S�HcT���D!&y/��:���j��-�9?ݮH�z0�|%}�D���	B�O3��sC1�z��:��C��Ư�߂擇D��� ll�\�M`E�o��X�@ݺ���%@��saK!��ꎱP��.K����`����;�^0�$)"����7�h�(`��Z�Ŧ�j�G�/-E_�5!$��W%�:!O�`ƍ�p���6�ԁ��U:�	CI�P���\O_�6h�� ~��g_�z;ʧ���!�!�Σu#�u���1b,8i�	��R0�M@Hε���D͎4�4G��E'c>����˻W3^�\�8Y�LM���}��ː�!�I�F���i���DK�"i�����V�^ |����֣4�C�c�*��n/&8_�&~�~n f�~����n����S�]kѲl�sw�Ȯ�Wv�I�ӑ�W��]u�������jn�7��D���#8��x���7 �%�Z�B{�2����S������G(Ӯ ����O�g�<��T�9TP>b� j���/�������Θ$V�j��b���@�"C�z$����!��]�<>��&�H�����V�r>$W!�TXi�K��R�	<��d�C_�M|����X�u�q���&"���%Ɣ.�nK*�00�T"���ѧ6s�yf�TV/̫� \�D�U���`3��`�'�	C��:��%Y=�<�������F�f�d��tk�fK��h���c���:��
˦��oV]�1z+�tP�'�N*�2_�g����#���x �TBe�B�U��h��5�����Xa8vq}^Oqx�S�Z�/�R�[�g8��G~A��P ѕ�@m�J��X��	�៧g���Q�(j���LT��B��5`z(B0�2��6J�����<]kF��ߡ�{�+gp��S��<��ͦ�D}`�e��K(�a������Z��&���t�������f{V��A;��N�ہB�Ù�fU9�+@���w�Ns���B��S��_r����� �n
����[�SoE~��Ȥ���9�J'�>6k�l�Di����{���h3�S�$�r����J�[̴)IX7���q�� �.�?p>p�D"����}��0���*�6
6t����a�>fPw�n�WAd�$�"ac9������kh�S��e�����V��\�T���p# yRF&�	�w3�d�#�L4�����	K�2[���T�#M4<��e���<��n����) 4O+�/Ǚ��9�������aqU����?��'�Q,:<�A�3�,�,h��
�s�t-�t�N�q>��Ys�z��'H.�*[R���Q"��lbPڂ��
'<�`1�*T}�Y&���P��kvA?
h$��-���,�\�r�y���O���D|`�4���� ���M�җ��0=8'�6���U��\�(k�dz�vn��c�	3�1�WAS���q����'��	�r���juO'@l
�QP[����=[�8U @�� �SV�����>�5����������G��-�R�չ��6�B�k�W���m[E��\T�����~V�&?l�G��43l.-�G[;$6,���k�Fggq�x��U[XNY����	?s���ժ��P���N1�z��!�Gi���BH&q|�p���]�gg��qǢ��m#sB�Q¿[_��<�^ҝ��kkh�N��_����X����_kj�Y�/ML��$`@@$\��Ϩ��W���@K�<�Yێڙ#0U��{�6����:"�H���3��Ѥ<߂��:5�3�4�b��� ��oʻ8g%9�?vQz��>㧎�*�����A�]��t9�t��P�YS>��rnq�l�(�2�lX���po:sk�Ɏ���~�xC
����9q�U�a[B" q>�����H`�2}�~�qo�]#�rp��g�Ja��թ���X$��C��s*�B{�?ܛ �2Ǎa�l����r�3���Ё78G,y�ȭ��pY�j�7�U�(p��
BTìy�G|j�ܔ�T�Ȯ1׌c��˘&e#�����lG�%�0B�L+�`���Fi?OAW�K����-_�]���l��6-�N�m��g@�VQ�\�_��S�kYEOE�5=e���:C\��b�4F�:�M�A$t���-��)�Q�;�#sP7<L>�Q��8
�GL8�yt*P��z�G��h�����}"wu7��ָ[uY���UW:j�6�,��`�e,��:oP���1�	���]�5��"J�;��Y%����B�Ǟ���+y����e�P@JȻ�~�1���oK�����c��ݷ'zN7���P|��~�h�4��.���F�1�;��0ֳ������v^�q���Oē±��`��B��󺖵Ƀ��z*pp`�
���)�ʅx�~�E�ܯ@��(����Ca��
�e}�p^���=y���Rʒ�f�v�h�Ki?�G�$������
���i���=�j��{��g*��ΘC��^{��F�z@(Vh��{������Ek˯@���H��g:��_����$�-W�-4	К��F��6?�!:�WSZWNe��7_v���P�C��~vbb&Wb=��8�I������5CT~���/v�׆p~��M��\�3b�����3�gX��8)v�+��y�%���pX@	�#Kh����	�o�N�N��`_
Q�� �I~� �Q��Q*��g1�?�����T��r�s�uMAn�Ư-�����Ɇ�X�e����s�yGP�:�R2�KS�'@��sߴ�/���vȣ�� h�,�n�h�p{���GoU���*�#��7S"w�����F+RY�D@��7FW -� �Q�	��їo�ꥆ��c�G�k�v1�`J�a���1�+�-�MCܼ������׈M�����T��l�r׌�$�A��l0P��a�/|��h^��Ҝ7��;���oZd�'5������b^_���snb}b�{ޓ`,UǼo�
^J�-��c�CY��hZ2V����K���l�����Y8��}=�pƿ �ΐ�%(�L�lx�~�'�}oiz;��T}�M��W����SZ�Ņ���)G�H�٫:^��7�p�h������5?�xzI-�H�c���=�d;¦�I�&4i
e�]rhjvOo)%��3ő����0=iCC�[4O*:�����]�CGo�2A�Mv���l�fo}|Qʌ�R�ԃ�����Vt�����Ɗ�6Ncl���n"q!�8���Hi��f�p�mIØ����s�������5'���e;L�c=���d2!9R��|�^�$7��?$rGWN����b'��K�����r)��� ���Od�B�G���-���h����J5<�+k�����t��U���\���!�	
�-P���tt�伓ʝ:F�g�,d��*�I�WstG'��v1Úb\RSR;��/6O�7;��腡[/o%Z��0q�
A�*�U��.'Sf�5����7MG
�y�G�*��h6w
��GQ�+��)&��:�57:O���u7k��䧆*�~��	�g�Ǟ�fy`��'�`D�w��Ow����=� H&�>!��9�.�@�g��|��jz�L��W��R��i/�����cf>#�z�L}��T�j���.R/������	ӿ�6'�DK�N�=lvv���I�7�I��L��#�N�y0�V�0Y$RAL���+z�ߜ��vsp#v�f{�ek�.�!��r�w*�߮�a��y�e1@��1����XU/^<VNN��S)B��tvY~���#� ��pˣ�`48�����ş������va��4iZ�Sw�"b�2�6�]�� ��n�4,�&���c>�=գ��T������jt(r����,�QMl�配mݣ����[���[FH��-G.�ѩ�a�I��RqTrr�i��[��f\��a�`8<�~nn'�3�����9�)9}����r�K;�s�<KH��=�o��$_<0�8�0�4����'�2�-��{x�~Du&�uA�t��4Җٞe(��I��i΀
'�&RDZM	��S�{o15zD�zY�p��`�L�>��TP�3g���{�07k�=M!C��y<�$�O��� ���`sfJC�
R��+Ρ�S�gQHv��lC���Bhm�O-Ġ���U|s��8V�EĪI By�yy��9��wѦ��7�35�ۼ�(�zs�֐gu/+�E�cI^�|<n��ͮ��~�ŭ+*�	e�Z֎�*/7S�s:�#�,�VaF�B+J��Iba��[p��j�o_�S�ۚ(��G��N��\/�d�E7T�S�y��L�vf�3\+���ē�s_���4JCb��b��A���N�.o����DK��QViS�-X%�qz"a������,�4��_&q#l��}',�&P+�Y l�3����J�q�.�E� �@g�y&�1��uv� ���K���![�n�~���t0��?�o|�A��V3R�N6��`�+�u�綔��B��V����]-6��:���a�
MVU0�wV9��mֽT�����Q!�u�4�P�@�	)ʛ\ՠ��:��_ԨC�hxa��Mv��C}\��)�J��a���m�J|S��0o��(F�9)����lP��V�;?��.6���z-�������@\�� m�ܞ��v*��uD	
�Aio�o���(���g�3�_�"��_�xL�ag�H>r��`�$� �����l�Ӄh)��������>���6��3��Z���l�Z�"���C-ye��2��CH�5I��w�<������O��MA�|��-פ�km|�tM���*�R�_ʭ�xN��J�$�F�N��m�;Ti[^�E��d��ٷ0�t������\�o�����oگF��vK���1s꾴�Г��HA�����rv�.�WH�4�p"����P�:k*�V^�N/������dy��q�;=}�Ҽ햂�s֪����_����j��Ux�%�(�F��|���]���In5��*d��иF�򙯩��_"-ժ�s=O ��bK�F^�f4�����Růs���R���k�fa>��a
�V�F-�B2�fn�*҅�B
Ԛ.��%R�]�5�
��T:��@��)����Xmo��{Nj\��S������7��oꩦd���GW��f��Ek�x_nW5y�=^-x�_ML:B���٥�M�o>�����U����f^#Dʋe��e����.u�bH�M��
��H���'��V���ʧ��'����Wc���B}���C�Oj�]�O���	�-H�?��k�l�0�[�m��UM�_G@�~��Y���)�S�ۇ��ƚDڄ�ڠ!W �%�ƗRbxDv��޳��o� ��~����.�"��}�)�{RS����0��a<-��c%П��0c|L��%�9�RI��Y���pS�~';�����8�5f	�A1�*Y��1���E���ŧL�_[l�!��d[�@5� �����=^�q�p�����du���������(�H��J[�Z�o�K�F�ז(8Z��!h��1wt�Ϳ�HF��)Z�M�T��-^�K���Q��(����!㶊��k����7q(m~�R���~�L�!K���};���9���<A�'U�V�Q�>r�-�9"4H����n�v�FsU�ʳ&F\��45���&(�'�b~�D�s�9K��	�#~N���Q��8W������|D�G���My����9V`H �*O�۷Rc��R;(�M�@� -��7O9/�uL�KvQ�@��d����pWn~g}U���,�Q�>�'�I������Q֋r�4�%��NuT��͙Mǆ��������~1���b��]Ȏ�J҃d��w:yx: !�ġju�`��k�B����Q����
�ԿIB���3/ �]�k_%�������G�vtB i���4��k��+�3����]�z"�UO�`�6���d�$c�Z�v�d��jޔe�n#���m���h�H�>
"H��+��Ͼ�_M�� +�f�Ƈ���Q���R�@v�O�fu����~��I��7L�J�g
����X_ޑI3~��`R��C��e�UׯvYS>������Z�4�Y���σ)�����č&?�0i�`��>�-͜A~�=~tT��$xҳ&^����ҽ�k�� ��e%m����h��9�0��5��C��3'}��B
A���h��C������7�:Wz�#;�B� B��}2爣9>�I�~JUC4�Zp��7 �c��G�A���Rs�;�\��R��e&��2 �z[:�"��(1`� V�)�n	=U��I��ې���\Y`���ɜ(��P�h�y�dB�c�?�<"΅� O&3������Ս�l&���I2���lojhV�>A�\�N7�?���H�>�̇��\��D�.���3P�E܃��$S
mdgLJ�3������m� �J˖�6��Ѳ�\i���9�27�I�1�
륦�X�m��U�P�a#�0`�e��(l��Eh���Z%��.c
��:�}}���ض�T���ѮU��~,�e�ڃ"�j�O,!T���㿟_e?>��fiZ���a���oK�2�뗕>�	K����(�M���&og� �+��at�5%�9�����D��M�3+(�U����X��P�I۩`%[�cŦ)��t��/|����}�] �W��I�pMj9L�5���u�Ũ���uF;uZG���ҵ�B4ف{�L\���Qk��ѵ �����
��!�{EX�
Y�qјO!�ȁ��y4(?M�K��W^Ҿ�[c����V�ȼN1��Ѐ��f���������N��G%��
6�I`�"���(�"�(���|�I���dϔ����6�@��;�7+�a�A���K��� ��^�
W���J���0�)�C���N�RG�xcs��"D������ܶ�n)���4WJ"�VgZè{t�g���<_У�D-�q��ka\hV����|k�$7�Վ��TB�Р蚎�N����@:X�<F��~YO�<`�㓫G�s0Ͱ���B�D׃�
�hs���d����|���So����@"D!T�1���N�7�Ac�*q	��-�,�,Y����:�vBk���P������,��V�yrS *���c��(p6�&���w�Pij��H ����Zp�ǫ�%L���DW��z����Rreߪ���-~��Y[<��y�Ǡ��ԏ�c�ַ�N+�eH�(��7�z���X�X95��v-��Z�A��z,o/�$�H#lp����%o�\\�g�R���1�>&��`w��F�R��hB�b�?ߣ��@��b��WZQF�;$``�R=l��݅n'0�X��K����H�';��%0���Z�7)ό�%��>Q��sMxiZ2Mp�e�4�o?�Sq@Q��*�մ_W�i#ƌ�l�p-$hW�@�.�1">0aY�3�\l~ ��km<])8�"���*+L���=v�G�g��`؈ �1���+w�V���f&�8�.�J��G��k��
sȹ�6�w6����ɂ����3�ʞ�b)qE�!�e	�$�>4���Bߞ \��é1�r<�6�l�vW{R�/��d �5B�^I���j�!&����<�>�X��0����eˈO�]v"S���:(|dY^�omr���nN�-[!�tC�6�	0̸a�<<܏������;�I��<�v�|Ĵ[��KE*�|���������_�T�8A��Y\�Ff9�8��<Ky,��A�{%T&����K�������V����ӓY |�a�y�gPh����bo(�#�Ü*����M�m0f;��Vt���dd��g�;� ���IbfPga��dӨ��������'�]9y��<�%��_�g�� �u�7��Y�c�[#0���b-W�һ*��'ɗo�P�@�]/h!m/�����/�5� ��Yf�U��G���f��S�έDF5�L�Z�t����Mxs�M�t�"�XL��!��#Ӄ)5(���aB�7se�[cg�PX�DO�6G�Q���'Y��r��5�>�[�)v��Dn��qE����Ӯ�h_Cg���.4#�6l�*Q�g��(��WHeAagi`��=�0i��N�c�.@r��f�7R��Y,�{�i�`A�a��$Lt�e��T~�u�A��_I��"[�&����ͬ-)��M�x�eu{B����m�� �ZI�-��@�^�%��.uz��3�{t����祓��rd��1��ǒ!��㜘/����@�U@�7E%K�����uW>���FJ��$�M����7�KroWa K�5</�V.���'���C5���ze?Nŋ(G����Ee���;�	��4'�$ �kڐ����|������)�����"@��wh��Iy��+_��R�=1��e��-�9���K�b��m��*��e���a�L����ct�Ē���l�e�ڙ�W�C����3&=�I���)���z5��M��v���yS�p�Ñ$���F�s�*&�v*r0H����K�s�FP_
%v��W��L6���<�Ff�ō��6��)G�b��+�F%���M��CC9�& ��i���휳��~k��@Yǔ* `�6�Dd@ώ��7��K�$�Tda48��˺ɟ�f���>���a���SI3��g���{�C�R�_4;�V���+wC;}�tg�a��R|���ݖ��5B�x��1��#���$A�@�鋵r��������f�{�����o���wܜ�0��r�B�̚dΥ3ˉI�kv��>#=5��L5p��˹K>�N��k�8�Cwy����EcP�ɞ��{ ��t~�i��Y�gx����`+t\Q�%��`�y<����K�AB�Z�*sϴ��$���fi�rXƿ�l�5(��3ɎT���-.̊�T)�ё�~�(�ѐB�V�Ua��:-X�����8���?7�}�n0���A���)��l�G�('i
he^>D[��9����Wf�{�-��Ë2}�qY�ý���x(Q-K��?���P��@�/V-Щ�(
�0�sߜ��b\ͨ��#�:k+2�EÔ$,X�>�K\��؍�}�\85.�	�Ybw��'5�S�ű����F:k��"7�2�����bRƇ\�M��D���j�4��մ/��D#��h}��z*�Iz��B�3�_��`��`�m�i���Y���q�S�5�R�����	6�nz����&� *���/�Rs�˗Th)�'tr��L%#��]@B5� [��jKk������^#�,C�'�_���i�l�$
����Fy^����S5��|�OfT1x����\�(�4U uU٥%�zb������ܬl%�c�����Gw�~2(���*�e��e��@9��f=%R8�f0^G:�<�q�σ[:t@M<���)¸�0�#}]�g�`_k��[���(�[ש���Q4���}'8�F\ㅟ�Mz���5Qi��4�yD��\i^�E�n�ͼ�4i����7��<^�<�C�[?y��x�|�C��m�n
����}^�s-�P��+��ʹ?c[����m�*�"2�b�B��¦Dd�+�B����J�������p��Nƀ�"i�ɕ��F�u����%B��e�7��漣���}�n
����?��r�G����B�K�"����Vk.�BW��^��0��l0p��1D$����_�"�ʺ����p#�����;�
3J�]����m�S���\w����Yu����C��q)�>x�M@@�����M����B%��,�>D��,��s[K9�?�,:��+^��L`���	�yܰH��o����e�,���^m�2�*2M�G�C�_����(�:H���8����v �r���H�B&2`{�M��PN<T!�e�
�S�52Q����R. ��˂�p�'<�-7s�y�;��q�Xq�W���{[-&�q_�]nHEP�-�O p?+� fHKW�M���� ޢ8ƙ$|�e�²�fl\�������(��z{ռ�f�;�2�@�@�@o�	�q��Ke�Ke�����tј�+��8�t�#z�"lo�RHxxt(a�l%c���0Uv [I��-�pEL~�����x�j1AO��k\�>$b$��h�q�8���;�[O����]nj<E�^ʟ�?�J'�m���`Kc�A|3�����b�ckIzcgd�J)�H�H��mN�z�Qe���DzHFa>Aw)�p"N�uu�]��v6��0o�� ߃�t&�~�9O�u��hs{�<�D"�ܝ��	Y��SU4_ �����6�蚳�QQ܌L��H��D痛7ޡ�ހ�j�����גj �󧽊g���Gcw���e�7���Y��Q۝��S�����1�1�����^	����z[�.R3��ދ��b�"�5]���j>���`󳐺U���m���d�vU��<2�6���}��wj:�Et��<��]RX;`7S)Xjc0 ���R9C���J�)]T��]�λp������ק��=��#�|9�<�j*Z�\{���9m(�|�G��[v��G��4�e�;�dn15�t��P�F/r̈́�a�ei�֑-a]~Wc� ��y�)j<���6X���o�S������CP�ǜ(2��$:A;_���&yν�E7_(J�h��#���ԋ	ز�|Ta� �k:"b.r,Z
ْ��L���.C7R6U������;'� �X����0��t	-o�Y7K���6 M]A��	V��
�xάܷg*ff_��S���6u��f�I-�D��)���쀦�s�Ī�#0��u�81�q���$�ȧ�.�s�7��Af��P "�T��;̖v��W�r❢}c�8��Z��XQ�j�W�-�r�t�N��yP �nJ��8T�yX����*0�
����K����?)��8J|���ܻ�&`,[�68T�7�6%�<��jk��h��f����R'��;�K?l���{��*�����)'
hwz5��x�X�18i^6���Y���O$��ew����`�O*�)pL���b7���GROm�VÉ
V������G��mֶ^�(��������H��a;4�q�XL��ꂍ��� 3W��.���m���I�4
5�|2��X��i4�c��I����d̒�[Z�J���|i�S����򳄄i�j<��:�S}�MZa��[h���O�c��&�nN�!��8����h(7ʉFO;��H�((�?U��
��EW�E6toZ`�ފfH���2ߴ�Udژ�k-�%��"��t9�0A1�1�q�#���s��n��T���.�fH[f �jj:x{ �!��{�����ɀV)Xk�ev�Z~���g.y4�oZ�Sk������}�~(mT��q!L7��,��+q�i>l��
�u34#<>.$}��3_$k�~�π�4n��(T�S�İp`�+����n���o� �.�!z�%�E�J8�<eE�ڶ�=_l�3~��:���{��t�T��;�i\�p}!z���RF�3��P7�Dz���2z7P5�m�t��W4����}��as�"��}�Yq�2*Ket��
�~(�u}�1T�e����_�!ё�4��W�����c�.3��!�*�H�����+t���UI�^9��x�}��y}�YCZ&D?=gVGN���
@q�Se�2M3�	ӻ�D*������z��mgŝ5Hl��C�B׭ª�v����_��Awq�i���Cę���F%�	N7�=3�n�����'&� �2���̖+����1:�	h�c�@W�ȍځ09�/	�d�p]��[H�T�e �X1�?\	���U_�*6�7l���e�Y��*ӷ���RV4o�WA�ьZ.t����E�lWAt~�,��Y�g��O�e��:ߋ1M�Y3��u�DIe|�B�:$�~��O�?��ry���ny_��G�[�?N���@X�fظ��. ��^�F(,w�c`d���O*d�%b��ʦ��4{�4��ӛ�b���HK��Y;�0V��X�#gʡoQ*�VĀ�u��}�
��p&�P^���t�iK�s�ũMo�iY�G,�_�`���!0���j-��ޅ���~�|��4O�	��T��9��"����N�Uv|��������vM�w���p���-�L�	��o6 �τh��jQwJB)g�2tD���N�^>K���Τ�w�[�0��"2�+�}o�{!OX�t��jԛ�o�����?j��G*��K��U)��k��ƶ�z�lF�7���Hz~p`%Q��H�4[=v���	�!�P�;V(��U�LsEl��@�+��ˋݝ��9&7�b29� �(FT៪��6�iC�l=�]�e4lWWS�v ��?y�C��L,$�����X�A�-gQ�����^��)��7A���!��)0pc*f��`�����N�OO2"�[�@8��m��W7�#����&s4�����}���\z��߲ڣ!$'����{��_�?���5��]?m~RLz>Ri`��e�Z��z�6�|�Р��Ve'Y+4��	��s{�}ܸ��z/旾KAa�M3�[����6����G'B����:��.$͠j~] ��~\�/\�Z�WUy@�*Io�ث������̰x�CܴJ�w/t�Z.��*��S���U�������{�sp�D�%׿����A{��~���D��"�E��^��~�5���t�j)�AN7:�V���)~�'����2�q�,�
��i�`;s���Y�u�#~}k�-��X�@���iM��z�c�чu��}<�V�������OD*�^}�����.1,ޥ���A�*���.������@/���ؙ�פc�Q��<�3�ΰ���[�$�g]�q9��;����'��(����������iK!u5 ��=�_���ma�r�k5ŢxC񮩆�Íg�6��_6c3�p�bO�	��6$��>���3�v�tYl*7��l��%�%�S��ӷ��p��/�3�-��@�J���a��Wr2 m.}�d�0#	���|[[�����M���e�@[�e���c�b֍+��&6�Vh�?9�raz����k���K�N��J��㿊?,��iK��/�:<͘�x`�,��~�<����*�1�e�}@�x��/p"�����0;L>�h�B��n��-T\�24ZT�^���I�s��^��%���V��|����l�+�}f�G�^$y>J���-#�x�.�D[�;Y�(��)���b.��ME��.Y�}ٯD�Q��G�/�Y@�"�3���ֺ�ތ�ަ�ƶ<�]��ˏ�(��������/e�82�3��zE�f*yl��ۅ7H�-�AUp�ڒ�-��ԑD�"G/�����L�3ʿt�������.���>f��2�uX��xQ�(��ȱ8�,��CF�"�N	��k���2؋s�l[U#b�葫
���a����"V=ub3*��T��|�����O�L���~?+z��
J{7x����I��/�-1X�ஷ�
k�{.F��[�-)�le��V��(����Z16�£���4����F��z�2�=9�ߗ�^�י�Ul�]�t�IU��Uc^����(��2�,[��ޙ���.����GH��S?z�#'��o����� ����m9:1.- �I#���Z�F�Fȧ�����V}�}��Y�]&җ8r�Ou�����w����q)�6����l���89J�G����4 ��z{�]�= ����me�ک�Y��w�ۊ]�u��N�����b�Ĕ�]��H9w\�;T�ۺ�B�jQZ��|\
Z�·Z:�y�s��������cEeGFk.��e���>� ǌB���(8���%�_��Kh�1ߖpK�0�ɓ7
����1O9��Y��ِ��(@��y��l<#�F�l���E,������3R/%�G3�D���&��=^>nq<��*&(���ٞ0��Eԣl�ƈ�Yv�F\�}Ȅ�����L<��o4�U��jqJ����꩎ ��|���Wib�5�����V(���O��c�N���?pyXNd��k	�k��?�#���;��v��Kڰp[��7��&�{��UPOM�������� ���sYx����C�Bk"��1��N� ,[�=h�q��X�E�>�%�1l�?��o�P%���/L4Q�l� 6*mH��3�W�^x0�m�εP�^G�F�9$n��{�!�	�A[��NM�ڂ���-�~RdG��R@�x����U����P�0���y批�7}
�����յwo�I�>��=xz���R�7��HY��a�C����%.����I���K������6q9Uؠ˃�����7��D{'���ݡ�"r�@���v.N�Boz��^C��е{��b���Lf���:�c-C��C�(~<ϏsFvB�u�����V?Ǿ��+�����Q�1��,�Ѭ��,F��j�!�^^\�Р�Hv�sV�0b���z���Ľ-�8��*�/��qo��#~^x����j���UbRT����ܥX�+�~ B�78��W��j�Y��?��[�|vN��;T��~���������/܊�����e)v�Ƞ�~��{3'U����("�2;v�V"���Ǔ7�la���lq��4�����k�f7=��R�/5��G#2�EvM���fu�t3�s�}s�7����D1' �W���u 	Q�Z�~�[�I;���H���#��Uo�cʯ�M�~�f���}�J7�6���-Dr�R��Q���C�W[%	mXK	#�P�N�j�RcQ~��bM�kK��f����x��z,��l�L��<���~^%8u���� zD�"��-
�1!2����!�:*D��R���v���pI�t�͒�{��	��]���5[��}�'����dП}",�	�0��ŋ�w��df.s*��C���N����@����7g�5��W!�E���������k��],�� ���.*6�=y�щ;���ٿ\8��-��]��β͎�w�/r����Q8+��AD�\�W�'ʝ�z�{�����@f}�kR��Pq����ZA3��A���`�R�3m�ےqH~��o�^�##��-Iˆ\�V��Pܶ����3>�dP�K���H�[��~��p��w�`P���I��WX�Nf����94��v�Y�9y�B��7K)cƗ�ִr��PF��O���x�[$onf�8�>BH|�g��s%��-7� �+
��7�M�F C0��e�v���N� g���]��	���~+9�N����}F��?YS(�`��g4>��.�(���'��qcd�/ܝ��b0���{8&�H8X�����7�"�hk����W�@|;ed	�rQ����;5kѝWgG�w��=���ak1��
&�I���P��Lf&�Ʊ�B+�&�2y��`���=��M��֦���j����#��?��|�75ft0����L� j��{	
�q-�P��.�Q �0�xZ�	�m�CgK��-Ԇ��1�Ū�p�@�L���+��b
\ݰ��$��E��V����넆��XH�D�}��k������
�2��6dm!��4^���E��%V��"�t���ږ��5:y����	P�_�%���βͼ&Q[��6n-����5�5�]+Q�����c��D�Rd_<ٍ+}�*~7P��C�H��)��BSTuLL�b�*�ɤ��1�����ͺ���C��u��=-lB�	+�.h��fնר��>�c����L8�>����k�f9�"��ui��Y��d	$���f��F���]��`�lJ.�1uWL���**�t�1>B'����d&,��[�4.)mЃ�(��z����8P�]��J�c��E��h��0��:@��K6�������l{�k��eH�K�_<�$��^�4`�����'�g<s�!Ŧ"��q�1gȬ�2��`�Oy�����:4D
P9~?���X�N�i�s*��D�B\Kb�[�ᶈ�<>2�lX����PH,/��E�{� oп�v��a7��0��/@tJ�,�P����o��!N?@�nm|,���0��m��O��V���ڷQ%���{��ebߋ��3jq��t^"%,�0�-!���vo�|X�y�W��|Oq@����W�suH%v�4��.�,ө�`�g�^Un͖�Z�qk���L��?�1�Fęz|�n��nVc������(���W��nCh�"���S���.��^��q�4��J��ș�̄�����9��=fGj����MM��n�6�u0�-k=^�5�D�tl��������݁w�	�C��͌	����u�ZX|�z�V���=�~l��^���� +�/�.�Z����5*<����zNn���p�@��ૻ�5y٠.�G���������S�g*�����_FJ_��l��֘�U�Skp��fF|�&\������n�r�+.�Kd����R��68��G�.����6�f�ݺڜ\���T��|�w&FV�}P*���|g�g/�]m�T��G o���-��4�A�_�2NO�v�	Y�� ��ph�x�B����@�t��3P�l����<�#ilQ� �&�9:iЍ/�-U
�&UA��,�X,�VJ�2�:�ﳟ��
~uU"x���V6\S�;<38���t���mz�T����� ��
z��	�/C�ʠ�� l���ݣp���q9�;�h�;�o��'�hK|�[n|�i��ʏ�A]����%�����R.������*?�A�/�\̄��/2�c48��ŉ��Y%4p�&�%�1 bBƃYZt�;�Ox�����]P� ��Ѩ�n٥E(c)�lS�uy�G:$��߅;�w�B��+���Y.�o^����2���q���#�V�|�F�sET�����%��r�Ƨ!$�� {��l�ŷ�p�Fc0�m��ᔒ���M`�>����r�mS�#ř����3�pV9�9�$�7�/��]�ʀ�'���s$� �NjTv�����j��P��M(`�\?�i!݆�l�vxx1%0\W�`J�p���rL>˙ţ�"������>bq�?!ĄP��x�9�bzO���$J/� �%��e�KQ�j=��xn��n���؍f^^
�Wٿ,�$ݭ$�I��n��XO�w'�so;@ੀ���-�K1_I���r;Uv��tn~���Ӗ�mѢ:��F?҃��[(��?Z,fy>��ffBN�:s�eb�nH�Z�[dO�Cf�U��߀Z�����eu��)#hߧ�ރ��+���}��4�]�n�^�=	�����W���%��I�-n,��x!��lYH5x��9�ɯ����y���	�(FaC�>���lþXV�~�����N\ƿ#R��������T��	BA�;yus*�S��|�A�U�wfC�H[My���gÊ[]^��$���g>^�~���XI;�#Fi����ȝY�u���/�D�A��g�D�ݺ����3 ���og6蛲���ɳ�|"�Vݽ1�"ҭ�/�u��-rՇOč�7�t ��&�Vi[��fi`j�}��G�m��0��R���Y������b ��q���a��"Q�cBE�� �	�"�����\VJ*���K�<Q�Y��#~~�MTۘ��������B������t�����pyx�����4vA���i�����u"��(J�*S�f󟏾�O�yx��1�����`����5��0I�o�I���Tn<�!���&�_�n<k��&���k�h.3�L�=_x���Ў�S���G7�^3�Hfm[J�]�[�i-����vQ�?�ݪ�b��q�|��)|��~�i����)������J(}f�F��x:C1`��#k�d����ߪ��-���sby�%�-�٨��R>PN�,�(�7*G	W2�T\��,�J���S��eW��?�j��kqJ����ڼ�0{��/�/���\�W��} ���4���v�'E]:e�r����h�H8֌��L�)�ԙe���_����4�dQ�|�/�LO�u0��#����Bʔ^�{R�ha�պ� �U\&ev��Nz�	��B#~Ze$XO�K��ݎŠ���f�u� <CdD���Cr����-����� A� ��A�y�>���� �(@�S�B�T��-�A�&����᳝V(�iA-z�+��;Yf�Q�tk����C|��6`���%u(��&n�7�?���� BQ�ȼ9U���_��&*Y[��kOWt$���T��h"�bP�j���e�CZ��f�a������y#��{��8�ǀ0F{��&Ȼ�0t,�q�oX��3�/My��!�������{,'�\���x�p븆�4>q�}�\�Kh������ �y�6E�z7᢮��gAo��Y��TҜ�`���(���M����ROԱ[���ә7���Q�QS�b�&Z�5Jkdt���	�X���`V�����R�`��?�zN��z��t�k�mǦ���%yG���7��G��bS<wy��~U�#�W�ށ�z��*�0%ڲ��80��6�h��W$Ý���vn'�"_��g�C�,H���0�\�:pU��_$6�m�ІhP���*��y/� �`Ҟ�Jܔ���9Dރ��3oQ�lV���L���M�[���~D�}C�����\�]6�P�tPE���g�����g~.��Ã�F�#�i�A1#��65��^���@��4���걕�2��Yk���I���T�A�ڔ��A/�a�S6ºx�T��[+z,2�mg)o�M��8[��&s�)�����+��Zs�L,>ra鍆HM�V��y���l�vO>yl��h&��ǚo�"fM�B��];�pI�>��?�q�i�!c�b�n���!�{���:" _t�����!tF+5��=��2�?�jkdz�;#�H���A�.�p>�#�W�Z�����_�I(ֵm:��FgT:��S{T�k)���C��mSC�ԾKH^��^�~�Y�W����;Į�4���-zΆugyn��	U�a'�L2�7�i�D��S�����*��V���TI���!9x�֐o�� Y\dAY��j�	T�G��?cE����o���µl`%���&@�l�%W+���j�e.��{��,�}h���'�����n��*����?���D�`xp�,�j+Z�T��$��͎��Nn]����:]�&��<+���x��o #T�κ����4;��_ө��B\�j��BKܬ u \p�A��~V�X�g�*���n�ש@̤���M{.q:��M�jAG�cު]����Wл��[�s����>!��,��A:6��6��Q�;�n��ªK��s�K�����>Gùr?a헠z�mC��"�Gi�6��|-���H� 7n�/{��׆L���l�wF�@~q�g�����}b�w^���<�NK��D�טD�{0L=���K�ϑ����3�<��{�����t0�.����?�4$%�ؒg�(�ؽ�,���U��^H|�N����i ����N���@/��}�p&'M!�:Jٯ��F��j\�V(���;�#Λ,���=�����hw���{�)�ٳ���:#�S�ܹ󦭧V�$S�A荣-����ڂe״����1��9�z]��Y��M� qܫ��Է���HA�q���o�$�Pk��D�;<�f3)�lpa�%�x�MD5͵wP@o$.#�-��E���j��";�W�����;��+Mw����wA�̌Lu�r@sD��@�g�t��ƶ�!��8%��<��.?|�g�k��3l2����Y�H�hc��)��ڐ��d��_�;s��B@z�C#5{��zv<`,0�:cWZ� S1 !a���ߤ_�@Ժ|t��hi��Kw���������ܶ��壃o���������R���@��Oo���C2�&7�a��&��x	(h���t�G���;�Aw��ߒ�jlK�x����!_.H���O|Lf��갅z�!N�n�Y�Ny�솱g�e� j�GC�Ր�9.��x��30���ԏ7mؔK�^�+�����58Vđ��	�@�	^�!�N�q�����K�y�8L��ܗƕ!g��b���"Ȑ@F1FD����.���@1�Us����5yf̳���>v�N�Lj�<�+$���ӣ�z�L��.��[K�X�ָ��`L/��@(�ט��x�Q��� ��d��vT��C8!���T�`<�y�� �cwV��b�w��eA�{,�p�"�K�P���>�$���M�{7���U����O|:��������$P� T��"��$*�]y��4��砣���b8��ސ&n�d��R�1׵�!ĲJߚGeƷ���k��@ckJ���ԗ�cKɶ���a��+�|�FՇ�f���}O��D	>��o( D/G�ݘ5ZUN�ݮ�q�LW1����v��Rx�t�\�iĭFy�䂳�$"��{&U$�}�!L�N��������Q��T��})g�f��M�G��D,�:_}�����:ZQ�V�W<eSP ��T,X~���#D���sR ޤGcQ�_&����:�}-��Q7����f$���ܰUuKB�	���]U���J6���#�$��N�����-���Y�X�]l4�]9����b"��S��N�K�/
x��4��i��],��Hq�L�R�2t�U��<�$ 7��2`3H�"�I�)Ǐ�U��;���MQ���KPV&	\�u�~ ���Im<�'�	�c�f�s�$Nyv�����F�[㌕]Wum�l:�7���93���M�R���k> �k�^:0�={����s�XF�R�}��L�'٫��
� "��|
"�2��m��/�x�?��fM,Έc�o:'4�;�٪H����#x��ة��Dc_F:�!��oH���5ɏn��J�Q\mV*���#ϣƓ�"jz3��R0�5uuA���j#�?j�Z�$��IR�a���&��>��Y��I�Kg^HSw��Q�$}�RzPjkT�
���
A
�ZJ��6럦� W)栲W+	MC��.7�9L��� ,v�S�Y��D�(���(��V��=A�ߖ���ˊj-z�T�.�^��>]��Ec�Q�G�ƨ��0ƽ~)EK�[���Eʚ�M4�F�ל�x�c+F~u7e��&q�/�|Q��� �~�٪j�R���JF����	O�u���T<2�	Qb��N^x�眱������X�ٓg�fc�\�n+&f�J.�Ρpg���V�S�Zb�q�̀��a����;l�u���ݲ��*��jw$%̺��}b�摖�X�tY�F�Z8ϰ^ȍ?�>:��q<	s�x�(���K�����D�O��;g_fc��ך>E��)܊N&���-b\UňRU��A+���9t,2���#�¾)��������+���x�$���)i?��}]��d
�R��J"�=s}�m�g�O81uZ����0Y���g���3<\Q��Xn��l�a�ΘܕVs�t���M�J�U�@������x/�Wc{�C,�%L�'VgG�@����#�C��Þl:�h+��běx[��w~X���n�T�B}҇6������t ��Նn��\��y&�E{�P��D�탫F�n.�L��i)���O�bl��Yl�{u�*}��Uh<�B:!/��9���Ҝ
�:k5� /�t��m�^���~Q�;�{����Y�n�\��yؽJT*�h� p�!�8m"|c��E�BF^�j<���|�4�y�{����	�!h�	��_�r�mwJW��;ʟR�� ~h�+��gW�T��70�oY�� ��u���jh
�x��*��Q����� ))�K�X�q���j��A�H;/���S��\M8�Ba�6��֑����b�Q^�)�t��RE���0 �@��h���Yu�] Z�-�����N ���y�&��\��
���
$����	�&%mH�� S����������Ia6�3(���,`L�
~E`t>��I*���3�$��jx��M��f#��t��q��#������6��;��R0�b�'�'/�)@)��	����-��I@p����:{���L�c�������Զ4�a�4_4^�*�=��\��0�9wN���E�\G2���|U�-C( ѡ?�μo� �喰�e�bĨ�pu�� 
��H���1���Y ��+�V�oh.��@7�Xd6*y�Q:p�M�����E=��GIp�x b�mTYSɤ��Ջ+㑧|(�hE@~��Ê�9����Y{jf��Y�	�Y���o�wے���}���m/��v��JU|V^�ڑ?}����H^�B�����'�%����L�>�S��G{�d֗��iF�v�E-��{ki~�jcU�t�!�ֈ�1�t&��01W5�2���|*�3N����� ���F}&l���&��q��:��iJ"�F��ψ7�L.����n���.#�}��sB��o���%�hm�������#��c9�������\��ꚝS*��Du,�z�;�T�2���a�#]��C�'���٤��[��m�e�v�u�f��_�h=�w��pcxP���xC����E8�ŕ�r�dI��%���z.t�縭̣St�,�6mr�9t<�b 4�a2���-��|"�Ѿ��&�mK���p��D46�_�������9z��/�
�9+�\���8��	��Z�u0絰K�/T���ԟ�`\#�(��9�Ȏh��{"0Bȼ�nn�J��0h_��߶u�bQ8�T���0�Q�t����%��G�lU����s ���N�k�zHJ5)!Y����W�zl*׮V%J�ؤM>~���K��±�,� �G��e�=��9b��:Y�m���a�~:-QT��k��8
͇^��g�qW(%�l�s��U�O�b?��L%���k,βn��B�+�ef��S�{� u���O`����hC>@31�ܫ����u��٭+X5h��^<������φ�RG�AQ��y�;5�0نp���3�R-�J,R�����	�W^�$�q�݋�]��B%j8�U�k(t,W�'��d��M�ƪ���jGn���*`&#�1�[���H���H�����Qp<v���8Xt�<10p*wh��P�*u�v�;��!���8�Y��C��Ҧ*�?�Hjh�}�^�*|��B���Q*��x�Xp>9Y��'£�ؐ>[!�EG����5!Q��:�r��)����B���t��bǧ���@e�\�P&�|?D9/1�̤��z�Z�&ǩ�#:��A�$�-S���L��S��	�\c�� kǼ�q�o�f��ấ��	z����r-Ǔyac��f%�W��֭��% ���@����'f�䂖V��Jz��q�}�&��y�������Nΰ�9���
������b�o�iI�f��.w9�|Yf�JcS��������:��n�:��n�F3~U�/c�������U��elW�����j�R���L���K{���G��/v��aD[�m����.Q�j�P�(ó��#��)]G������Z���V�+Ի#�td�Xp��[M(�ןΎ������u+R����6B�_%�D]m�~b��9�B/и������ZW�aa�4D�`�
h'&5~�OW�z3&f���V]-�uY��.���l���t#���"��Zx�}�)�l�><[�w��+(�9퇆�#P���뿏YeY�c��Pdʲ �2�泻�����6�@B��ߗ���W	Q��ִ�/,��|jP�E1�
�N��U.��V��$*��������q����!͠��F&2fLugQ���?�"l)H�D�V鳪U;�EC2�P���� �O�'�w�ˤ3;�������ӯ���"ūi�N5�xԵi�I�)I�CGk�2i[�wmA���r�(�7�##�I˞gm/��oZ��S���-sEK��u/]�W�CUrR�Gc|�1�A[�me��gy��`�$O��jcH�����r!�9ܩG�Ԝ&D�oT���$h'i��AUKx%׭ɢO����SO��7���ӹ�+>=ʏ�4E�+��+O�X$��X����S�P���3���>�#��g�#Ը�1�_��X�m�*�Utb�D:HnV�(O�A����ì$!�.hVi%09W� ��]����9�v`��r��sޜ����H�Ќ����Ł>�wv9�U�UZp���|@EY�G�AEiL�=��)��T5���u\�� ��&ǉ��\�6e""t��šI�=o�)U<>��y��}:�~��X��t��ܗ{��H��t[ܦ��!h�V2
xR��ͳا�(Ii��B�&ux���H[��[���&+u��
��:�խ�P��
�e�� �7*8�
���T���	�^Xs>�K� �����=�bV�p2�� �!N�>k
/�'�f����S&8�	�?��g$��_��J0#)}��,�����"Qu�7f��Aoo��:ԗ�h��&q�r�(E�/�!��)sM�M�?a	s�V���=\���W�]@*9��O+��J����%F�ϙ���)�u�'L�#kw��p�0��I2{�xlQ�=T��b��*�g�8ַ��-��Fo�H���OC�{e���K���
e��^$� S�5}����@�F��~2�D��4���Tz�iF�ءy��C�0��ݺ�V�h�9!�iS�@�1cb�l+�9��CIŅ �,+��+mGj~'QO��u&��OÓ��u��la�,�u�d)�M�ֲ�6��W�f��c-�r� m�h�0�؆�e?z��}v`�^�ػH<_���ȟ��h�	���|�s��+��dPŸ��|��	ѻT6IPpe��/jn���+-��{�Z	�*�vB6<\�t3ϝ�ש	�5
��N��؀>���[ޜ�l`�������VW�W���X�w���D)��޹Q3�S���H�����[`�Y�I�,�˼���i���_zM�f�yS,bG����a�mjC^�N['k��⢫�brr��k��� �]�����þ�"C͂9[:�t�K�(�魇���a3��EVw1{�~&�,�q�1���H_,�� �kn�`�g c�&A��b_LQ�Ǡ�A�/I�oq��]bn���QW�0狵��K.��/�w�#��K���$H�k9C��KZ<�qCB���Gǅ���of��L�Z�3a� =T�����\�J��6�c�S"Eї���'���ق1���7��P��2�"{�cH�cȹg�XeVn7�(��q���Y�ח@*٘(����M4"�y����M�j�?jz؆��0<f�L�\�^�ћZ��x���:�a�U�̂���.���r�N������OP�3��ԯb��Y���JB����fc$�A�r�բj䗾�h5(��O'0����u�0v�TYBf�sHc���.?9�辍��}?�W���M1w��Gf�"�9�N��`��S-�񞡱)�4�*��cEG]%J����;�����f8b�]��U�j�Nm��1[S�_gnQ�wkp0�����1�=��E�:��z�bY%v*���� !����.n^����_\x4��mT���[E��U�rMg�Ek礵����Xe9�����$%p\~l���;�M���ZD]�"�n;�%+���~�_f脔��)��RPz+���N����|���LH��؆���"��$�� �B�ʒ4�?�����s�� ��r>p7E�J��(�[�q̫�)B�w=�9ም�����)��5UޖU%����*}y���C�
0�V#���U��c>� &�T,�삀S�@���І���n�s.��d���C�zp�����yGQ]�>��f�_�S���wۗ7q�����n�����ϛBm1����$"�p�".�|� ��ϊ\ A��h�:KYB��#��d �w���Y`��X������g'��wCV�Q�m�٩.B�@���f<��?�&��7ˀ��$%8�7�?=7��E�>�e,��D[�gBU��kI�X<�V�[�o�B��k�A27ѭFoE�̋7d�K6U�ݷ;�K���K����kѪ�q�o�)�'�ʣ6�`�����NQ�u/��.����/��GA�H2����-It\����1x�R5aK ��s����Zp}�Z|�W��f�1G<h{k��LE�S}p�c�#א\Lf�vq@���V��)c s^�⟌(�gb��:Nw��&���/ݫ���h�}�����E�eD�l�<x�L�?��>#hno!#%�+V'1c���7�Vy����1�^��G���&A �����LYzk�6~��j6����1�W߭��$͆)+�6��ReP�O��xt&|�����}�9փ� v6�HR��&&��s�2�nv�_Pv�S�+�{N-9IQ<e��kk�R͸e���J�����`��V�oE��J�R.cR�R�=ip3�sPd�(濩<._rZ�d��;gЖ�e�䤉,�g�9���zK��u�)�f0�ڶ��!���)��f����i��H����a��\;�^�:_���?	(�`�(�'XZ�9
(��P��5Zmz���B{���^�Oճ�w��|&��uz�u�F 1k藃�W�S��W��4�7%K�vX~ƤJ�WM�S�R]��YYV��]"�欄X������Ӗ�O���{J���y����&�=�.*D�J�H��4��uﯝ��rr�U�y^�*d�A.��y�T�H	�8°x�V���)������Z�b�=�#�Rx�T���0dC����#IZ�}ԭ��l^L���2��J6:�S�6����ׁ���F��Q���4f�E�&�W�]k�}���D����=x,i�ڴ�
Y��Ъ�-e[_j�.�e�m����� �w��pXϥ'��68y�K�o��q���1C	�x��?C��]1���*1�K�B�M�r��f�%Z}D��{&P���t���@pQ��U����Ip}�U�${D�[00I��N�1~Vȋ���nKC��B�
���Z����ۿ�y�D�k��h��Vg�d��)�y����!��_�y�uB�+y��,�!�P�|W����Vojj%G���Rܺ4\��*>uI7�=���S�h{�F��T���&��Ol�=Q#��A�(��4$������6Ĉr���7�L�y[RO�jm��f��䵞��ޠ�����ADW;�^�l,��c�E�"-�����q&�RF���V�
�H+6��Sx��ob�)X�,9��އ�zΆW&P9	�3����n@T����=�����b����*�r�=�hK|:��EL�)�O���X'���C����Z�Ϣ��rnQz��Sc�h)�^O:�e��'ë��#�N�	vu���&V���i$�3�@���.��c�4;� .b9�}'5/o1r8���e`:r��ߧߏ������O��x���O���i�v��
x<٭��h���5Z,���b��B�#8 ̩;��%�T�X�k�௥Au�NCE��7����{�B�AtU��'.m:EKu�V��mD�F��gs�`����/�6�.��o� �=B��s�����4�6z���T:GT^4=�|�.X߽2����֏�??�=-�6⯎���Ƕ�^1(��ם�S��bT�s�ym0��;�����s��A���XiV�
ՠf����|$��m0-칻vc�C����F���`�q��~L��,�㕾%�:Z�+����0W�
�H�#����*f\��u%Z5 Q��V`� ��D���x���Dq�D�b��S�.t�����j35��:Ц*��DQ���R�Q8��������|ʛte�߆`�)5c�
�?Џ�N�[�?�'a��x�TYn/�����
]��.���Ƚ������t��.�iϠ��Q���݌���B���h�s ��-v2Z�Z7;�����#�\`ފ��l(l�*�E���;�l�Ki5�O\u��U�����lDUٵ�t�)#=�0�@�JT�򫕩��N�o�??��RD��Aj 8�Q�)0[��Ca��lc�34���(Yr��G/���0`]�<��T�×����?�3y��d�4��XL�W����V�BA���69�YT�S�A�&g����|�<��qjz{;�~X_v�ô�?�/B�hL�6T<��X�<����-��� �w�i�Гi��*ЏNpl���R��"��Џ�-���rSW�F��tZӄ�G�93po9��B0���e�>7_����Qj-������:W��_�8��eEz��R�X�ږ��^4�U+��O�����]~6�W��g�����FuV����������6R��Ih.���w����2�"0�df���&�g�{���EQ��Ǩ�k )ي�xR2����i��L�feӲ$�Y�Kd=���gX9.0��p�"bcZr�3���BJx�挖zo�`����bl�5*��x�OWG�:�p�zz"Mhw�q���h�%2��v��Z��?�oZ&�J���ލ�]Υ�S}��������+�ǽ����n�?� `�]�+���H_):EЬ):���^��3T����a��*�⥽1H�֩�r������O�L�#�����$Iu3�d(�S�=�ܨ\�Y�軦tշ^g`Ͽ�'uL���	���Ȟ�@K֧Y7s��N��d�����gwiA/�/�����El�;�c{����v�^
�#9�c�����e}{��rz-w�܊>��O��^gr��ӟ���[����^!2��|Z�~ҀZd����G�3̻vH�������'�����GV���0�̐[��":�x	���1�&��ѳ��Q{ѩi��1�1T2�;N�X1[�[m���$�(�9_y?��5�?}�Z1G��!G��ݪ�?%o�-�8 hC�²w�����h7}ӆBQ3�Ƹ����j��+p��y���V��,��)ArY���eu��ʹH�`���r�N��5i���x�1����څf��Ѓ��0*ئNWJK�7�P,��Pb(��Wj��T�=�C O)��8y�ʲs�ǲ&�`�~n�rr�n��T���~�n�9P�K�m�y� "E�f�q�Ew���2JWv�sƻ8_��v?8�xg��Տ�LW�ڔZ,-�$VrV���pe���+#ޓ���S)Vz��Cj�x�s�%i��'t��(պ�bU�Fl�a�t�-��b�T�]~�vOR��\�i����>�K�j�Q�3�=�q:�Q��= i25ū��!HU�����oR���R�f�+�\w�EJ���Xh*���K%p��)s��]􀢭���u�y�՛��x�h��H�� -��R�L�aW_���w�Q�ѝc8OM6�|2����Wt���3Po7�����f�%>�>�!ƭBf5cfG+�sxJ���s;�d���8��h����VE9��C�1c8��ѧ6�s
]�Vu�T���w��za�y�fM����m�	�8�ӑ�to#�0HM��;����K2���YR���4�ܗ"�0���}	n��⊬�
�K��.����l�?,�+�t-;�.t�ウ��(e6^{N#2>^꒺Vɗ�3�qڜʹ�����6���k+
��م7g�������o⑽�vP ��.�*���E*[��L.�V�ϐY��5�ɡ�r<4�
�d�P������%�Cyap��t�Y �^` ��w1M�5�3�@�W�G��k�j��i�Æ�L6b��lTs [��
��֬f;1�p ;������u��#z���Z7��@�+`&0O�_rNc��\��u`�!�$ڬfܑGh�˼�����[Phq���
�>��@ ޤW6�)�뭪�Z�Ϫ�k���H/�?����Z����*9S�A"'��GA���4�[G��@K�R(�����#�!J.��_��9=�49>D{*"����|���C����._��%��D$�cH9
���L�G���c&0&��=��$�x^'���mvs��\!3=#`z M�CZIӋHf	㿒Ɇq�cfRv�|�!)���I<������f�_P���J4�}q��:��e��Ų�|^�6�g[�O���\$� �<Hy_�%���!Q�|�exo�S�AʔM����UQ�&A����'�3VaH�dT*"�2.\�A�d��T�.��+F�P��i�>��pY0�8��c�g�\��W�,��n�rO�W�Ψa�?����	s ���WnK��)͍�dr��Zj�-�`֚@7�H�bqb��|��'h�w�r�L�T����vs�3��5�o�O��G�����~�^͹�\���'�XPC����"�.�I!z�n�=���6�}��2p"���
��mZL�Lb;�^�m����n֗Sׁ�<ؓ�-6�hIC#���Dl!T��i�T�����v\��5}��C wV{��j�Y"UO�i��5������3��#�d䉩U�[�;�|6�}���wre�0$9�w~"�u��w��MFI� 4��ycx�4�`<OB u,Ao�
��s��ŏ�%& y�h���}�i�|��3�������	���6#r$D�B{��mlNE�!���v]�n����6}�<�#S��K@Vs�E������/~io�Y��W�f,l�l��_��`<DP��ᳮ���ѓa�;6s~t�	�� ���m�ܸNN�<�x��`���˳���6Ph�s|�"eP��b���C�S�s�|I���<�ȋE���m@c�y�B�m �Rm-��WYXQp"�!nG҉?(3��l�+41^k:~�W$�U`_�Ԑ��#���t޾�˃������!{%������)��� ���EJ�-��\ 5�{��g���~�!m�4�q$�9w�L��*�z��ZKڶİ�P�7��V����<5!�Ե��������%̏��,L��`�/����[%�}�X��5�fƆC���{�n�X��qo2�f��#
W}�|�����A����@z�jl�B�s�컆9�%c�t�W �⨌����h5�F��)��<�g��J)�;:��5�<��Mu�Lw^�Z�c��X���2'g�p�E�5Y=�U��j��,"���O_���1�9����U9��c��� �p����Vb�0{�t;��ې%R'P�Zw��{��� k�N�/VQ ��Sxl.�D�v�sQu�h:���/�^���Gs70'��������2����$^?��+�:�%CQl��lW���OCǅp������L�$��S�� *7��P-�~7��$��1��s!����&�HȚ�7Np<H��*Yy;��Ԭ���*�2�Rl�X�6A������3�yﻢ|�������V��HR���yM	�"�c<s!�� �^����>�I��0.���Yk�C�<���i�T^0�+[��C�sk�! I�4�T���MJI���J�Cme��+���EF{���+���7>�q �8�˓�؅D:�,�)\�C�3+/��j�G܉�G�u<�|ȡsǽY&��
m��zpl��p��B��0A�'u����_�A��jӲ����˶�U��^f�K��zsE��$���b���m�%��ʹ�i|K�M�,��ɫ:�r�s.F�D��f���&��0��쁕�i�(�oK>[=�)�!-��md��@a��y�L�4��6Z����pf��r<�R0r�6�r^�.Z��K�c����o��И)�3�*8���L�Q�tN�'`��5�{�>ko���&w؍��I��N���P"������sΛW�ot�-A���,4T�ڵ��!��hM~�>���k��zGOz�2+Z��nyĒm9���J�oy|'X�������7>#%����R�`r!.ߘ�c�fY���-n��bT��%PJ���K�z���F�4<�v���Nb�<�-Q�2?�������%,�ɿF��r���;vs���]bf4a _���a�)������)��SN`��qJ@�7����i��o\��7��Ut8PԈ$�EbŲ��Vp��E��!�t��f�e�a�h[����Z(}��q�"���
U�����ŷ(��3�	y�Z��U[7�1�B)�� �.dk��O�#�/�#�����I;7l�=��uQ��|�t�zX֦A	�W�E���&���w
�*���������Q{�x��Ԁa�]VO�m��m�Q0`K����r�dhz�n�w�q��<;�5��>؀b��A���4
�I���>��H�<���d�4V��~������%�a�ayz�5��k�V��t�֕�9�p����n8B9�;o��;�B0 �j��|�^	���(�`��� ۔ (}O�k����_w�M���=�'��}�#U�ev�ɫ�=�hܗ�Y��%�����V��n@��z�`�j�FIfM�h:#����5	�v�^�d���8�r��V.��?�V���}���m�K˧.[�������
�l�c�{�p'[9�n�U���9���}��Q���6��Q��ZC�A
-J�)�ݖ����l3Q�^�L?ve���Y,}���� �A�m�y�$E}�=�ւވ��N8��e+b��Qj�<|��&
.�O�K6����2���Y3��
W���16T=�JP��՞ݵzhŢ�Z1�'ޔx'���8�&/^�z�[��}ί4������h���&=�>����3o�Ô�[�宑�b�����p�e���Y7��9r&�H�����U�5���E�)aS���m����J3����O5��^0�T�v��-��f�:�9�N�>�ZL���ɔ���lo���d�UX?A����X�s
���e������*y�����;�����D%��;a���Z��������=�j:�0�Ӣ4X���%y�㽱{����v�s��8p��B����=�a�h��f!e=��7�<ol�%�e%!��,��+�BG|��\��M	n�B�d���H��^To3�\�@=�X#��$�ƂA>{H!�c��̗��>�HN��~�wd�����7�ͧ��qU�����w�֕.�PJ��R��J*����S3Ob`rW��;��3�`�8QT�;+0����^�� H�x��֊y��Iw����:DO �r��+��#��g�0^Y*SY�Ƃ��b��6�Ο�_V2����2Q�c�M�"l���I.�<�Ŗ{@�&F�o�~�|��}e�V���3b�����,!�zp��R�����.T�w�(��Tba�x.�f��	����}�06��D���wω��{~�}F����u��\�ۤ�nb+S�
\����>I��o�T�9q�<�Ag���@�@��A�u��p���%C� �bY��3%�楡��_��k�����nq����l����)����儶�&D��E��O�\��:-HM:��#"�
YGU�6YXQ�xf��߬�^k͝T�6�c)Ά(�U����ӂ���Y,��W	F!iܳ<7�Q�3���²��>�=8B䙍�\p�V9A�
���[c�%.-G�I�H8���|���6�V�8Ζ�^B�AB�G�f*�`�>6��+D����V���ގ����5�=Ɲ���l�E�R-�9�7r��߄*��Vr��i���3�,�I5�ı�P�sO`��!�Yz�ئ��3���Y!�H�r#��mZGk��΅��O���$������iA�0<���HX�j�I;,�^ݘ+�h¶���K�4��'+�����Y�oi3��t	�ѵ�q�wZ��� Knc_�+ (hf��ڨ�����]��ؕ�� ~��=&��X���{��2�	��d��m�S��y��x�fKH�dgM`�i�9�:������u1����A	���=X
��w�����������_�
��
��Mh�j(�|ck�Y�}��q#�  �l��PR�`�=,��x�,��k|�˷��Zm����ռM�H�f���'��~l�Ϙ�F_n� ��M;Q�0�Ǻ��*9[��`-T�x�<!@�T����0�O;ډM��= �G��5��w���9"U*��bm�����Zrs����W����b����9�h��:��P�Q��_]�z����<����{z��n;�6��nM`.�>8�&���eI
l����}}/��W�0.-�\N�&Ȟ��鑩��ی���m���$!�ސv���{�V�PI*�`�!f�w�3��З((qDܛp��F��gu�r�~&[TB��¨n|$�'ڸƲw*�O�Ӑ�nG�J�l����1u���dh�~�k���7j�O�,7X���4���J��e������@��F�As��42��z{��o���~�]Q`4-�$�����v�o�~��p^�蹤�N�Z�6D|�ܛ_� ���)���r��o%���7���]̼R�i���G� ���di�C���7�4�7�=S���Ɖ���N�[0��`ҩ�?�VH"��b�䚮��>m*^���9���^
�d���ϑ�@e&RL�|Jχ_�8��U	���e�h
M�l��C�{{L�?��pq��[�A��D�ܱ���p��/��V4\b� �/��|��nR �I�2j8e�c>����p�t��&_��] h"(�,�k��@3 ����90I�k��,3����O֦�����QYo����Vr�!�0���F��2�����泈���h�����r�~��on#�>*�,��提��^&Շ�ӌ��%�<ń��gćxsd�POI�V��k>R��e�h��֗�s�gxp�@�d�9��'|�nGZ2?��ЍDٮa���o���$Zwu��MN��=�7����P���;����ʽCes�����ӡ����e�to}
���4�4@����k�[��f/��xz����w��W����3j֨���i��-k���x�3C�
��p5�ܸ;��:�����^b΁��Ԋ�⛰���7���k821,�o#eo1'����~��Mgv�w������ 	���cH>g~j�3�o�r���/���D�IE{B�[[�������\��u]�}����Y\�#�,����D\p!���>ʙ���h�?uD���*��
�܇;V<��,��*�ڎ����.�� �y�j�lЏ���M��K���4�o��nI*j�ŋ��+�@M��>R����2@�|;���g��A���BE�RK�MǞ�oh\Z���	����� ��1�xd�ş�o��#C#�>�PAh�!�@�m���	�� W.��F����b���o.P����?�F�sr�-�xnI�Y����Pr7?U���H7�~����Ǫ둅�xk��U[�F������=C<���cm<�!R%�'z����٘v)?׳^�q�S����w��t<��"2"bۑ�SU�Q�_Y��l���f5����N�ѽ����a�I�|t�����c����U��j��p�t&]��e����Ҙ����
϶�iWw��~eVc��nIk�$�ŐU��{QdQ��Y
�!�� (O9D6�܋��<Uob���w�Zs�Jf`�\�v�MQ��$tau�be.q%�O��t���vC�pp�k�7��
�/쏟!;��a-@��3h���Sh�%�D���b\%�K&nj�?�џ�3�"������q�,,��'Kgg(}mϷK׽�� ���G�5��
��̀it9�AhՕ���E�Cj�ѭ���=���zK�[K�o����"uf�]r׋C�&T�7a�.jp�T�$�P�]��'4}����@C.2"�����4�7��S�#?����K'�HX����]8w}���d�e<D���� n�OD�d�8��[��#������
��V�0#A��=���ʩ\�x��B���/�;�z��_0R��Q��AA^Ag�Ǽ,��F�6Wxk�&����HQF:�b�0F#q���X�5`�D%<��珉��T�L{��v��ԋ���\M�@���݌�Us7��q�7	6*�L!s�-�c'2T��@��kՀ�
�����8,�0��6��ǆ�o��s��
���
1�^����9J'�g��b��kn��h�����;45�@ctElէC�d���%�C@;=g�y�<(0Y�ǡ��Qq֏��8<?Ttr��c���^=�r:�ʗܕC��眂����/k��m�Y�͍Q�����I�oU����i����mO=��b����"���׻a���"\��MPU�9��������q��n�>I��>�"]��uCl��}tο�����"�]rN��а�
��IiB06Z���q��.oc������"�����>J5UP~M!�,��Vjݻ�Rz-������b©>���x'�������3�hI�uN��SH2];�M$1��p?�TY�[�'Ɨ�Ō�L�u�:$&�E��}��=�Dp`&w���K�)�UZ�@���=���V�yҳ�c|'���Mg��>*�hWI�}Tl���G��z�u+���%�gpF_;=��"�2Q T��f-n���� }�ƿ��FKe��=Z?I 4�X�|���`�D?�����mд��t��=�cv'��43�/k*tz�E R3"3@�4��X�X4,$�0�'�}��#��Q�?���&�	#�_6���YT��Z�Υh�c��;i�[ͫFM���Z��Op�J�IvجBm���� �h(����\�WX��ک�)�������� M��R.�2\�q��}��`�B���Ki�|\��O^�UVƔ�z�P8"���ZG��^y�M�ˢ���cn����J�/َs�����Z�5�� �r��h�M��k]����HO'zS���2�����E;�zoXbLV�ӫj���FN>�����
KΈ����^5������R�R�� �>����3ɐєP�؆��hQt`&�v�އ/SS!��C��W��˯�Lg��돁Ǭ���Rn�z�" ����i�E�N�R�bq���$H�L�Ԫy-��v�"��";��� B������"�\�^�@����5X��ַ*�!w�ʭ�g�%�4��K��I�̓��&����f�Բ�H��@6��	��=���]�,��E0j��F�*HQ��@�55nkh������O'�q�1�u���bܘ�V��J%j���}�;��3@h��yX�nz�B�,cwՌ�$�d��@�f���ʃ�P�\6Зh�uX}�,�:� FݪHF����R>�1��p*2��b�r���&h�`/�քA�ǿ��|�0a�&ץW�	8U�ĄAܷ�_�%�7n͏�����jj:r�
p�.&�����b��NXv�;XC3��I��c�{�u�;�e��z#��P��5�p��@N��V � �c"��&MX���DN�O�Յ��	b�?z�#,��H���YEc
Dh���
.Du���o�mAG�<!�siujK�kϑ��b��{P>���&.@���<_w������5�p���i�v�4S�B����}����C:�C�%�^�mY5�̈���h]7	'������{��|�z!��=8)��(�p�ψ�%��nn�R��M�%]�
u
�t��(cRgO
Q���$t�N�����wԪ�*s�3����9ʩa���W�@����h��d��l������d!թC�́F���E����'�P�[u��=1L�ـ!�f���ͥ�[ax�2�uЫ8� �Ձ�:�u{����=*�r��TO�V�`"�!@ǈ����D���l�O�([�M�����-`��9�=�T�Zx.��R�� �&�����p��G���ff������K��/_?�����`z���R�/�����'D��w�VwD'4���]=i�����?�r3/-�g��N�iׅW��i�C�﬐G#]o��+}p����2?��6�3�ڲ�a�C-���y����{{
��@�X�����d�� �.n��WU��MԳ�?�p�zk���P����!J�r�Ч|�g��}n��U�����^���b�m���7Q�r�����蠾�'zB���?�bA��Rl��_bCKh���o�,=L�l����uo�ZW*U9��"�y++�V�=�G:��x�=o�y�͡ȇ ���3�ϭo>_�SOL��{��<���q�����ZW���ή��@�S��3P�5�NJ9�|�Xdij5ڊj�;b��c}�Qk�ҷo;
d�?�y����w�w�C�Ú��O��F���fn~��s2{e�M��"�*���ZZ�ЎH�0�y���wȃ�>:-��G�A�?:\�;^B��$��w��W�4�V8�������ic�KC4��9��k� gV}p��"m�XnJ˄u����^J��H/p�Q�b�o	d=7�8�?��͗A�`1�C��z ���"��x�S�á�]?� ��G���;vm��v0S���0��'����~`�g��K�k��I9fg��#�&�hn������	���9EWmR�l8Z�f�P'���������ަ�m=,�%+�;btg�Ye`�hr;��?/��1�k���^�:<T��m2�������6\P���ؽCb��o]��ig�I9+a��V���F���-���#��Y��*�g{?�>G>�(-ю��Β%5�HV_��Q4A@��� x���E�Ud��ӂw���	D�\	<6u��M+4\"=��4�4�εʚ�h3�D����B��F/�l�A���ĩX��Vzl\)�{R�K&#XƋ8F4�����z���Cz�&�!�����Q�@�^��5�o3v� �jy1��|Tz�S
f�_��!u�*��|����X1�\�l��a�@II�{��k?�G��٭?^ e�e�W�p���x��1u4�dG2�"k�&G���K,���̎uW��?�u�6y�{;�,GƔ`�y��REglǚ�R�m�N!8ϘZ�W�"�M�J)@��x�A8>N6:��Xώ
Qc66�2���-O�f���:��,LG���I���*��Li�(@@_�o�ؑ�$�գ��5]��l����F�����-г�`�Nٖn{�z�(���P}�ڋ�f�5��I�-!'���!�,_$%g<Oכ�K��Q2�P��qC3�\�J	��kIq��N�ϩ-%Ҿf��������DV5��}& ����O�����́<��3�'�G$ɥ-R+����Mӎ�c�Q���D:�Z��l�(ؑݼc�yyu1qP��T̅{H�,d�'�4�f�n���Z�y^B���>�bcJT*k�Q���-�Us9xķ���?� v��d�ű/�/=)҆��BkDd@�{��ý5�5�g:�Z0���m`�m�ܰ�P�����i�����;	��kn�i��(A�`�`���t㪬�=�G��UI�kF��~~h�����pWmF����#���!|���Ec�\4��O����_��W��A�	ͥ'���!��ft�ٸ�HF�)q�9n��n����#B{��%�A ���̸]�9�/`�D_�7��$���bTo�K�[{5|�1��d H���ā0�.|<� ��;+e���� �&��3h�YCS�1n����*�vЂ�G7��RS��M.Z1�L<g�A֘/;.j��րD�΢�Ă�2��f"3�iz��1p�)��O"}��x�!U���3g$�j�6� ������#S��v��B�R����ʻ�i�������Y� ާ�A���m�u��:HEȫ&�ڽ�\�_j"�1ϵ�K��Ȧ� ��H��]Hk�����y��y(��CJ�u;z`(�S���07� L[�W�rY�G��
��0�T��RV���<C> ��-�(0��t�ox�2c1�x�&C���^�;�YIVy��NRN	C�m&��f�����j���=�����4b�)�[����_;��M�Z��.�y�ۑGl)T���4Դ�*��Y��&��41g�i}d�n���>���?�Gо&�&E����/ic���:Κs����\6t�8q�����`c�;LӁ��q���,0-�8�h��j`ɾ��*ry�e!e� 1R[-�c!���Vj��;��/>|�b�k/���1�(�;W8P���}r��K���@��%b��f���4p=q�K>
kN�<%Cw7�,�"1o���-讒�$@��؛cp�#�/�5s�	R(��kRR���7��aw�%�f#�d�þ�����{&rmq%�p|�=d��3����w�������iqt��,�2����)�%�o�����D6�0Z.!��$�;�dd|��|ۄE����f�����P�����ƶVIE�qwJ��C��5����Đt��w!P^�pJmFU<�	׬�d�iT�P�C�4�}������V�X<J�M[�0ַ0H�_u� Z�og1�n��1����Y�`;���3����w�z3���3Q�0���wG��Ѕ�e�Q�E �����	M�#ǽ'�\֯!p?6F,��Br���"V����k(�q`��T�5�u��� ($�{�ϔ��'|��- އz��Ի�&�ܜ�����p�1Id	���Ο���[9�C������3��y�;���?K������?����X�K��@ؔ������+.RW��Q�����[,U-�gi�����X�Z���[ɾ��W=��b�-d������.En�J�m�H���"/�
-���N_,Ga׉���]�TzNu��rPت��o�,�����s5
;�U`����(��
]�d��A�=��V��}�["Ȇзw�#7���