��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�+����Rq�����������+�nS�U�F7&���S����"�M ��U���@�˴�5��.� -;P�~�oa|
)k���BЖ�@�o�v�4ߘ<��4�l��D�4Ak���-.b���mC*��D�i�M%��%�k�~&ʳ��0!����nY�qe��3��ck����o��z"��,f�ը��%$���|�;+#�0f�UhOǃ��2刑�Lc�����|��|����Q��Ol�pf��\�4Y�
A�Y�a@��qnNAz�pד��ݮiF�?��'~&{�X�v����H�	���Gʲ���dӤ�>v�� ���K�B�x��X�[#s��W�V��.��f$�n���:Qn��24"M��<48�}[�� �(�5��t�L�6����ئe3Xa�|=�X$nD�H"ď�Vl��⼞=��5��n�Q���6;#٬"I�L���P����/P=�}�㟂���C���?�ZI�r�	5��]%���ē�2FTC�Sh��Ds]鉬�@�0:�?"ܮAۙ�>���?��i+c��$�vf�:��P����LX�Z��+�'��Y�}�G��)��q��ʋ�X�]���ۅЅ�aڴG��i����(ް?	�P9���y�
�����E==6�iS��=م�gU����!��8�د�§���g��d���B�Rx%��E}��8�!-�U��@=�R ��s�/�ǥ�;,'�f��|�<�\W�21u�a���{-��������k�����@b��G�9SK{[O��Y��7�vb���yS�����	�63ǲ�Sr�,B�/�t�(��� bc";W���"-�����?�1\�ؤ'

`�x��4Q.�H����E�l���5��S���kd1��{+Hڔ�խ8�|$�������؄+����)���gn��+砯y���>3T��Xw5ӗ<,�C���   ̰�78ys
7�s�m�MO���_���t�3���d���*�۱�)!܃�9��-�J���.��qkT�*)�
0�Fx����t�g#@p��s���(��ܐ�q��U)ײ�Zƚś�!����qp� }�̚ޒ��	�v4����l�a�+|Eۺ�m�%��~�K~�u/+Em����	����������O�����閐��q�p�4��H@n�� N}���dv��m?�:�>!���GK���7r�H�0O��ߙ�	�N,���;�XG�Hw���2�d�lD��
�ϻY>�R���`������R�i�[~�~�<0�|�8t!��l*�,p49Ọ�2Vj������N~EG8��!S�K���͙�}IjV���l���1��Cz&3���\'(��]AG�0Z}?���=�bLϛ�A��3%�$�[G�j�fuA'�ٰ0�q�,����\�I���w�%�7pc�/ ���'t|�M�-�X3U �������fܨ�ZI	�:�:͙(:��}$@Fۢ��q|Le)Q�>C���ӆ[�1���E=A�	��j��WQ��;9�L�S�V����X�,�`������DY,�m�?��!!vC�yu��Ȣ%������S!G=3��i �t�2h,q�&�"���'+t����L�G��_�/QNvsN�UK�@+���[#��yfK�+�2)��/� =�v>3�(>r�'�(Abz!8{��>�G��Y��ϕ���5�
aiY��%ZӰ^#�KJ�7�_����r�90�"Hf�T�F ĳ#4�˟��?��ف�2@�F���Ƃ����M�]>�6Sy3!����=,C Zʺ�}p���݂�<�\��	kI�O�>�~�?=�jXF[XX�� �\)�h�\�v�GE�hOZ��y��6*I�(�ϱJgٕ6� {�� �l``;ʟ�`F�%{Tѱ� ?I�K�^�?�G��V�}t"��V��oń\���V׿� ��{9q_�� �\���F���LJ�����tn
ǏK�񍱖��}c88+¾R�Yd�]���R�2���W�+�Pw`ބ�������%[E�J"+�����q��0� �Ȏ��vML�צ��g֒��3��|��`��&9} ������\t�y9��w�*���k�[��x����f�!��캩�G;�ǻ
VA'�XS�B�g��ҼG������~����Np�*�G��F��|zH�3��t����d�'��Lk�p���1�~'QB��A�v�ah�[����7a�yJ��ӻ�t%-�0ۘ*�
��>(�޹-�=yG�?KK��:K�~�� 2���j��Xv���d��=��|�8Z��F���약_��䋨��8E�;���I��|�j�+�����h.aC�i"��j�T�y�F�>��_qS�,�j�*9eG2ʺ}��-f]g殺���-�hGk�ViR��q���~�l�_��WX^��"����{f��h������ԁhQ���×���uC1���������������6���<q��L��TZ�r��|�&�ҫ���|}FJ��T~KȪԅ�_��H�-u�x_8Fg�<�2���Y �CW�tnO�HZc������}XD���u����M��r�!
��pi��R�����{Q���
����ک5;G�d�Ƽ�'Z�%�����\��5B�P5��*J�{�r���N��J�vlF?�/>�V	��Rf��)�2�RX-���}&�Ө�AH�t3�����Q�/iӢw	wۛs1N���#*_�U�A��ڂ�ہH�a6H�^�Ѐ�}����Q
FQ�2%�c�T�������xD���#H��H�}C��K�ܿ<�a���-�0K�#�����@PȖ���B&�����A
�@g��~�^���XR�E��Z�'�=�8�v{���Y�^���"(���2 ('�a�7�ƬR���r��9���s:��<�."��ʌyP�mE�ۃt�^�g����y~�H�ヤH(3)�k�9E�J^�l~O��'z�?��v�I���LJ���<��>�?�k���U�m���pцpbV �#���~hB�t#$etU�m��r5l�l�5U�v�(_D{���q�����7��˟=��2T�d�s�K/٪7ԓ�^��� ˠ�?v�jץ��)Q����,�ͽ������8��9��q��v���H�͖҃0��L�-Õ$7���()?����n��P���7Nn[igx����ȡ48xm�ɴFju,/RVu�0���{k��̙���?��И�}Q��ے+9��_t&�O?e���K�)Fa"lx��&����P*��e�����"�U/1���Q*j��0�Ö��"_�ֹ��goE1
l�P	�ދ�걽69�щ��	3
4����ﭙ)�U���T��H�dҽcͺh�C_�t����,�,����4��)A�f�=�d���\���x9	tWU����h%�p -<��˷�7C@�f������k7`ڋy}�!󃩊p��窅���V�LO�6e0���V� �*�Y���0ltδt��74�ϏM��j
*"8Xkr�e�)�W{5�#�+������M���Q0�mSZ��8�{�[��kܨ��h��N�/�;����h}Y�)_�f{p�o(@��������c88bUej�`o���|�,�#�P�&��9���|�Oe�;���4	�O�}�ẎB ��Ԫ]-.�Y���A��_A������2}rO=���R��&��g68l�6\�!�n��YJ�О5�q�t"�tܣp;�t�ctд����i�����ԏ�
0v��%C��	��!}��)��ͫ'L��q�ɿs�����d�6#�4lr-�}�m�뮭������B�{��ON9v2������׀W��c�����.hi��g[��i"�Ш	�q�b�Ct�
��s�|�A}(Hs��(��p�R@��ړ9BӠ˔�]�`$�-�K�C���;ɹ I�;P����x\\Ȣ��*,A����j'�(���N3�3֑�ǣ�jF���]H�&�聪�:B�I�
9��L��U5�.�F�%xD���1�Y��A�۶�U.#�I/p����D�ף���B�JQ�C�
<�/�y�����ܤ����|��r�:�~z�G��_�MO�K�m��i:� 8θ.�FUo��V�'^�ꇩC����9�UM;���^{�������˺�E�Jmh�5�]��}�{#(U�1\N�+�`~�1���~�:�SМ�B�>��HاHB�_�uЉ%�1�>�5]�w��rHD�V�c�egeI;�/��6&98E��b�e]q���H*�$ѱ���{I���\�dhI4���O |�ś�t�uӕ���	���u�Ղe��.�?�ڛ;�.	j��!$f ��0I����R���[�#519W�/��]�<	 H�[fhE4�Prs9"J���F�B�/��|᭒����an��L��
4NV�(m�ݗ�:s�xU�}�쁆��W KK � ���ޯ��['>��9��:��_�VV��/�Z_�EYd�M0e��]A!/�m_C�����z�m�ҽB��Z���q��(,L�ˉbj���H
�������B;��0�Ă�Y��p�=e��9�
乞1:���X��lj=��L�IR����q�q����=�����Rah�2I�k� %�h� ~9�)�������aQTn�)�P5n�~&�d�F�y�j�>�D����v3��،�W��C%��p��Kn�K��\�a�pY_G^�	݁;☽�{:���Ig���[�;2���St�jA~��ld�G�Gd3--z��Ii8�*�
�t�
��.Dؙ\[�"?�Y�#&M{�-�I��V�܁Y#����G7qDc`��{�l���e3��(��9�?���A�x�YD��� [\�8�à�k�ӂ���\ZAH�G���җ�?��3��4�HI�sy�c�P���aӟ���9���dx�%	0︣z'��zm (W�s�.���Y�a�B,6�,�3?9���`�PˊQ�V5R�B�w��#zs�YK�l��}A����*�'�=�Ǔ~) ��AJ��8����q�:O
_v�bK���<,?^�.	3CK�jQ�<�41U@㥑���"n�$��9]�,Zy9D��e��>�H7��J���te>��e���R�T������ٓ��ܪ�P��ɾ���v+�h|�@���Ѧ}���2rΞ�>�ͨ�Tk�h/G��,.���p M��>����8�K�}c�H��i�JuO�p��s8�x�f;�E�&�dj!1S���j�q�p\�Wd��F6�mjsq�&��B��{�������X�ڞ�<|������.OY����xL聙B���w�T�0y��37��ƚ�60M�Ӛ,ݢө�
����Ϗ�G���|�����;QX���}B� �[�z�љ�.7_A�03�e�ؽA歚������Ƒ`SQ{Ԝ��y����e��W�ˡ>X|��[b@M�qg(���FC�i�ϟ���v���@T
X�����K�-��{3���{�I�$NT n�,�qV�����X�QO2��LH>���+�&���k��n���`��~{Z"<�y]7�2v�p��مx��EDG�P	��G��1���x��ʷj���Ȣ����Sg}G�8̃����̪�����|�i�-�"�D�]�F�S1�F�Ư:�5Q��Ζ˫��R���a�aB;�{�aO?mF|��P�u516럧��}y����ނ���uv�o�E�h9��6�yt�[�2>���\��ug'*3�{�b�@���G�76�e��<�t)y4}Gg�~��8��IͰ|7���V\%�W�qЙ��q��M�~�A�1bKu�SoM���M���TWp�緥��7ƿ:�nˡ�Cjq�(bͨ'Q���J����5`����Â^��y���$yA�l�S��jc�Q�8�u����21��wQ|Bt�k��8<�K��
Ouj���IH�7��]<E�sȷ�6��S��_�[}�^�E��:.��tL��QD�]H۸n&,-����g۱�:��J����r0�4ohQ�u�?jO��Ҏ�޲'��I!�jE՞�r��ZZfsgc��aF���Y���n��E�8�0L\7V���]�����:E}�]�&ܨ: ���ǌI�x��Yi>��r����[SsRW�z���L!�9.zܒ�Z%,hFk����9�s?d���`��.�rSl�����O�ŕ���*]߁���I��8���i<��Ͼ�0̱�V�[�9�̹I�-�e�SՁ���]>��+G`(����Q։as	�I��_�L�Y�h}VV|�T��@�B��5�f�|���b�l�0,{�.뭺߰�c����?:T���UJ��i�ȑ�gĔ������*���d-�Hw.�e"Y6ng���p��.���j �iz��zwr���o"�N:�K��ɔխ����1��&�a��n�r���ױ�:y����fU��pU��`-��';�-
���2�.{@�a�kp��"ϡ���8�e����xP��(M�,Y�mH9k=�K�����<Z�b}#���j���t}����k~q��.= $�˧3�
���z��I�Z@��R�c�E��t���	�I���H�џ��e	����)\b���^<�/�dk=�
���:n�|�����b������o��K^?2�aaq)�~�`=�[�0b�>|���M��5%ǈ�����s��H��Q�j����c����[�C翷7�G�6�SJ��.f�c5��?FN*�D_7 �f�D�Qt,a*��.Oºi5�/�T�n��6"�d�38��J���5��/2٠"��Q�1-���y�c[��d@��öF��9C7���@��=��_��ޏ����J�I�c/��i;���>�.L��yT�15��ܴ-�.t
�%�������L*�>]�d1�H��?����!�z�x�no���|�SPL�=���I�],���Y
���?����/�C��J��Џ�(�`�5Gjg�>ʁ.�np�Hݨt;�^�A�9gQ��Qv%�D��Iwt�h�=h�UP�r�����ޯ.>���r�\m�H)��<�����UY��-�S�?iA�� ���@8�sL:�$0[����Y��[�o
f"B�5�=Jg�eC��A39���Օꠖ�ݘ��Rο�ag���q�8�F���Bu�	��j�Z�؅h*ܡJ�;�y�w��@�s�r�5���k �c�?�uW�R�v�|lG�xy�*��?�7��j-5�59dT"s�X���:)k�m��
�T6��Եj�J��  ��@V�o4��;�M	uZ�Xe�^k��R�$(�M=*������[A��(.���t#�;¼XYݧ��O5����'#ht\�n������:�����Rs�->��4�s#���M�(�y ��H�L�d��?�7�϶�����22"c`ؙr�HAg���R��P���w8Yz��<xW|tD��$T�A���w'l9��3�k0dyy�3N�1�A9nP������Y��8�rqrX�����-�G!C�ϝ��6��6Iu�X��~/�(���Bq���=��+XD�0�%[��b�Il����\J���5t����g�����K��b�����-)��d��<;�C�8���y}���s7c���C��0�Y|H���!2��w4�9���I]�U�Q����"yK�ڟݪi�"��KH�t�8)"Q��|t9V�A�)@�_�j]��3>���kISձ3��}6x��E�@�=���|����<l����[��H�U��.u%�;q�C��S���2�����5yo�#�M��p���{cV����+N�P����y�?�J�Fn�H����tj��T��1�O!�����>��`5!�r,E��!��E�oC �/��H�*TL����0��� �ϝ`���_��ck8O�c��Q����/�Dsw|$ҡ�&�T�/>t���b�U�����Da�u��;
B)�ձc�6��m˻O�m��#%.�T�8����Ww�͂ն>�[��icx58"ij;�??�y����.���p5ɲ�2J��L�e��ژ.:�(/�
������
��ذgiJ�g�'��Uǲ+�3<�ރ1�hϗº�-����:�y\�y������A�w��-�8X)A=߬`;�ҢԀ6���L-M�����=E�>��ݬ���>��(V|���C��l�����`���IZ�!^y��H;.\���̚:d�%ȟ��}�}L.�ƯY�e�y*��V��3�_~32��7k�/�ʾ�Zݼ��g�1���������'�n�Km}4�1}���Ê!y���xf3���^���Cm��B�=h(���R��).p9��]0�H�>�,������"���w�惻�pt#���"x�9TC˧�ۍQ�f'?;F�`�N����<|!�5�h���� ~�{��Ԕ��[�1�|
^��zɓ<�q��@��]�e���x�M�A[�`���1�Jq'I��3 �c�C�q[�V�k�:sō�\�z�}W�]�G�0k�G�YDUǌ��t�0/}!�:�����r8��1ú��� �&��}�!���G�L���}C�y_Ԍ'����x��&�Q��`DOI�c��3�#J�,��[	%�_��(�O�_w��X(-�/�r���2�]�/grB��~U[�M�&D�IW�c?uw�թ%u����1�\�������&Fi4oW����ۘlSI��)א�<��]�&;�P��`r��5����5�K��Ω�ԫ^��Tn�K���q�|���gԣ �n��="���)�״c6�dk��^�~��z��m��cJ֗�nM��
:W��ݺ��&�
F3r"�ʆ�qÐ�Y�
���:-���p��ƍ��	,A��1����3�^�0�����TRl�����'Ca1����Bh�'&n�*�mP����/1�C���O��7A����0�m9\�`���%���|�S\	(X��ewn����������j=��B����`ddW�$��ө�(�}&#�S�D�w��\��챺����I�پ'B�4��z���ԠX�K���@$�'����q6-5�DF����-�X��_bw-�=M6��>���֩ԓ"A�_W{YO_�/�ύ�-5��j�?�`t/r�Ȏ��2M��� �7sנ+�gt��{���F]J�� lb�� �Se(�u�3�� |�.������&�T=M���+�A�����V���~��`��+�sX�QXQ�v@5�/ν�G�)�|�C������6nܿ&�$	���j��``U����
��5��P�C �t�S��L�Ԗ�RIB����d^�� ��~��ྖt�}_TX�2bϵ���������vw#ѮE��*�d��Q��m��?;y��q8Ë��eD_8O�I���b�JW�Mj��='����r�GI^^	D�v�ɬih_���b�1"b���&#V���?	�����3l5��j��k�~�7�_(q^r:q0z�x��$����:"��[�� �:�i��v�椷�nL�/d����y�	�l��$��ם��-���k=�0+����0U�[��\z�Ȃ�ʏ_v2�y�)wَ�OƦVs��J'5'�x������|����5vL
�ޝ���#�ד@�;�FO�]@�"�Fo[����bPmͣ@�9����m�E���[�[{�+��J}#,!� �<'Yv�ߛqqH���o�kH�$c%����ߓd��\�4Pb�@C��h�������ȑ'9ׯ�lhQq�zj�-/��ԥ�^ղf_ͱ�r�.���qƮy�jG��D��6XH���vN �wLN�XR�������͢�E�%�E]�����N}��G�+�DSz(�NF|!EHR�zK�X
S./��솄�@v��)ݹ�Z�陵7���K[�w�yF�_z:%8ךX=�i�8w���=���;}ɛ}h�)�A���U�^�0Sw���&�=0WJ�1����_ ��K c�
��k�z��{"M����E/D�?���m�h��;ξ��Ӯ	N:�fG�Á!8�N����%#���9}���`�g�3��7�q�"���q7����ǧF��tV��[<4�J�>Z�Ȗ',��.�}9��!��w3�Y
��
�mC�v� Xy�$t���{��,�j\zx\��p��1O��Ê,k�x�TY:+����G?��z�K�1�����r 1�[:0Q�r�>��Κ���RC�xn<�w�������1��S����(����, ���p>ǠD�Ќ�y��[����(>� 6ZHv��-D=�P��������ݓ{VϚ!�+ �����8hŤl-wrKh��CNHA~f�c��][Bp���>������0�r��b��S �:��w��u�r�{E��l�@ �<mZS}x�����wi�|��^��Ut�v�~s��'��;/Á1kC�eS4Y
u���"��_V!���]w�koO�@�]�$��eF�ß�K���<�?�D���O|��%D���D92}x� ��60QٚNi��mX��ǜ�d%�o��ȋe��Z�ÝW�rc�zz��l�1c�͏ҧse���ժ���J� ��1A��r�w`l_*}L�ei�ak���j�0B�@}Yϳhg_�$�uH�sc�U�=����פ3�l��D1�be9]6s�7ơ�`5���q������䊘~k�
7'��w��wo>�G��x�P0͞y;�/�^X!��RY2v�e$��i,�WR��cN�ya^:�a{��%�s�́R��+T��>dN>�9#�����~u%�h�ϟ��4�-�||�ð�4�	C|DM"�wb��1F�@<)M�3��u ���#8�t��MĖ�"�'H�r0"Ė�ꮞ������)W�u�~��4T�p@j�dӅ�t�5}T݁w�Ĺu�꛾���H.���v�݈/6���eTX��~w�&��&�~���Y�e�
޺�}ں�_4��>�f�tf_� ��c�-�*$��zG�3)S��IE0�q���W��_<w�
U*�L���-��w?L��t��y��-R�h%C"\��m�c<ᵜ��7f�>����x����]���v�]u�u��ų�B�E��Ė�w�~�mt�W˥����`4�G��*��ދjށZl'���0A�ě�\S�r�-�3�Hg��`&�`)a��������-N�Q� 0؇�ST(�%n_CCv�� �UP�A��#���]Zg��'*�!��a�?i�U$��K"D�}����2��g~Q�+���&��J����L������杄�L>e�o����z]1���{�����9�l�po�v  Jx˗��$Q׷k��;H3���D~ ;bϪy�]��t�F�6��oBfI��%;պ�BH�M���\� �J���՜���;��^�����[i (S%	ne���߬�Ƅ5�����e��<Q)�F7�l�Ƣ��La:��oʩ�.���F����L,����!1��s�r�Nl=�*<8� ���j.��G�q3M�Y7G�������ldg�a�G��ی�>�3h�Ȉ�'⤰����K��c��m=N/�g������dzy/�pf��L?�:~��wr�����լ�R�L�䮌k�,�P�zK��!�Z��/k1u�IV��!�<��Q�R�4��3���`:�p'�FJK>3�\��FC�>\i����w7#����6�F۽�x
3��[e�C�Y�a��j�!�:\����j��\լU[oBʛ�U�@�Pj�������H�o尫��;��L��E �6Gɮ�F�)�KsW�!ev���4��݇���Fe��{Zuv��M���2梉�)��UI%���6ۙÅ?�Uy+����P����Y��0�$v}���ZF��<&�F�#&	!�1(b��IV�(�e���0��G���Ϣ�� y�&+n�N���p6J_�n�A$$������[N�IB���[!�j�54@��lɄ$�ƁB��P m�S�]"۳��;)�{�h<j�t���A������b<��,8��Jxq���cH5t�1˙
�xDD�������Y��Sr�����}A|b�����U��sv�<ӽ�#t�E��KU�7_��^l���c13~�@Z�V�2I��G`�L`V"��~Ǐ�Z���?t晸����_wO�d��;���6C�$����ڃcy��~��ZQ���2���M-''�ejˎh�h���s����r�����l��3��� ���
��w�b�d��H��O��<l�|�,��ջ+��O��N�,p�����р�uGb�6I ڍ����i�r�/�����[�0�!%�e���?<F�f; Cg�xU��Kdj�����*4�Γ�!�\P_~"�Q6���yr�p�|3�W)���7��4��y|�#20z�t�}��-��ۯcq���X�yL�*�&ddz�.��,e��l�8��H7}�"�n�o�%uN��\t�Wh�����4����`�r�9�4u��wz�kV?��s7��m��C���1O��A�Zq�m�J�	L3��󩓎y��a5΍���K��Bz ���_E9�I���$�$�%�yɦ5�4��}�kP�X�����t�����<ӸA!��Ԭ'�{fO��T��E�	��mc�(��)��X����Ruy�9��qYsD�"�0�N��	,-n<Jag ��(��C�p��k�H�\�	�AL$0F�^�d���}Y�$t�ES,lD��D�W��K��0C[r�xoY\\�p+F��q�Ȃ�n����<��a]�I��/�&`�k�di� 6�T|<פO�@u���k�U�a�;E&�,�)C�A��OO�XFf���������an�r�#�FwP����&(D�������%^H�ek1`������0#�z�l��1QD!%	���t���u>(�R������j��*� ��y�(�,S�0i�@d(4L&�כ��f������~,�u,��h �V!���ѺaR&�l����@O���}�a�t/��F技�Z
�n��h�.O�u���j!������CMdd5kܟ��������5��S�ˢE� 1 ?R&��M��g>ek�/�:2Ga�ǧ�C�Q�v�%�<9<uܡ)�߰��r��|�2ޑ��Ϣ(��:ޥo,���0����s~�C���j��[C9�c^�~��U]=�xƽ�Y6SX�1�%��G�)�pUg{~I7����T�u��T��ہ��%RaΞ��oz��Z��}?�W�PѦ,��nB3h5���K͏ ����5R�|��i*�?BQH�D'c�����o�aN��8��v�Ᵽ��7��W�C�H|[j�2-�9N�9�,��n�<�9N�1�:`{��ah�[�f�:oY�5F�F�Y*��蛓��=).�ө 1=�O[�`�b���en�j>��y�$�PՍߐ"�g�r �*�![�օ�����yVp�m�P��	j~�ֈu��5£��������E�۩JZ�5�qe��1z��j�%ǡq찡G�OS�]�`��I�4��Ш:�'�ҍ�[�'�Fu���>.�ҏRAISyhJU�Q�_Ug9�D���ER�BĈ��T��:=���3����&:�\ZC�6�m���vB���		�h�/�=���kw�c����r�B��Xj3ȗ�E^\a���<�����
xߦ�$w,��"�H�R��?s�x��n�C!� �r��T��DܸU]0)?yǐ���!����G�fJC�6qm�$| ��+8���_p�*w�}X�r�K�AD�����ٚ�@��`Q���:�6[���|`?��w�H<ce���I�L��i��H�m����M���R���M���Ң��N�P2ت�!`���>�X�']�fθ�*�A��x�&ibȬ�ZlS��!���� ���������s���2�lє��9�V�&�ε�7��Y���ލ� R�0��!_�u
� ����Ο�Ų:�u��X�����Z>B~k���l(�����O��sv�Iջ�NJ�?o����f8 ��p/�6��,5ƭG��'!8!h�X�P�	��������9Vtvdt��Fr�Q��s��/iA���@5)'�<%򓣸���R��g�xu����e�HW�@��BF�(xm,���"ەn��R���Е��O8Ch :
9��o��8�����2�Z�"�1�g��AR��w�1�Hx��q�A�^�lG��+B�oh�6���ܹܘ���EH���9�w���V`�/�
h�^�w�Z��<�����'����p��������M�����xCEu��"S7]ډ���x�o?��w`4��7��m��N�R4k������~�����^_B� j ��l,f�RFE���9��޸&i���4跨^�dX[�ȍ�*fnqU��;'4�ZK���MB#�a��1�b�l3���.��U�}���^}غ�DF�B�ˋ(��K�v8/D��+�+9I;�̅*�ν�:�n �v*Z=�|x��ox���>��p�B�p���w�)|��sQ�J��ZlKY����/^�V���d܃J��Ƒ��<���G��<��VFA!E�?��
ռI�vp����� ���SM�x8��q���@j��4�io\�XG�e�cOk�9��t��|<k�_;�+�a �n������}xoD�T�0�{^A}�A5y���;��v�?K�T�����a��b�<�'���I N��F�v�`�=
$tL|�N��K���i�����+���;�\��j�F��=��@������j51�Sg��m!	�z�Q��k?,Y�+��t8��YP�v��ὃo��u5�U>.Bl���p�d��~�0R����yOL��`%s�I�C+����P���v9��6��t��BWMG�1{<&�ǵ�p4��I�r��ޗ*��{D&��8�AG4��{`�B���\4gKV�K�����i�{�+r̳��5�臚<����[bOǒmT�Nf�썆p��x�wfg�G7:���
Ê��Rm1�	n#�(�,+��P���v�y[�:�K�C���J�y�K��n����Dc�+:6Ӌ��R�V�7�4�������43Iv&�$tqԒhBF��G�=�<W���XY�N�GaM&�8��M9ѐ����$w*fw�L�G��sLG|v�����)M%]}��85R*
�w�]ⵔ��x?�B�.T�M~���	ΝKy�oe��Gѳ�jia�M���71�d�_%lz�����#&�RE@��SX[�?�T���}��Dd�/��i�6�������xy�BR�`�b�_��.�H�,_"6t��Ю��:��	~�_{�,����׍C`� �L�p%������SI�l�,����[\&�۩��5������h�-��ɼ-�o.�k�&��1���gq[<�&�I_�a�k�9�3c%1c�>��``�7����4mL��B���a"����h�wD��ʸu{�B�m�p�%��{��IQ��ө|���]�H��Tr��gW�<�q�;�@{ya�eX���o/?}<8^�9� �Q��N�1Y��_�����2�LM2��%2"L�".ӡ�,���h���G8#1���,_�I���3����Y��Gd��qw��K�>���/�q�yw��Ϻ��q�^�9x�:��R`�[��S����If�u/�Q��M=���M���_r3k~$[&�F���M�A�܍ɯ��X ���f�<����������v��5�\#��.�Ҹ�3�{Y���U�t����o������Ҽ@�i��Gn�V����4:��"X'�]�t@��c%&k�a�>V��8��P�:��}<�@�B�K���y���k�tKs�j>�Q�e���iq[�OQE��bf�h�Z���^�,ⵦţ��"`H2��LKը�1�J���<��.�P�=��@���ˁ�"A���x�:z��\	}�w�� ��ɰ�:O��H6��q������X��Y��! >��S�e��jdߓ�\,[�:�����8g�($/��|Xn3�+��@�`�Àyp��./J��=�����O̠l� �};]j0s��#���1���+���������VsXg+��%.��n��C��3�U��'��@%�ul�̙� ��ch�˵�Y���Ď�� �ԑ�{���BNL`4:��o��#��OƔ�HH�@A+6~�ĄT1����1���#�^���|q�X�
��6���*��#�.�YzM�����EG�����0��H��5Heg�_�	e�#h�N�K�ZL*�5��<�z��䴊ۻ�Y�
�d��ͥ�������h�?��@��D�*�6Z�]#���2���?[��t[���r�i?�	A��S̶����_Iz���s�E@Lg���Q;n�g4���b=��t9�B$��K:��H�u�C#�9������=����,c�LϚ�?����IW�o�5��r��k֝�n�UZ����$8B����A!p�2.-#��"�`K�8kXj������(���#ckF�'�G�9��I@#�&�44wA�^�{ �����(,�Bd�zB*��V`���$����Io]=�S�����B��X)X˸`��� ��|G������ ����zvk����^����j�-˔�P�Gm+F�R}�J�$J��"���t����I�	d9��!�4º*
��n0T\���n��M����!]�~ �)��%^�r�Q� ٹ��6iUs�a�%�o��OJX�)����?x���fR�H����ח+��FḘK�� ��k|����b6�3@�)v��;��N9��s,Dk�?���z �����ZR[�4��(ـ_�Ђ����vH�(���LK�Ր��_a=*|���0��Z��#c~Q��㐸 %��'+��	����^i��n�TS�n�,�!�:VO�Q%���=h��
��<Fg�����m�|'[ �A���D;e�)��<�b��D��|��4^_�{P��T��E�	�rdx�G�s�xa�)�s�S�g�YAЏ������%���]�'lG���t�a�
�Z{�֊b�U��mA>�W�#�n�0�YVoi[%�%�|��|�S������p:$�	�v� �9!IA��k,I����ܸ,;33�J��}�  ç� ��al.��$v�豘HY�������fl��˦�%�M8�A�6��+�O��=gI����O}�T�l]S�	���[,f���C,g���ӽ�2+mC�����*U��í�>z����hi�z13�:�Z�h�t� ���Q*V��n��P ϩ��7Y�q"o���R�B<^[��0��v�~F4Ξ�f?���J�͉�Yi�~��u%�3�L���c�U^�'ow7z~[����2��z��j��[?��U��k���ĭ�r�'�$�(:�̛Vt1��>&sa���j~
�Ri��̎�U\��]��B�8�2��O�$���-%w���(7���zK�'_���{\�0#��h�Τ�1:w�dVU�J\�����:�|݊�e�-�(������Dk�,<�) *=US/�"��7�o{�>E�Ԟ��_\��j"D� t��-�'TOL�y��(������K����L�u����O<}�5,<�\�ϟ<~���+�J1�[b��C�wo�,�|Qg2<3�̟��<�{�_3�:uf��Ǥ*`8]U������Ɵ����S��z��-)G ��m_�8��m6l1�Ivk��g:N\Uj8���ڟ�}�X4ȕht]�WX���呬>3XW,Ԡ�6���S.q	z�r�ж�dH7!t��Y�ǡ~]B�!��(x���$`�Dq��v�JTv��>(��R=��=�2��-p���*�	%%��MU��K�3�d4>�y?�ř�V���k<5wil�0,�Nal�۰$������vh7u��N�j��a��HS4���{}��^9b�9�E����jHT��	�~�R=z�o��_-%���w�m�f"�r}ű*�`���vJO��v�v�'o���>4>���WZ�\���z�h��#��x�3��f�u��J��yF���n�N�H�`�1m��{"�>-�P�U[V����.U%,��4'dfg���2��I�g7�nj��:��5g?.�Iq���C����ً���?��USK7p�W6�A��Hd]v�jK�ig�I;����{�꓈k� ��$c���z�C���`֢����b;y���!����|��''牴����_�v��L�}��摞��#r��ne���D\����a�)�h�ً�8��hp�t�y�Z&G����k���ߒw��
����;A�*R	�\�0�R�}�UY໦!����֕`���Gj�~������vA�r�?a}�����=ŝ׶4FhO�.C}��)�c�P�0�B��/�Kc�s����}	v�RΦM�S���)v"pxK���g�Ӳ�rj3T[O�G%��I� 3<	<�S�[�zAl�Ȳ��q]�R�Sm�*S8�3��5�e�����VJ�n�9S�����v���J�<[���w�FZ;������3b'�P�j>J�3�S�F�,�K�KF9$L��p<huψ*چ~�.�N}/�h��c� ����D	��.�U�`w8���G�ϒFW��ϰKa]�S��
R,�����?��sw9�߳�O|�lU�XY��͙����<�>�P�c ���L�L]ďG����T�|�b�\O��/�&�|/��,�~$g)������߾��X�Da��4���d�eG�H>��}�1G�����ZaZ��Z|�O��ZF_��k���4��g_��=��������j�L�3%��vC5�ҿ���/�+�%m����:K-�#6���� S.P9�\��f�r���1�1{�����G�X=�!�4 ڴ�d����|�=��%%	����guӾ�l���$�W2����;/A9�Ð���|���Xhb��C?��h�o�1���6岴�0�OG�~�Ì�/����P�B��,�Q�����}�z��,y��Hrf=���F��\� {��-V�8��2E%�N/���7D�R��d߭�'��8ͺ�`5��,��]���K���z7s��@q��\v��y�S�.B�lݹ�������,	pb�琝��.��9Xzj��AA8����RT�H���p{��Bƞ��1���)Y YP5��B��I22yqՌ��+�꯽2���=F�V�q�(�;��Ʋ!L�A�`�es�aU�@oao�Y�]�E驔�h��2I4{�x�B^�$;�v�KF�E�g��@�)}7��'��vm��T<<{�Cy��H*^��=�)J��]'�U}�� ����xD����xDSS4���d'�%�2�{�5%�ؑ��/�ap�n�"L���=!b��٦:VJ�Ue�H�:t5����k#V��S�.�r��;�����!:�:���{!l�[�cꦨ'}K$u0}���D�Q�6^(�^J��>�b��=��h���rK�>�����DQ�ܑ�A&G�k%v�lq�O6g��h�.�Z\�T�Y�j8���r!��Y�P���O�P�:]I]������lXJV��g���q0Dl�Q���i�YF ���ۙ2ߝ�X��N��ڗ�sd���ǤD��A"O)����D�N ��NO.Z��)Q2;�������,�QC5���|c��g���|�l�$#Z�#�9��mzh���7yF�X��pU�9��=*�GV�R�$���8���1���؄���1��?ߔ	��|G����Ѕ[��%����/��-��u��L����1k��
��.�c��B�`��$0�G�r]�Lލ��
"^�F O��)$r:�]�^�-S�,R�iۼR}C	[�%������v��Bj3��/��	���(<Svt��A��w�K�nC���pV�=�nR�9Jo*��ڕ�;�qW\�a=�N�������ْ	�{��P�`��P�C��u	m9���G�x�|͗��m�غG�����s�,O��A�C��V�؀����)F��25pF���ٹlx]�ߝ��g�V���BY�	�hq��Hl�ĭ�����6�r}���r�yF౺Uq�OKhS���
eOHy�R����6g��m�Q����[Ū����J�*K�����%����h3��q8���*6�ﴏ+�Kv���4��T��ZѾ� �%����`��ȕ �◇ �/{�~�W���y�A�h�Iw���Bj��%�e䌛F��ɖ�-�ē��u�z�d�k<��)
�<��[̷�卉��"�j����z�+��#ȹ'md�+.���i�޲;͂�Y����u�0�"�&5pȣEy/W'���e����O�*�� ��|v2<9kRa"މԊE�=A�x��0�W�"W/t���r�׎3ՀA����v�΢6�	��w�2afZ�|��J���o���r��G�u�i6���A�t��X�=�Nx�ӷ��a��x8��V�S�DM�5�?e}J�.��Ew¡�g��E�_Vń|(f�������)��}^�����U����RB>�VN���?���jy��cWqGFFA�+�ʋ��7E/�؍@��*�C �.;E�/�`�b���۫���Y�E��J"�I��U��~=��Dx}k��V���� ��2��>��cN��X	f�L���S7�@�1*uf�R����Vg�"Er��T���R��7	�>��Ϳ�3���ʶ�a��Dn���Τ�a6n�Q3/��C��-v�2ol��;��;?D�u�{��g��r`WK�+��T|ӑ¸[��:h&e�Ȍ-�L��S�v�a�B��A�i��q�&�y�6c��v�P)�d�B��6�6��� abF%A��p���=���˘���5R<��eM���R\�G�ϿKU_�Ja#��b?3j�$�\�$�F	�1�ȍz "�V�ɆpՊ��f�<Si��ʉT�Y�F��|�[��3��+-F�_���њE���?�%>�L�AD4%̦�� �3�_��b'���������к�s~ցg7���0&�`������G\7ϡX��=��=��I��r���]_L-�	i?���hQ
(�S��a�	��ل�ֈl�UuE#O%#�s��L�GW�N�ޜl�܇�֋��d/��X��XeG.'3Z��ͯĭ��`2�A{���>�F�ǒ�d,W���<������>�^��U�@��dF�.￘k�[��t6��݈�W�9�Xg�X�TBӜ�)�Gw[��:���o�Z]�2��Ы:�-�"��H�����d6L����xk���W�6����X]X^ƍ9U�' �T.���oҨ���8M�5}I�W���$Z����[V�2^K�JrE@O�W��`dkZ��m��4�����R�簃�kΝ��pt�K8�3�C�r/�
3���ޕ��5;�qEpD,.񇽠�2��Μ�Ѣ~ꦺ$K�u������~����k�IΆL{�1ڼ��jo����\z�J&�����Qz;P��.Q%VN�r��K�1��ރ��!u6�5U�o[J�_D�� �J�ݕ< 40#�;�����.���7�E�
�f$��*��:~�6HXGr��_b���<U]�k��߭�d�^!^����BSmP�[�k��6F�/[+�L�|fQ?�0R���92�Z4��|�����Y{�C�/����AG|3�&_ܰ�맰 �����C��W��!�k*�5����a�_�EY�Wf��?�pZ��� ,���} ��6���]������Y�/�uǴ�Z���d��>�gx�C����!���F���#}8�[�^JP�a3[�K�3 JJ:��,<�L)5�@x����`�S�$�N�9!��i�h�$rӳy!��
��=���/l�e�kmo��a�˲_*":T��́b[��{�� m�̭\3|aR�eR�裘2��1�G�^�O����?N��B>�������'�JF��k�|f(	h�t��\7�y�o%�8�u�\�\G����1���ďp�����h.^� �&-��E�]�/_��ט�^WZ��YFх�0<2���l���&�|���a,���q*�Ӵ,Ds�>�g���Z����=�4R	l���=���Ko2�S�|���s�,dǙ��8�`�������R�gkxݨ�5 �?~J�l�;��1h�O�_�0ؼ�xK9���Pﯖ{~�Ev~g��4/�3<��	m��+�}	+C����u�����K���)�����C�J�*�Q{��A9%��4����iX��5U�rq+C������BjK{ө��RR���o�"���%��Ȩ�
�)̫�XLp3i��BY0�Y��*���|�I�pi?�N�"j?Y/�=��������j�㒛� � \�}��֝�o#�9���O�����pt=�|	�zeV�T�K�ƆI�B��:�@_xQZx�e��Y,�<��Ɗ�1�"E����z���D	7�[?�x_ɼ����^e�BM}��i�u@:A�VH���Qy�#Q�c�r麄�	Y�k��Y7��>�L��L�B� nH��|qP�jm�� %�5����M�=C��th$ǲ,Ż�C�U��k%⹁�����!u^�-���X��5-��zVa�?���sP��wS����v#��?Ϟ����B�IacԶo�tب�_0��7�v�Wm����|QD���b�i[XA�h��k��ap�8�)�؇%"�eYRp
�8h��PV4`�-OHz^ e'�'I��}u��#��E}]w̿�ȯ$�0s�R7l�^�@4�ԙW��1��ʯz�� ϫ���cj�YuI��TX�30,�rd)�@�O D`Aj���c3��ppT�j5��~���+���Q��#�"�{�۠�G�'�;�&�����������0���5ӈ{�^<4�GJ^Y���I����K��@?<�{�)���>/kyT߈K���0��R1a�	�h�A
/ѥ�=��7Q�v���|�O�QdҤ�Ks�|{��7�L��E�G����k��M��E��<x9�
k�.U�0z���u|���K��%W��M����Z
v���r��K�N�z(���h<�>�R�H��
Q	�9vwlF����N [8��=UC,��i�D�H��y�(��5������x�Ռ�S�����3ٸK��l8��tIB#�SV�#^��u�MF�^o�A) ������^<L�8�����P�k-�w�P����;2{	���MΊ�a��굤������r`���Vۙ����PuQy��mב.�m���d�*mc5xZ{�-$�M�!�Y�G��W�r$u�}�u�gxƪ��f����@5�4�yw!#�([f��Q_8�ӥ�:2gi��D�_Mi��h�XF@�i��_�e�)I8�s#i[�hϐ�f����%���{6��2�Yq�����"�}@*��z���,A7�a�a2��?���Ĵ�k�VL����O��'2���1�,������� ^����C�Lz�ы��$5��۞ 
�;V#3�!� zKQ�f#>V]�DUiycܓ$y6�~�[*P����P�D@��
����4��o!�	3d��(�;�t�%V�UR����)�����K,��k���1��qƻi�r�Z#�;,ϊ-�D�KW��@�����$Yy��ߡ�.�3R�&�-�]n���R��� n����S�k��΍�\�Q�!�lt�k4(��~8ŗ>�\����V{G��G8zt�9/�Y$�id���	���K���栀Ʉat9�;����b�/�P8|7�(�s�k�����Q���p"Ā������435�_"l��C��L�&C%Ik�s6n�&Y?�#���E��݋��Pߛ�k.�W���d�[� L��u�ʾޘ47��,�!'z̭-�����y�#�y�g�0�i/V�벪{Qsӆ|\�JO��P�,��nLa�&�z����w,�!��[�=>�k�(�G��fo�c��mk�,�&��8�ه[��� ;���DJz�RБ��'52<�s�}U��&:��b��Sw�΍�xy��6w4�c��^�0��U0E��y��f�e��X��:1>7�i���y��ZoG<��nkz
H���+u���]����+���Bm֊����Z�=�\�K9��x�]Z~K5|�盞9Il����
T��PV���Vl��Ȝ�N�����^&��+���=��|,(�����L�b]9�L+�%F����,
����4��4�����/��;�c��!p6�
�i�	߰C�h&�*��;[7��+���ڧdIL�j�=ۙ����T�
�밻�;�����zBtא
m�-}�c�ڭ��A�C���V�v��={E�T���2��6'����P\(����(��*p0XK0��1^���ND[���rq	ZP�����i��M���8�n�(PZ~uC�N]��(��+O\^N��
���}����Z��^n�r�Q�}		�`f��i��&�b�%��{hs�};`�'!���o�l�A7�G>UC��a���ZԄ�T�Ыc��Ɉ�h8q�������B���!E�PO:��9�g������X�C"�(^L����>�?���̲�g���GL�4-�QI�.��ـtx[(�����O?ZS�kd��u;�xS^)�C�wQ������|έd�(ņ�������?%{Y-�	�D���9Z��D=akʷ�vfYA�T�\���a��g�f��Q.��Y
&�?�b�c괎e_T	�j>*�> ��Y�4>��Kx�(�ca	0�o����X��F)��d�sש��^u)�����i��S%������dI+j�.�����?��~>k�߳X��
~����A���i�X�n�����7)!`�3}�Iĉ E�����F5�Z$GY�W+r�H`��6rb�?_�!k����X��j�!�'�H:J���t�B���hleҶ%�ϗ�T�16��q�����w[AF���l��z�����.�L���';� ��^��d�6���˟~�1bA�Hӯ%3 �Q�y��1f�@�y��Z�_�T��T�\:�����]���7"�pJ����A ����9(ox_�1Oo����%�	��Q�`�\��gw�gL�5�f��BZ6���F�	�����A�iV��d/�^�z����b��ȶ��ʾźK����~�{�n�����nb��;���\C0��I�I@.6rZ
H �R�N�_l����*�T�2@���U�B�ӤF/�om�Ds$Ab���h� @A[u��ݱ�oz����b�q�R�2yz]�R~m�V�U�߻
�z�.�1f�l��o��@�D�e/{�k55�B������d�`���i��=M~��ߏn�"|Z�H0�-��h6瀓�Y�*�* �|�4�Jo���cسg��жO���3���ʺ�*�'���Oq��H�K���\Z�D�I��>X�{���W-%�+���h�@, ~7���j�vT�5mIV>ye�s�60Q#��T��	���t�Hq'�A�]�>AA�n�0D0��O�(+��4��* uMZ])��C�:�?�����=��{#�" ��֡��u�����#g Z�sȏ�5�`�)0�X2�T.��V;��G�\��}��Z��_�p� "ܛ/��d�7��5Y���!��0l�������"�IE��8}I�5D,�t�f����� %n$K��U:b�t�.�gS��<�9 ���l����k��~�rj�WY��Q��l�.��������Kʋ4�4���B".U0�;oos
@z�T�u���/VV��	f�0���@�
��JBt������zޔ@�)�����tz[Aљ������P�4_������Ç�� @��E��u�
��$�����)��6���] �z�XJ{��:��G{1��k*��۳N��WX]]����M�$�`��+
�����C?:�z��j�M6d�g�7�a%��#f��C���)��8� �(�"�jm&ʧ�@�'�n}*h��؝x�v�%�t=� G�&4�~�Ac̹1���
��1�޿���&���]�[g�*�Y�dfXt�c&����0Z��<�E�ѽ|�����מ�A,aȠ"3���/3�Y�p]��mU�l�<4�τg��æR��V���CV�rq�k���s�sX���I;	�^�?��|g0E_��Ͼ6^ۅ7���}8��vj���l�m�0.�c�����u<^�P�`}.L.�/�,�Bpܪ$x��BA=IN�n���?^l�Z���N�ؒ�"п��ƣ��H��#܌���;�|��^�?}'�/��]�\Q��Yn	%߂���CO�)k��=So����ˈ������;}Abӂ�@�
,uN��խ�!�E%�1-�Tb�H�o�z0_YaA=�� Y�ÐQ��d�����G[r�T�/��m��I�P�Bi�$}���'��(y3��s@����SEH�S�$O�	�\6��s�D=��E�0g�=��<C��ʒ��皙��z�t?��q����x����]�4G�\�b�xru����?�e����gȠù�J�r�K��'u��|�M�y�})�r�F���2��A�^��������kyi�L��5d\է<B~x6�Q��^��g���!�մ��Պ��4�A���Vr<8��ї��h�X��\�K��<��,�gɔ�(��%����Y���GLP�L��E8�7����%`��>� F/T��E��+M���3�k�Tk�IK��r��a�����n���wiL�n���E�Sh�1)�(�(6��G�N�Ɠ9�u7t�wmD�kX�x�	���`􍘼�%@�*A�w�iV�8�c�D@z���	)em)ްkC����D��Q��0H5b-"M�g/��o��Oj:[��M���IjB�RlJ��)/���(�"�b�J��_��Χd�eQSO(,�%���l��)&#�T��c�@R���7�n��.+�IFX���p>7��}��d}�J)��j�wV���69���?�?,N�9�j�@�
L<$~�W�H��]����&A<�Z6Z�y���.}M�0���?�`�<����E�禬�'�.>DW}8`�{�D�{T%��ă!?���������ĉ�V���� {& ˒��U�6�{�F��PF܀�$�"�3Md<g��N�m��-�z��5��9l���b}I�.�z�����x��OG9s��L>X��1Ę�,n�� ��j������l�/-���Q}Y7m�Ď�/6�J�.�t��^��s*b̖vX��Yi�@�nK6Gx��]�"����E	ܼ�:��'N�,7!	�dz��`���It�j(�Ǹ�xa��B�Xf2�j\@���"=���8O�5���-U']ӑ���-���@�3�M]B-9��/�k!�x#����~K��<r�����`qg��� 3�`>x�KT/b�h�f�r]��,����:�m/0�ޥaX���}��@M��Zף�wO�6*��EEN�y/��^��B�8�H�?6S���N}֥IK�J�m�H��VC�~OӅ���%SP�"���KA�Eu���p�4��kw�7'M��#w/�g�0;+��\^0!�h+���3q��a�B�l��w^>v|&h���)E���@+,�+@���&k�̇!9l�7���ה9��L�C�(L;�$��;�*���7d���z��Et����+Dɟm��z�����cV�w�i�� �7H.�V��[���������#} e���so�
2րƧ���T�2j�;MgE�5��穭�²��g#�o��F� ��0s=r{TAϒ܅-�+�$�o
�~�酱{�}���n`mX�ѣ�����#�X]���j�wn���Pe�
��;'�HE�D�8C.�5�fF2�-kܯ�dA�X��k���%":�{u|N\xV�.�]� �f��pב"�G6F�}.0L�%1}����H�#�71�l��il(U}��o���'����)z�����FZ0�d�I�u+���lЇ�Hc^Ԃ��8BF��:���I���E T]'�m������=�͠2�����q=�32D�:õ[��u\���	�Ď��
��XlK��ܔ�d�'b��HӐ:�y[�8��n������:�p��`�7׌� }E�e'AyދG%��s��-�jBs�M��%o�xJi�y��E߲vS	@�&�R�G��C#�o��T|xh�>�)���&�]��ld�b(h&Z?ѰzB��]�z���֒]) �x�xGP��ag?�T_+�d������xձ�R1���։�1��7�5$�e��)ӺtYw5;�|IB9xy3:�{i�u�@F��b*��;Q[�|J�
_�":�,�R���R@JD���xYBP���Nd�7>6�e$�]�	�i\���/�4}8%j����PEj�֪cY~����]&ι8�WЧ-����{������ң�����V ���-r"�qC�z��2�o&Z*+��9~�E�C.����iv�c���㘟��dT������m}DKx�����D,�4��pl9���Ϲ7~s���hp8��Y5�����?�/��&,��ex�veB1�7�5Hui�n JT3��'3��`��5�h��mť�H;]���� �]@|Ә�l�����pJ��+6.���C�.�*�n%�B������T�׀5�GAq�<Ņ�KB2����#P]"��L>�^�Y$�=����ak�#'�r��jD���O/0)�s�j�PU�:���X��R�dc�� �;+D����n��G'��He8�q���c(��*d&���+�TJ�� k�UU���ZA�����զ
�2������P ,�v�d�m����F�[D��!��,I��QK�]�¡_n�haZ�v5N6��%h��*�j����Vg����kD�g�[�ҍ��	Cz����=}�+{W��4A���yלA����{��u��>y) "k��a�f](\�)@��:H�V�Sg����Wz���ҫ�1�A�.-��ދ]�r��dՐHm!��FZ(fp�>���KUG�"�ȅm��cġ�p��X�zu�����z��$^��f��-�ظ�ni��[�@9�}dR��e,��FE �����v��Ʊۗ�]�f��{cz&I�E�Ud(%w�;�սΤ���I�Ib�֨����te���iJ�^M#$t��A�z��Z� ��$���jB����lM�+� .\��j�"��Wh*�u*�]bK��/m�����C�*L����&�=.A��IiMl=���ͥ�Z���<�k�R�;�G�L�x�ѽ��e���NX75'7�����N'A~=�eҷ������0�7?�?#���x'��Bw-�[�ñ�;��`�V���\j�5��qz_�K�v�r^W]��,m;���t�$�L��E�f�V���"@���_$�r�s�˞.�3�B��d�]��u�e`��'����|�yD�W��ʝ^9g෼18�R|V.�\��A�:�*^�r�~�Y3����s.���*?��ǅ�{Qj=Z� �L귡Zy(#�D�|�y$]�b�{5s=�@���*��\�4��=ـ�|[7���� =9��(�W~���w��n�jv�໣�'�-��S� WO+��|���=G$��]�P�)��E���N�L<ͪ�P�E��Ě�����?x����܃mu�^E�P>O�O|@��{�V�	�dk�0�Z@�B�t �S�C�=��Ʋ�\S�<��b0��&��%���#� ����(l	�c�¦<������Nc�9�.Y0��a<�xH��08Z��;�q1�\_W6ڇN��p-}η�D���ff���=qr��OR��g���.c�o���m���TN��uj��U��7G�����N��*3��JԄJ$(��!*����Y�R��x�=!�"��c8���^enc!��̷�{��I��enro�[�a�*�����j�?h	��I4V�^Qi$�9^��%�;���	�}�%��x1k�Iau��j� t��T��x/��L�5+���|��!�4� ��2��.c4�!Q6�Jh�3��pu�9�]�!n&Y�H9�m��T��h�VsG�I����_ac�|O�J���EI?x~\�x|���v����0�b�6��x�W�2f��㚊u��+�D�oå�����"�ʈ_'its"���<+%���6�&�t%��7WL�ѩAp��Y�H�D�SJ�+�@�ρ[�@��mV�3u��fO���|�+oƧ7DN��S�����l�;q'g�a���S�r�-i-~�ЩG�ܔ2	m�@+(�M`����@�Vb�ך����T�0��w��Pzl��]��&�QL״2�����w��~��m� ���d��/J0��O�z#����c-�H�Gș)jvHf�+��M6��B���3�����_�c�K?��mJ0Y�Օ�������Z�^�&����p�V봱A�q�pH4 �F?�v��-�X\�%�oU[>OZ�d�X�z�Ont�q��S�VIiz��8����`��r�<�ڿ(u�*}���հa^s<�XF<� �כ�V��P�U/�o0 {Ƹw~a?��!�7�����]��R�����Į�3�1B��E�S���a�KоA.�/��5G�!����&.v�[aݩ��L�7�z	��Ҝ���D���#����*��-���͔ӮZ\�
�08`�rV>���S��걳�ldx��B���:W'R{���3$M�ER>�P5^-����٬��>���m͙L�M�<�5������*���6��0�`�N�1��.�(�Q2Z��bDiwk�K���I(��V=8�f�|�����l�7�9�X.4Ɠ~��Q˥b�vݨ�������� Ε�¤Wa]6���|�\��tƦ��:�k������%����F/O�#���D�[�\D!9���\C_c�;�-].C�ԩ9v˂͐��a��Nǐu�X*cr���3$N�Dk�so����r�ߋK)�f]f�O�ϡԧLʕL��� �B]�k(U	ne�
#Y�)���ۮ�[C � Yp�v�����]����U/3�	�\�e#�&��D�KW���N��$q��-�\����G5�嵤P(NY������2=���A�2����V�+�����; -��]�+W��8FPL���Lx�ݛ�A����C��^�%ﮪeݨ�f�6�.���6���%�6��;SҨq8*K��!�	`+|<Ͷ�t�l�Ê;�z4fƨꭢ��B���/�]f��mű =nvdt��<c��u�/x-��S�/���������r���@	��L�_���!���Zܼ6"�����&��|��~2��IO��0`Z����rs��:�C<��3P>0�~r5b�+U�F]�ۯ8 �ɯ�u��
���2�G@�=��F�VX��d�f Fx��!�{w������ 
�H�o��@���c���L���G����jƒ�.�3�M�Y�pk�/-�ى N���j�b�OR�1U��_hy"����+� �� ]�["JL�d#���x�(�'l[6	:���7H<���tG��'e�K�0oXp�(ȹM�GI[��MD�;I=T�t��B�	�/I#��������6 $w>RXeR�����Щ7(��B�:���"ؗ��cߤ9�d���1�m���\�Wn�-�G�sj���O�_��I��Av^������Xa��'���*���t}���2ڹMK"� <�-�x˿*���!��_��<�$�w2��g��F����S7��>���z8Ɲ�����_p��P$XSx�5�a��3Ã]�kOF	�  �@U;Ja
e@�����N�4@�.>��6`�`7jaK�Ϙd��l�5�ȐP���u�J�m��lcȪ�p�^�k�	u�̾��d8jZg�#�Yf�#t��:�J�<[���L/P񋱶64W_��V5�)d�=��%'���mLO��\�w:�X�"�
_�Tj�����u]��ߧ��e��]�� ��7�!G�����"�a���
���A"��Ԥ�X��N"F*i�v�w9O�jxK�a��(�9�ɺ�E�v�gP�V�8�F�[DJVo���k,Z�r�x�z�;�J�JY8���5��?��[���L��N❛�v�7#����
��_�+�O��$����ۓq��Ś���0���鈍jy��̓>���>6@����ҕ�G�f�lpO�C�f�������NǑa�kP<���A�N��^k�sz5�$�r��ܳ���.]rJ+V,��"�I3������v�����"n�.r���!H�9�w����$�tx�c����ڀ�k���]�Vy�)fyk��K��%#r�iR��0�E	/t?��e5��j~����1&bdw��p�w�Juk1q��{4X�֣P�)Z8��iUiJ��%�� m-��;��}�kr��:lD{L#����b5/IHtqS�`ag*��*�����yO��9@V�ۈᡖj�'��^��f腗�%1�<�m�
��G�F�ZG1ړ��B-b��X�/m
θ5�h5^T4��Kd��$<FC�t@jZ,�Jd�m/ۑ#A-Ҍ���2ߢ:��L >gb,6����#ۚڦ�y
�?F/���X8F�b,18R��)�0�Y>u�pԫ��'��#3����e��o%��7�|l�AGF�^��;���R	q���T��̅X`R�~��Z|�1���=������7��O�
�!D��yHO�Y��b ��!f�qU�j��mj��nS�V�ꁗQ��F�lH�������;�N�r�d��T�2�ϋ��rZR������1|-���č�$-D���sZ�$���]�zu]��շ-��"=�:y����*='�p%q��_<���:��U����eI����y'���.�"����1��� ��x���t��,�!�|�O�Y��u:�hM�6��E�	xx��8߶��q���Z�B�j�'�� 줱��b�aR��^��$���Fl\��f��Un`�;oԟ�_���n�I�	|�1�q��d�9����r"�y�/�ۻ*Ӱ���wqY)ƌpl��Z.�|�&��VFu�ܻi�h�ļ�-SQc ª�m�x}0"�p����>}+N��0��\4���ig|!�[��8� K��Ø����5lpY}I �@u���:��=t���,+�j���R��>3�K�,�)�k4%��!���{;OcgE�|��cd�,׏c[|�x�Bx�M�(��p��>A g��^���?&�ދ�Z���hZ̥�Lߒm���P i�#}�Ad�H)�
�=�A��:/jh�D�Ysi_p! nW�jCF~����ۘ��9Sh����K^�Ӥe�P�{ז�5r Qy�b ?e�[�A�����60����j�y�p�hU��dΌS_e�Ц�.�em$�����(����9�LO�6G�+w���!4�F�~ �d5����C�I�k�����l�|�\�w��R�� =�%��o�?	'F�m1�H�,����J[�1�i0�B�ͬ{*�A�:Pr�����ẶR/�O:i]�DM���b���ph��m�ċ�Vw"�kS:�qF�fn*��gP��n�S(��h�DK��><������J�:�>������,�B�@ �u�z:ŗ��6rúg�������8�6��3������8�9Nx*_^��Y�bo����eU�d�g����^e�'p�̢3t����슮>y_�

�3oT��|i��ş��}B�l���}�
�Ԥ��@Y?U�-v��9����;���$�g xj�ז��K���^Ӓ����wC�@��:�_|�����Hh"Cɟ��t��7�&8���pL�Ӟ3�������b3�FxQܬ�N_����\�������Ǝn�`���M^�a���Yn��K�#u�^��uo�f�W���y�	�a�ݟFR'���0��_j��`���k�fŘÍVǛQ�0^�[�e��r�}Ѡ��4����]Ϋ�&����g�}�x�z���l��y3pY������	+
P"~������"�(�0ɹ��@��P�������d��D�7���^�{qZ,�V�'��B4�k��.itX�ŷ6+�絿��S{����_�M��{�n9[La�-�_�\>�C�>av��ǓG�<������ݢY	ݔ�%čL�#^i��t`*?��3`��E�a�iz��gɱ��ߎ`y��o�[X(�k�����B��(X�y��Y����em]�Zul]���WyĨ��챣�/��n��{N���R(�7շ?�Bb�����i�=�w֘�R�kXɛ���� =[l����G�����8g�'yP0���PK��Z�q1���(�F^��3�j׌q���Vj��ݗ���-ʞ�$�3�SS[$�g�j�Di#�Q:���l��wM�5Qa�ȟ�e����l�~�%�6��J�4�܀��|�N���i3^ 9q���/s�`|��&!v9�/_���
�[2}hZ�k�cY�6�BIp75�7�Ճ(V�p�DG(�3˲�������eYZ.]��d�O!�����)�Y
��A i��l�z��u�ްnXՔ�Hy�
&w'\�@P�͵'���bK����J�ƀ��P�g�u���4v�\Q�Zi��-2	.�D�r=��q����d�i:����8�eq"�lC�O�)��D�fC�T�0zF��_E��"M?�J"��o@��g-C���O �:S�m�׸�`jk��|��}� ��<�I��^`.5�V$�����G��N���bD�
�MN��dP^t0�϶���9"R|Q脵�^]#�@��q=����@^����q�iE�P	o��@��m�y�߇�\��&��"�YT��F�Ϯ��LC��R#�CtA���������z��1�O�3�G��5~�8 �,�2B+T�J;�ݍ��O��L��5���i%	6�wq�(�zʂD�ȵzv�9�m��To�<Q�{Ha��ol�{xH1N4�}��m��n��K��:����X�tIޚ���N���*�3^����_oz��3Bb�O�9P�Rd�qf*�6J���r׾t�)
��s�9�?{�MT���URd.ĉ��T��)�LU�<4֢̳#~sTD�7��0����5t���5Х��^���ք��YS_>�$�����:h�;c���%�Ť@c�4}7ij��8�*�m�����l ��n'X:�CKo^��fW���}���
�l �Y^�T���1��?#Z;Һ��~kd♡gy��R� s�d�7�٣�(��IZs�&�YrsF���hO{$ba��{TDJ�M 8^�R�ȗ6O^¦��I0�
���GK�:^�\1[�.ŁiPM}��ux�L�5��c�@�}�]����C����x,�T8嘩h�o ��ݛӇ�9y��UM,�<L,m=�fv�~0��i]j��L9��E �-H s���ٓ��ӑ@�{H��<�7[�lQ�]1J���ɴ^B�|��:yA����a��$TxTJq�vg�"(2y"�]uv1����AOL��̖��依��l��{��Gx����!�e�������_t�_p�+v�C7��,'ӟ�=p1�r����!VC#�olsG��	�o2��s��c4Y�A�����je�E*�]��#�Ƥ{�Vف�T>�jJ'WLx�}���ͷkr�Ճ䭊.�8�\<WU_
{�\=Q+���I��K�q���ɥ]ݩȐ�Pt��ﻋ#�򙻨�BށDiIw�����H ��+XV3+��vt��P%gTa�_�;C���.#Du=�4�W������Kg�Ɍ˄Z`��a۲�Ke�8�0x�iۨ[Bw�IxX���w�tS���{��&N�싊q�73@��]ਤNi���ا�C\@c\�/D�Ѝ(��p���m��;�����|_��V1��Ŵ�IBZ�T$�j�o�;���Lf�w��U���.���+Ұ�y�S��QT2N�xLoM�WM� �;�bq��=����F��J?�=�?4�6~`�󺋑n�l���K(˱8Ŀ9�~ju�X��e�(�	X��0x�]�iMe�򖫙L�p����Ә�8s�g;���tu#ٍh��}mI�^���ԯ�)��m���:�.;&u	���]%�ٔ�'�'�yv�=��f���"�ZZ���Jb\��G�fTmg!Yn9���F��p�?��d8u$)="���x�2IL�.�3A��/���'Q�[M!o�*9@-�$SH����8?@���">�T`�x�y+�U��b�{���d�7AA�
<�
x(����\�E�ׅ�X��{17k��ZP|�6��f"�h��$z����K�a��i+�|S.��5�#���!󐆔4wF��Y{��ȯU���7m�SM���-��o��I�����"�?ޙ
$�Z�Qqu�t�7P�ݠ���,�\���w���hd�G�S��#��"�����Хɇ�7_�C�ۇ	&Q�/h�U�� �7v�O1G׬#p&/���� ���ђI�9$���J0�Z���r�"�h��і���@�1�BD;�L~2p�~�1���ښ7�����'t�~J��X{������V�w�Q�Iɿ�g�� l��Τo����3|4����ׯ���e�`�r�PF�2��whl&��{t(w[�SMb��5:o�%_��PڤHA��~n��]�î�8A<Y����`nĲ̖���$<ܩ�s�ށ�TW>\���k��jU{ʾ���(�=��M�,K|�� �p-��J��C�E��9�H`Qhi�P0�g�$�@F�a�0(� ��I^��x����F*�*˲�ܪ�Q��ߡ���\���˃�E\E���!��4*�64KR�U��wx�T
	^�3�SH��a0�@
���+7�#��qg�SX�Ep*�/zS�*�l�g�DRR��=*�_I]{p6߀W��zr,�X����H���IL��D�� U(�l�)Q�}����!l����)�6V���	��M�)o��n*�r�&����A=p��d������E�, ���)�w�>�b�F�l]�)V���Sġ��F�� ��^�T3�D����T�K�;0_��-.�a�,��u�"p��]z���"U�/��'c�F�*SA&]Z� IrQj�L��;4�mys�s9nh=P:��Κh�@��������z�h?b��-<�kX}&�QU�=���}M����W߈�z��Y���A� �Z/.lЄ�C�}l@U�������1��0@z=j��Z��/!��I~^�)<+ٵ�C9�(��̪IA?s*_�}�Ȧ�|�|p�"���Z�k%�mQb�쵚�V�h.9^�Ynu�}�^����s��jd�?� ���m�୥D/#V�peV��*D�κ��w�tk����t��<�oa�u@���{z7�B	��p'e���o�|��{�4�ج��%�����W&��{D�`����^:�uA��VwK�J�����3O������uO�F*�9��_E]m���R�v�'�����t��Ɓ�t{:�!p�'6(�o��_0���mًc���bQ�S[(�1�Q���7co,^VՇ��m��B8P7БNb��6���n�2#�>k����+�����Uo��F�4P^)%�=����3ƃ2(��=��u=���%d��Y�L*>��7����L�H5)��?��&W!,$Ь�� N�O�Ǵ@f�� �+ �Vrg�A�|,�f�m�z��8�d_o��@��lC�̢'=5._r</�S�l��X�z�L��M�����!Q����U4&-�X�s02�(��+��nR�.�H�Z{����>�<@���x��"k�M4T�]�Ω��w���H�k�]�NR�'�5=)��^�;G;��`�̝	�, �x;L�u�IR��H���@W\�n�]�11Y*���v��X�q�9Z�ҍ�@[0��gkb�)�������v��k���z](g�')[��3�1��@ˇ�Ȗ��盶7��Ώ�P�0�'7�̈́�Z�C���Bm����LCI���F���دG�|ި�L�Rw#���4C����=����\A�BCK�7�N$� �]�}�@����� �v48�\Uۨ;(��A��^'�>�JH�w�c���Vl܊�BC��V�H=�82 �B�	���V�´�c.y��rs���S�WM fE(Έ�@es�ҭK�o:�#^�.Mz�~c���ƥ�����eY�k���j'�f+f������G�ť��!�P����m?q�������O�E oz�A\F���#7[�6�|a�����F�f�"��A�S�l!x�c8gsk�I�5
h_��_R̴5��M`���� ��w�lm ��R(˔�	ѐހ�K��Z@%��Z��Ӌ�#�L�'f�qZ�v��G����$�w���caB���ǉ�g���k t���m`�te���Y}nT�9A���b@
p��i��?KX?�ϲXe���|��Cf_�e�E���O�>d�ǽ�R�	�G'o�kJ�pDx	�e�L�6�C��sx�Hm�sSj![�.���X���
�1�����3�>.0��`_X��P�C�q�:�vHF�ni�c%� [���
�^��t��-����E�8����ip��0���{1ˀ �ʆ�<0�r���39x8/���ئGt���S���3j{�Ƣ�_�B8�g�jư�)��AY���"�a�ل ,�?!}�6IK�M��o��������f�GO��磱l�:�\dc.�D8��O8&��K.Aӫ�����⡪��/2!�y@�������5�Z��<�[tK8߭�G.Y�㹆#N�l��u&3�v�22�N��z��t�"�0yS��YDtÚ�G$%h�I���6�%�ROL�vI�w�v\7qÕd����h+�4H�%���ά���_9O�OF��I��	ń��+{]oޡ��N��1�5��I�.=e�(t�tst� ��}s���ڸ�"�y��HF`	�k��h��v�����BF?4�(Xm�ଉ��Bv���>���K�d@p!z�	��ų�;�wKnK#��2�ٲ�[F X{&�n�ث|#[Lb)�iu�����r�U�$=k�YI���{��Y��xl��,�i��$QAT5b屚&�4,~�G�e��D�[�����Q=��{m�.z]%boYX�9J!+f'�@6��J2��V�l����!q���+6'��I�J�+ϊ�G��o�������	~��D3�'=>d��u��|�����:X�3"߫��FMG��ԃ��fN�r���I -;9�fֺ�q��~��$�p�ӌ�Q2�	��vi�W��a)!�O�M�/����Ԭ�O'�����\ԬcҶ-w��Is��~z8�p�� �H�.(ͼ��M9���)������s�0:'�*U���ڷ6�ZD���b����&�0��6�s��l�Q�A�Np3�Ĉ[��������XT��?�!��FV$Fv4�[�:��k�+�|i��mL��]Lc�����z����h�7u�ߐ��1���(�0�rX�z5H]~vׂ=��Pma���a�j�F�3�����*)<���C��ҹXz��<�����#���WH����������]�5����$�QÏ�rG<�(���A�[���7�����0���a���&�������L��_�2)Y"�:�k�K*���o�������e���G���Ӻi�D7�U���J|��j���A�58W��ґ|�����k��z��}S�m�i�8���������|T�N��<�˼�<���\��0+(���O~�GsS�f(��2�	��:z����2�PdB/D�FD̿�ih�x~���?g�R�qi�5 DUN~���CE��P6$@��s���Oj{�&�7�\MYw��_��w�	���$DY�dȶ��LP�M�_;ձ��~L�4��*~z��B�Q�!���aC	5��hY�i�<-�3��_49&$�B�Sd�#`�{���E�T��%t�N�?Gq�K�Xe�o���y`t�g��4O6�{{*�yjQC�R�4���D������V=�U��Q32��*�}����"��J�i�x�6|�'ﵞ[�Hp�_!g�
��k�^w���_���rj6���<g&ݲڡ���`+)���d���t*��&���[h�A��s�xvc��iO\\�KoWM��h�m�|ep�LjC�a|$�C�z����6I���ͺ@|��Uyw��m�
/,��<��M'��^LBo���f��OtH�T)3T�xF�r;���8a�@^��>j��c����.@ɩ1��O<�m,���(��q;T=�66���]Xti�����wo�w:�֣Dc�%� �������v�ׅoʦ9ܦ�/��!w��X0uRs�G΢�w��4��U����ޔ`�$�"���]��Q���4�k���L,�U� .�<k�:��I"��) �q���a��I�������M}��D���`Ξi5�������A0"���7�U�5pg�}d�jf��oHO{����Q�Qs z &�x�|��0x��?�w8d����J21D� )��^$V�z~s�?����J�Q1�ިc�ջ����Xl�Q�#�����3:��/fx���"t���cC4�Z?̨ �^��#ˤ�,���B:���.+�s�zR%^�����',�D��ԭ%�A�Xb�g�X����d�)��r/0ɷs �Ձ�9�"n)۴\X�&������
�R���*x��=)��O1��GfG�������8��(H�ç�4)�� �*�J}��ڹEIh�)�� mq�ե�T)�O`�c�F��s\16�Qi��}��)W��a�C%��C]��X�f�,H)7H�i��{}z}����r�	�@����ソS���-�����5-2��p�Q�W�B�u)����ӦT�#�'h�Ӯw��u7z��6?~9/�~;<Aq��ݔ-ܞ!�/�.�P�[[��L|"�ԅK0lT�IAA{���H��tg<RB�o�j���y��k�x� eTDW�X�g�K�!]|���w>�QDq�
�����
�=X�S���>�#(�n�>"����!%��W������K��M��U���C���g�D^�N�t��L��;/p����'�̼�����ϧ-n�<qk�eL�9�̞��Z��R$���bޑl�5gi�Q(ٵ1�NZQ?��;Q�-&d˳������* -���t�ʀe������E�h��b(E���Y%��<�%�?yc �.E�O�:"��PI�A�{�iM��v>[(��+������H$��j��aĸ��OH;ǽv����W^�K`~�������}���/�����u�ɟD��L�FHV��ǍK>bxp3੶ØNF�����@IM9F��x����=�\���<|��~?,	��o�r��t��}�Zb_�ʬu���G<�q��oٛ�;t�����Mf��3a+J,Y��>�"zL�.ġU�*}��B���P�����v �3|��� �Q�J���F,��(< �g���{�"6P.��t�|�VW��dD�b���;d���́����Ki��DF�������L�j	ׄ=P�ۦ����0����G��:���Yn�Tu}�t��o״Ts �X�ޖ"����x�e�� *@�G2����'��z��-��ЬO���	:]>~���M`���Cp�����j���s�������r!.�"�|OR ����]BʁA�AV���{R���@�E
�1Ǘ��W�c���;h��t�����W��)�]��#���e�G['�O\|��S���$/T9��p��0�A|�HBĈ��;o�<Y�eòo��8�T��Z�'QIKH�"��}�u�/��S��[�,˲�ϗvQ+�&5�Vn5!������m���-��sܪ�N��
�� �C�@G�`ai���!,s�C��C;��wj8�&W������t����8��F�@?'F�) �%Z�#��� �A���e
*�S�^�<�v����Y��!|":ֳ�&<&ĳ�W�L����Z���L9�di%�%���<��6S�jS0�s���p�|=�E#�?��?c;o���Qҽ�ىq�� XzQ�j=�r�E\K���X�x�&	���*|����Z��_Z[�l8�g,�E�Ч7��C�(Jd�z�@��.AA
잀]�L�#w��{.qJWB�8l�� �_誺!&ih�S��V3��I����;_�@y�(��0(Bqi�˗���>ti�/,��)��P�6�z�W�i=)�@�v��!�aH���3�vs�d�(i������!ѳ�b�c���3և��G�q�q��f��}N�ʉ��3X�ڋ�Ze�����P��{��hN��ysR4��o�y���أ�\��|�W/>pޯ��L�SJ'�^�D�1r�'��T�,�#�j��]!����,)��^��g0�@�����h�t�H�BW4%@_���IbLv���u�q�����L�4B���즙X���O��ڱ�j�#ְ��b�C枰���R��{�;�nCe�7�s�LaZ��$�Ih�䏀�|�t�v/^�@�[�9�r������w�T�1�Oe��.�r%&b[y��ۏ���j7,��n�ں	j�H���!f�p&Y$��4xƟ�#��ğ~��Hf;�P����ƀ��18�N���/���'�ظi�١�Qb(��^BN�T�����{S���J�`$��,�ndw�}�v��_����b�J�Zl�l�W��?є2�~�@]OS�`hN�)sg��Π�O
hm �5t����2��c}^�W0�	oٍ�@:�����\� �I����(�%���;;�'V�z;vc~Tr����������Dv�X�ե��k��N,�H(�<��F�c

MkK���D0;��1�J2�{�r�da��
��B���g:o��dR������F	�9>�Rׇ�
�]��M�>3$���b3Y�������+��&��(���͵ *T�I֩����>{�2�xB���ޣ�Η��@�"��o�3�ZXqD���^�O�m<2���?t��� E�z��q4��68�+3XlT��� ���W
і�.ka�z�)_���^{$:������Z������E݉�D(��|�9�B%�p<�^)y���;>\=]e5b��3����������G���G��U0�Y�@d"�h�ˉ��" [��QJ��ܕm|����s�c �!;�Xk;n�~������	R���%"k.�-�h/��c�V�N�u#���ڢ[�xD��oc�1<��f?0řO�<�����x��Q����m0E�#�q�#hI#�L#��X�G[������h'S�{t���V`*����\�t� 
mT��"�N��3��kZc�AO �)v���R�X�D��?���v���7�X,77)tvpd56uIn�.���Q�4��e�M��=��Y-� x
"��<�1,8b�"!w,?����c�?�#T&J�k����Jח�R���fB���xi�,8�v��gOL�ϯ�eߕP���$n�� gQ ̅0HPXn�#������Z�XY-��y�#�f~^)�j�n��@/���~�GFP���-�s��f9��v,7ȽyC2IBk��lA�Dr>�<'�w������c�>[�����b�Ӱ�aBr�_I%�=��(hӾ�.�Y�LFY3�3q��"��``���;��B{@�w`/L�F�W}Iص�[::M׫�!�?�N�(,�!0&�ދ�ܨ؈s�uբ���DJ?3b����c9�=7�ޏ&�V^�OL�)7.Nt� �twת'z�x!�ݖ�U+�"���#	����Z��(��r��YQ��(�T���28tV�ڇl ���(�}��u�vh*$i.9"�n`(�0}�T|�sɎ�M�g��*�۬��M�	n	��j��ݝ�T����9�U�j�@`×��UZʥ[2܃�E#�"��*5�fq�Y"ż�]�W%��wcF�W�W:�"Up���f�lcCn�Zn��NR�m�7����i.�ɱl�����'|�<������eLKa��fe�6Hf����d]P)?��.��'  E��T��l�W�\����0�(	�1�q� �
�Uo�~'��Wm�Q�&�6.��{�Qj ߟK�R�ފc���5��+e[�2��"��)���8���T~
L]�튊4�G�o��΋�����6�Tu^t������Nay�;��o�#�A�u5�EY��LS�	�`�եj�t@p�f�N�Ε�|�}X������/�.�yP���4��Z�eI@����`@"#�!3䏭����8Qq4J���_Җ��;sun?}@�*�x�M�B����(�iO���4U9yD{��Z��#JSIΡ�
9�B/�@�F+��4���f��V���U�A1~%�M�s��r���]C��R6f��Y#�٦��=�ԗ���n6�����୴�#m��v�j�~�f����R{4�W�,z�".�o�A��G�pMǇ�.G#K� ���K�>�A�8d��ο�Q����ku�w��)T�F'��2g���!	D�@k8K�i�\�E�=���U(?�~�~j;�g���� �SS�v�W��d�]A�pO��5w�4�������;���Q�P߾�9��7�WR��� FnЫ�۵$,�Y���e�V쓵�
XFb����8�S[�ds���#5!����:������xD���S���_��|�ي1��|�� ���[�do7��,�.�׫�̺R��hm��P�3�1�����>Tt��9�>�:�;\��q��hm;v�N�+�P׀��MA0��K�T؏!4���!S ��˟����������gw�c5���H8��ME���T�������5��G�@�Y��b�`����5w#8B�[ׄ���G��%��ջ?'~�5RE)�[*�Zc��k�z��+;x����g���ᾂ��`}B,xUȳ�o�'��J ��[�s��y�o�{������HS�۝��hX4^��%��[Dj\�S4l��͍調�d.l��� �T��e�i@A!B����e��C�����\*x�����>��AK#�[�l�[�Hg�)]�pC��5��E�W��q��E���l�]���"w~�ʔ��n]�d���x�W��Sz��&`�ț��0�A�����1����v��@J�#6�>��&6��9�٨J����3 ����F��f��F��Z���!d�c��ب\K0��ڂX(�d�liU�87c����9��08��.���_ړ0G��:�0��},����s/��Ľw�`�"��'���!a�k��sB̂�C�|�?Ü�&7���)�Fwk@��8^��"�P�;©�
��`F:��V�UJ�P��Ƿa�NS�X�3^�	�'���+Z/3-����6���R��-��ԍ|<r��˵�P��ր�r�Y1a���s�W��m�XA��q��[Q����Aa�����bķ Ռ�S�n~��C��r8����r��
mĕ����i���zQ���������$���H}�MzM�y���?n��`Vp4�ke *�p��DU}�������&8�_e|#Yh�LQ���e��h6�N���#E>:�?@v޸C��� i����Y�7����+��êwka����,l�~U=��;;�g"o�}���K�u�1h/<a�dBX�)F^r�<���K�+}�M����цJ����P���m�EnA���i��}����x��31�h���iۛ;=����&���j!�)�Ka�Rz���Bd་�-F���S��K�e�L��HX᧙�MdfJ�|{��Q�"Υ{~ؤ:�J�����g1i/S���U���d�1�]|�o�
�<ʞH0���ԝt$d���z��Tʧ#�����bb�e��Oރ���d���F!��oX�<�G�CM���a���L7��ろ�4�,��I�����D��f�4.祩��_���\�^�6���B�+#t>X��T@92�[2�*�c��	%$�e¬���XF��
�ћ�4'��;�Z���4P�Q�����J �rҹ�G�Y֩�+*�k�0�@k���:��pt�-�s��4�<ӿ>-E<S(e{�}����8��b�Z���fǩ�<q�1L��Y�ʲ���u�o|��)`��!o��\B�T��F�a���ARv�$
��t~�u f�;��D������!��x�9Y�����IZA�Y~�+������E:rg���|>��cGm|�鸙Of8�P{�Ё��ٓ�͞����� U˴,�/18<����:8�)�$o��I�F����n���s��. �k�x��wL�9�|@��@pđ$�@Ԝ6�1����=�W��6�0u�z{{Ġu!�d<q��r�M�K<��lT�t��:�I�Ԃl4^�}Wc� Fh`Cp�ȳ���\�m�h�{u�DQ港ql�іf���f�d��C�v�Ķ-�ڧ�5���kS�{�NR�U����Y���@�^͹��+c��"pxO��̣Vk.�S��K*J�R 3���{�YB��q�*L��X��)�'��c���Ӭ$mqD��X��4ᳯU��s�WQ��+�P���Axnj��,�N|�Us�)L�]w��-d:5��8��!k��J-�DT|���oP�G]T���ǝq�����g"֬{g/#�}�}��O\��9��c��I@�E�~ةdJg%�4��P��o��Ȯ1�ׂ[�0�_��x��.B �_��e��h�������^ړzߤW��n���7k���
A��w��g|,�����7>u���������X�D����ݙ� a��.�]G�����>�ee@[��z��`��!�d��Ʈ��\]��������-��T���cA^�����B��g:Qx���v~(*����&ݎ{-�o�2-Xjz��䞔w6���y�b%?�����%'��d�BJ��?P����)�ۤ ���ja�m8N��7(�����@�#�2��J}Yń����f+W�28��R�Ν��`5�o���Tܒ��~c@�ɷ�+�gN���~_�ॣ��p�G	��.%>;�r�,�=~��"��1�	�?H�-yl��f�'�O��J�)
��heB2}fYvJm	VTLm�֌9F�g� �ݳ�f�2�#�Y�)���CaO�E>.-S ��+�ˆ�
^U�M�aX�Y8��4���PP&�B2[f�6)m�&��1����]M�TM����jXH�N�C��2���u<C-�J(:��~?�ե��9�@q&�dPvs?����mP�	�|q��T�O�*X����l���b�G�$1�0��v.\����LG��;��Ǐ��8�Au8p"A��ngI��)�D8���e�f[&�.i����`��]���_����|� rLY6�v�\[�����]���a����U2F��������)��(�������7B؀1(��G-�T��é���$�7$����h*Lp�q��n�����;��@�Q�7O�S�� �Z�t؜@ �7T� ܦ��)P奯+"��Q~�ki~�S4['�I^�V�^�g�.@ٜ8��;�Y{GG����Vy;�9��^4
�����,��~�0���g���=+��,l��w���:��;�`t.3��3Ue���@�-��p|b[��I�\&�ÏU�3��3Y���>I���e2�C)�-��-3��\m� ���P@�2TF�X��cT������Bd/�I'ON��[��Ϲ�)F##c��d�ߑ�ƃ�æ�EQ�����7O���n2D��u��^�A?A��T�>�'�㮾?�t���\�JRe. �������`����Yq
�2D�!��U�i�7� ��
dp�~U���'��?aoLD��s�q��kRO
���^�V�*9�ZVg 62�g�k�^M�ٔ{M� �+aJ��K�d.jb�x��G1��L��[1�FϽ�
K��3��d����Tc3��kЋ�_w�\e��p"C��� �>�,D,Y*�K�Q.��I1z~%?~���^��-�B�ϥ*Ol�f�g�C#.�e91��枠�W�ׁO<�ԕT=���PB���	O�.(���a3HG	��A����m3�����ekyoH�g{ņ����NI}��.Whg��$I���#Q�z ���Q���	���5�t!���;�}3��j��bM^-����B����8�c�j�.���[.o��	^��%)X1�a��W�(U�zڏ[�0�|��Z����%9-#�)����}r�&��0�ȉ1�Iߎ��� J������=�KC����_��͊�$; c�È\�� a�oC������wœ�3�A.�9x�+DF����p��:��z)O���h���$f5=ۇA���q^�������vtgp�X�����u��6�#�ᗥ�Oݞu�!���κpHiE�h~�Q�&K7���%`,o��	�8�w��,8鷀�q<՘숡��xa�** X��#��D�p�]i��V�JI��r�t@��МdW�.F�j��[<&m�pn!Obb��}P�����X�Q�_�W!�DS8db[d�	G��#I�F�bQ�$sG��mNї�S�*�Zt����AZ}L*�,��&��Da�'xj�V�H�AJdV}�ٽ�Y�k��ݿ�/��?���Eurf���<�� v(&K�����PW�L�IN%��b���m����wj�BJVY��y"��ʥ�/�r�`���l��6��>�f�Ҟ����%��9'�n����8mQ���C���Ȣd]\
��X�/�'8��T�鈦40�&;U/\�P.L//U��~pid��{Y�A�e68�2]+z��xr��������ڮݓn�#���|��c/��(��MW
�W&,�;u�0
�̃�%��!=������f��s����y�̡"�g�쫼H� �3�����GL1��"�N�I��h�\�E�U�\�D�qK� L)dh��0�շ��,�2�s����:�/�;�O;�]��#7�K�ʴ�2���5jr�e��.�
�f�JB����Ѓ̸�.�b}I��5Zb����'F)X����l�������R�=iǹ��G*M<��%�6P�Qhf�ߤ�`�R#Se���w`z����Ɓ���D�����2|u���̣%>�����P�0o$1)�iC�.���@� �qS:{�n���Q^�%m6��W�ؓ�n)-B��K�	��1{�A2�������3��L�k����Z>ê33�c`�߄lR�f���j|w��
���C�Ƿ�@�Lo����x��b<�����C�)QN�j9J��^4s:;lv)eh���N�JKl�a��u�s�t'�=�F��H����`����\�UC}��]�!��	�){�=pل1��PFO��O�'	�9ʊ��iVY�k23c��W�NU����FN��g�R���8�<�'R���N2%�~�{ܤ�nF �˪I�+�Ff����#�OS8��Qt��p���q����qz�}��V�+��-��qJ��B�fb�(\��:-�{��.�F�j��.`�B哖��7ۂ�2��ź�����'��!���ވ�+�Z0z��"mS�֦�_,���$2%���W�	f-8rh�a�2��j#W[Ae@�'
�|F׷�{c�x���&�MZ�tI�t>���W�~��~^�xY����PR��	���p.�,E�\ǝ��0S�Em�9W6i *��Z\
��!�O�H�޺6n��\�eH8���ʩ�6N�$s��h��P}mn��Ø$H�+�e�8j&j�A+�e��Y O ��9�P���'D �����,����x-�G6��[��C}�F��'�|� ��_0!�>s#��F�;���V7M2���=�̰�h�EA{�c�B���:�ɍ��qsǋ�Ph-�&�p��F�����9��~���]ԕ����禽���i��mh�gy�	�)�氐��	vH����A!����Sb����!��!,��1l�L�#��_��xa7P�?T�;#�_�괡����`�Ѻb�[hfЏ��[@<�����ˑz�F��'}�Lk�,?M�V��O�Y	?6|b=O��	���챼�<��-Pi6���xi;��ή�tb=��>��,.��v*E�2��>�̮�0�ۗ�{��<����z�LD�j-���O�\.�a���q|�4�����0�[��+���]�ӡ˶s<������ �.�Fi?�PZ�b�ȑ�.Ƚ�_V����HS�/� .b{\I��c{9_:u�<%W��ޘvL���/�$�%6J�Ut�!g܏*a���й����
5��6/�jV�[d���0���I#�нV�SF�9�{$�!Z��ɢ,�g��¥�����J�]��~H�}�����Aߜ��������-�Yؽ�8к0�J��L
�CfN1���Ǣ �Q�o�8!̧��}�@�$C��=� T�^¹:X�Y�zn^�L�������2x/��Yņ��1�60C��Q�����+1�A_�H�Jb"8��[�C(�A��]�%�;���{����5[-r��{&��|�|-� �Z '�1-,�=��w��",'c5�:��}��[ɑ��?/tk��U%(|����j��������GI�Y�*D%�j0��iј�V煍��
��4����&�<�\2��t�>�ρ.��X(���$%�o���X���;�R�x�K� �!����kQl�̿]�S�H�6	+J���sinV:v���f���F�'g�� ���}����H��S�A����O-���bi�!�����d匕ޢ|�oO��=�TL<�Ⱦ;!��c����e����+R��{z��5q:���q�!�k�(����	ň�$��P�[a�q�C����@�!�`���$�LhiMc������d2�2'U���14~�h��}��L�ʡ_[ѢQ�㩓^�e���Ц��"�>�m�Ca���3$��K`���O,�'�몲���+���c_���y��y���YIr�R�柪¡���DWF`����uwOpL3n7R�b�Wݝ��r����м��I�s~�-��.k���Z�fn�zSr���!��y��Rp#\æ�*QX!�<94�d>��(���4e��Ӱ�Uw�̳~�k|4+������{D�)�2��/Ϫ��7C������q��U����|�>��ɨS"�ǵB�spMbF��>��^8JR���"��Ts�[u����-�X��ڐ�9�s��``s�4�$��=��`(?p�4]����	���<�������!}�*#n��)4Ѡ�f���A�C^m>��A����~���j�b�76ô�p >p�]MeQu"���	��2��B�x�$�f4�B��Fs�%\���������P���J��&�`���
�mB1׌�nN��-z�]�0PXh~H5iw���X���/?��� 'Q`�W�o\�8���WPX�jCųU�A\��M�4���Yl>9@r:2<��v�t�$��#�JH��Px$����f��\E�-�ũ����:�'	դ�v�Y�s��,����`-!����.��1� mK���N�S8IS*�����z4��e�0�!�bo���jޕ��X%�R!��̥^�?K�0���<�k�c�a3�1%Z��nnR5��!Z�6�?���暑�՟(����(��sԫf�#󩦄��jA�oA;uT��ٰ��a��q��a�(���,!���C�֟���8Z��{b,tʥ<Q���v��rO�Q��3�&ϧ3��B�|DJ�E��s)7De>Eb�<.6E�g�GT�����se�m퓚B�)j�j���)��2�I�̙�]��y�m���;V��1�@���O�	�<���?��(7��޲n؟l\���gvEuI_��`�M�0��iџt������U/�)��ZO/sO2&��-Y���.�2ٽﱝ^�8�F|`\�Ԓ/H4���Rm���0���C}ֺ��- $��!;²So��B����!VOgM�,Dp��B�o�6D!Fw���_�1�גۮP � ��=����bM�Z���گz�(|�@!�����JMd��`�ٖ7�?���^���78W9�j)!w�
l���I�Rm��$?�S+{q��YV����9�hw#x��|���HP�N�/��&���V��׵��JD��;��5�ǖDb���d��`O���A�R)b��SX�[�
�r�l�EW����������U����	9�b�ʛv����\K=�,ԾO��������k������ R�^U{|/�H�j� ��t4n��-���3;h�������*t��#](}Ϭ����pI�x.DJ)b�ϔu�%J�(��πegL�;�ث�֠���"�!m�AR�-������i!�x��\�q�� M Ѹmu�Y����<�ժN�V+�'-�m�8L�n|�kfk��蝛FD�2�����X���hꥆՒR-�ɷ�mm�Y6���Du���Y}E��J�_nN[�~e���{�h�.�ЈK�-���Z���+��f�J�8����V]�_j�V21�]�	�N��	Z?>�kF ��������{�|�X��J�;�c=/vVq���$a�"���,G}7N��'j�hL��ȥt�QT0[J���)\�x|f��c�����*���ߛ���nZ5�l��P��a��
���F��r�������y1�~���] ��x���Ǭj�Y<�b�w���O�	��-=9�(z����)� ��m�}t�n�4�vl�u���5������W
7MYP3�!Z`��&���=Z����l����������'X�����-���X�K�sbo%��8&D��{���:��w�7F�Gm��	��wk��7q�	Z��3�(C��x��W�gz!����{�x�Ӎ$vv�:��A v(g�EN	3Í���fF�Aĉ�ҫ���8::L��ZNw����o؇g
��b�����f����
r7�O�]t�f7l�5��ǝD�E}����p��L���E���~�'���2��M;-t ���U�����	;��g��nu�iMŝ��P9������-�̿/D=9@M>���4�t�@P���X���Xm��T�wG۷Ko�t='�;\9��#	����_;E��ev�:�b�)���$Pn��f�����هe�xAX�{v8di�~�x'"C�6�6�S�
W�B+�k���#;���|��xP���"�5w�ַ6�3m_���Dn�Y��$^ĨC"����ӦC��?�Y�����K�A�݃�q!��f1oU��,�/�Dײ��g��2��6b<��hw�R�*�HT��������C	>�XjR2<��%�oAG����������a����c�꙽��/��5
���掹��H_�ъ������ȷ�"���3��CY�L���_@��B*��Ճ�h��L�k#ͩ���*D^���
�O�k��{s�(���_��MWv>X�ډ� x�
���w���
0�����}_P8�����x��Y��(zT�����z�9;�e�2����Yi���]���`�5j�q&HԬ����p��;k�4
.� �$3�7�T����,���TV��F�6ӻ��x�4>�hӦ�k���ͣM^Ыth-%�!�Q�^��h�*S�w���$���t������pG��\� �!�v����w�(���ۮ�q}ly֑�|&nđE!
hq��)ɰ�`U"t��k�I��yڄ���Ra���x��"W���D&�+� �ݼc)��-��g�<�0d�m��x�m���ô
�P-�Ht��	$�$�p˧��%�z+?]O�&$�wd/�;���1#P��������w�L_!�U`�)�b����>�� ̖���3��L��r}��5�K��9�ѼhQ��6�b-|�x���c���I�ޑ�D���5����ͤ��	Wן1t0�f�9�rz��q�	��	�_"X3�g�8�x/;�|]�@�xʑ*� X ^v�@�����'n`�g�A� |V�]�F�FuO��)��t��j�Ȇ��+lʪƏ@=��z�ӹ��65��ޓ��\�u���Gq՗�tƻ���j�]y[������ձK��dpw��ضn+�߄\x�Έt[�6{�o�+�ɂ@�y�X~��+	1��I���l"�o���%ן��Ф�րHd��4Ю���n�{E�29,5�CS��;��K?hs��yń��.Dl!�{��g.y��.&��e�B5�`O��{��!�_�>�iX�ݬ��R(�)J�T��	;�Iĸ��w�C�qV��qd�ݛK�6�:�Q����U���b!HD��aX�݁N�$?���1ׂ�q>�,��u�G�1��R�2��Q���g���b����e�Ol�����
�jz�*��p�L�ZX�O�Uv�I��q%G�CM]�aώ�\`��,�!�r����!x���핮Zp&ќ9��hS��d�쎁�wV����GHZAkxA�=��!�s�R&�l��4���5$Of>��� �t�r	o-(X2�dv��*ەq�{���N�n[�K�u`-!x}و�
��ǂ�T�e�Z^�/����*�$���/R�(����N,���L��e�f�m���Z�t��Ƹ�%ba}��P�h�C�����W�����3jKL )_��?�-������[x�M��/ojBg�z�!���P�%!G�V� *�J�Gp�Ri�/,�������U*V�Gr��s؁�#��f���T���6�S�ܞ`�N�����!�k�&�(���O@����dХ0�s���MP}n�`@ڠ�� $8������>T�eF��R������Lb&vr�ձ?�Ft6�3DST����+����N����ś@A#J,�tF��<WF����H��N�z��;�#�ha����i�âZ���(l�$Ԣ�Vfi:r[��o��|��!ʓ�+��� �O��5N�;��IGk�A����Q'h����f�+��{�QwW��px���l�ܕ���'nH?�̳G��a<�����W�~o��WD��T`�"����F��_���A�*D��$�0�g�F�T=��x��F�Xwg�q���h@�4�1p�dn�Q֭e���{��	�A�(X/���(O���U�[4�h���0��b�:7�4p>U����).��(��Rj��.Ej*i����������&\�jࡃs�#�����^>�j4j>�K��%E����k6ZY��_pA%����̍T��ARe���g`�mm'�%X^�����uLM�~v��V�-�\]�_m��"���N�voI��*T��d淋�{������_�M@���1����M�}�����O��a��s���_k�]Z^jU6�Fo�I#���!��T�b"����'�����ȈJ����R�'Z�w���$�d�|֏��g3�>��K�i]��6���lxJ/~�CFBy�Dj�K���\L���/���$4M�Ӎ���q��4�S�f4:����7��-�紑�B����
~\Q��xˁA�G9���Z���Y��l��� ����g�!"��gP��Ouo�@1�Ҁ$ �bP)��������<��ۍ�j�X�}�<�����~�<��|�!��ޯ�[r\[��ݒ�˦M�~�;.527�`8��_G.P����;L���c���1�<����tA�H��=3�n<k�3�x�k���W'\:�A�P��k�3���!V�������|�⋆q�K��6��,��q}(��(΄��!��b�uV���o30)�X���+��]�D�gg�!-i�
��e�ix��[[/i���ry�Ȝr��eC_)C��)�0�r�,�ne�S�Q)�n�I�����m��_��r�-�O��W�J�!o:
.؎�{Z�s�C��^��to?�Z��wJC�M�^E�fPb
�;n�7:�* �>�a*0�8L���tڲQĂt�����f~��)���,~����sDU���I<��W����n�^�!I��;䞢�̵s�G�Q��
=U(q�q��E3#��5�*{��Huͬ�p*cz���JT��҉�=q�)-�*�Ը�	��^.����p&��}���Z)zd�����{ׯl��B���
���?/�Kc�6�K]��! �3��GH"�3<meథ�E���Z���)������{�p01^]Le8/]�d�Z?�8s���	����b1a)���1
X��e�*H�e2���T[\G�Y�t�����2��)���&І1�_��t ��!/j(����#X*t�������ە���X�Uݞy_���\إ駦����!�9��6�����.���<����g�|����b���"�f�C��z��8읐��yr�,���ᑓ4]�t��Z�qٕ�jP �yΥ�Q�n�'@J�E !L��q��\������P��`u��/�������4��R�����(�:�E?��'��Y�T��%��ߗp��tKKkĎ���V�B�t��j�D�����4{�؁1	u�1]��ᝦ㸃t+���v��V3n�!
�=�6E��W:ڂ^o�xƣӕM F��s`/�K�]��B�q�Z3�>���LRuE*�*��S��P���#��0JE6,j`��W�k�;Gj��r���w ^_U��+��븁N᢬<��6��7��)oC���@s͔Hb5Z���K��W��N6L�۷ej�G������_����J �>���Ԉ�-�2r����U���t6���+6'4�fv��
���w4�����|��DC��#�~���]ʐ�S��W��dT�Ւ�f�*���Cn��kӻ64)+L����7<݈��eE���{fU�Ee-��7m�M�(�����^�{.���j[.��o���7��'3��mk�z���.$7��pB��ߊ����c(�J}d����d�: ,�Ǻ��J�OD�����6���0ߘ���(Y˕�^�5�v/7�Di�'���c�I�;$�-�'ho�\a� �Ta#�f�U�����ϲ���oS�tMIs5����)�;��oX��#��1��mee3���� � &�n���mB�@�Ťd>t�P��-ČCf�qj��'Ѝc�cs0�ϗ���dv���״yf�ec�[���e#ϼ���ppV�m$i�0�ҏ����B����F|��y�Ͽ�LYr7b�.Ɣ�_�xM���4f���I����� �+�e���z֕�R����M�G)Iu�  �X�9�=�<(d�{�$�AA�O �wk��Ni)�k��b�MU������zۼ^�U@Jwy�龴k��:XA.9�t3��a��(4�dz^X!2ii��T�M�����; _x�ώG��-��c!=��A"p���x�q:���A�J�|��7���kF��2Q�e�7nQ�B�%@^�T]���w��s?O�����!j񹌠�"���S4�Z���*Fy�I(�˿!�Y8�\[ջ�(���Sq�E0�H�$������*\s���k|L�l�B����Q�ƓF��A���'~�����t�[!@�?�!�H�����.�(uJ�|~���4t#d~�;�ˍ(�2����2�o��A��s�'�{�lƧo+�������/������'���S�l�a���S����*<��B�(si�����ʾV��n!v�1�ї|Ho��$	�ܪ�Ǡ�(��w<-2y���q��\���CQl�m��'�G%,"���ᒗo�W7�f�-Ĺ��VhX��_��Ҵ���6�P�R���*���L�!o����}65#�d+�χQ�����,]��bfϺ.֬�������+��c�>gWѦa1�d�W�Ñ֣�f����ߒ
7�Opqߢ��(��1�$in�2Qaw|Ő��yܚ�Y�X��
֟�}�����z�ɵ;��Z>���h��oKU��Y�9�l8����I>���=�#@��᣺�;�]$��oxX�)�"�p׼,!p(uj��ȔV��a�0��
�W�������*���"f��p��h(w��3�6��^s��{L;Y(1v���*����5��$��}Tg.9�^�|�"�C]'I�P�䩟�+�Č�9�Jw���+AB��Ɉ@��(7�{�JV���H�'�r�����)x?'ۙ��D��vYj(�h���SF�ho��4�#�L<$��@T���4��ɳ��[���d)���+}Tn��"��l�
���,8�����Jܙ�֤7�^�h7�c�m�� �u���'sk+'��Q�i�V<��M]��ڣ�`|܄g��֧�)9{�UT��`F8�d�i�ÈE�s�_,�&!��5�C=�Z�֊6�VB�zY���4@��D��a���Ӓ���{S����o���{Mc�᣺4� ���@��/�0����l��1���"��*��P9+,&9���[�y�\�'���O}�G�EZUk��UB]�,�ݖ~b_�i�]�#V��>}5�E'0�~���� ����h2Ya��0�1�����궔J]��@D^����`����;x�8�F��;��m{���F2Uڮ������y��;m��
ժ7d���2�L�+Z�A����d��si�47G9�Ko���H��%�S�t�[���P�C�KS�__�w^o'�["^3�VF$�6����h�����A���o	Z�A
�.m�T���wj��>L]��ݹ����_���Q��ˣ;Ŗ�`5N�qԭ�4��E)&�����x�?��k^.�Ò�%n)ւ����Sln���C�슓�a��=}��xSˁ�ٮ�lr���3\��x� ���19��}ӋӽV ڧb��;�2+�W��V@�]�Fg��Ay����Y�#�u���5�����q���#�0u"�/9�&�qЄi��OSq�trKl'c�\��N_ɏXR����oZi����V��մ�a}i�u��n�Ns�����
�ܶ�\E�;�իc]�d�O�x��ǤY)*�<�Jߔ��|���)My�ǆ�Y�����w/�>�d�.�3��Ǜk5��M����N�P滱�`�}�>aA[c	���^��#ta���r��؎&����M0C]\���0�'2�Ei惗'�a��Г/�t��QN����]_@��R�I#K���l2�݄F-���cI�*v���K�g16/��dڰiX�&����A�4�ի�^�g���Z�|vS��Ey������;�zi��.����В�-�Afb��������y����S�O���)7�%� ��E�GF~�"PO��@�N3�U�t�9��j�L~T��՛3�,����~���nV�gޒ@�6��Ц�Y8�������<�)��f8��cC7}憨�C+:N#&�Vd��$l�3o���v����͠-���`ۛ9�pn�ǳ���E��"p�r�&;E�u�FTٕ��w�C�^V�[a���9���φG�'��P���Ұg-@Dfj��qnO�����(;��d�;UT�|zoݓ���*,���iS�d�3�]���}�`�$+?��X0��UQ�^V/�9�b�4/�@��^�}��ƀ����lhEbBG��\{����C���'��EN��޻|�.��e^tj:�^�	o�@'�����IqǊN&�7���_�?��O-��L"9�;;��=R|���a@k'����W����N��z��q�g(�䕤뀢.��fC��sRUZ�zV���a���A�w����%ZhďU�@��6x��~���@ң:�����a!��	+{�����q��Bi n+t�7���/+��VjC����^��|�7�_r��W�8O�.��\�j�r��٢�%�l '_�n����gF�/]���)�$)��4C�aې�Sy�lZ�Q=2�ڍ��P�P�_���j�V���+�3V���mU(�Y��>���"��`z�_�@�`� �,�l@�}D˕ě�>��iY���Um��T��<�F��ZW���<�]Qݳ�m�p�BHx_��|8�ç�7D|l��t:��l8�)���S����u1Ǯ���ٜ�iK�m�*Ws�Z�@������H�kKZ%����<���PZ��³�ԩتo��J�*�:(�|�������E���Ǯ��u-!����.�c���G�{�CRKH=�Z�z�R�~���N�:��G�%�[�/w����9Ne�
�WW%Z�	�f�~�}�"|���,��D𵏰��9e��z��>Nz�8���6D.?]����m�P��SL<w��.��=[%��]b07���Q=���>1�j�%A��;�|��.�S���2��1�>��7K٘y;K����/�i�`P�O�^�Va�?"�eT���p7�[�%G9������%�����*�ݫuv#��b�l��A��q�S
�����Bs��S~4��l i���"�N�� �SL;T3g9�BN���-����9�懠�3���@�e@{G������!&�B�(�&���!ź�ݳ���t��\)0������Ϙr�ͮY�����-5!���b��P��3`��VP�J7��H���U�:j?���E�<A�ۀ��у2ݪ.�v��٤1eU<�Ě���^L�.T�aG�wh�֭���)g�n��3�蜍����i�!�����*]{C����0(X�_�{����wm��;)�����rʷv6h��Ce��׸�u�����Fl�X\ U.ّqRk.G�c^�C��&�J�A�[?.2��I!��՝ܛ�ђ%���x�$kt		�g��\S��va�za�w�q䓹��q�9ܹ^F�\��HB|e/"tsI�b'�P��r�с6��w��iےm�eQ�vVz2
��B�|�7�+m��vz�s���y�q�I��aѿ<���G���*tLq���%[45�U;�*\r2�$2���W���?w�,�;���Y��f�n\G��*���\+>q����j����a��Kl�T�E|�8<��hg����h����-y%��T[��F��s@8�a(zq����opr���U�2hfܢ;	*��G�pD/��j��Ѕ��l)b��"�����!$��_M[�3�r�\R`"�_:�s1A(П�g�>�"�#f�ɷ*�&��F|
��]�]����nv��YB",h6�7Ρޅ�{~]��ɹ$~�c���x?v��D�1g��)��h`sN�\{g+ɴ_ "�qM�.r�Y��66.a53AMq���mu,Zը=۟�$�K�9a�Q:u�F��+�#�$�k��@y��Δ�o!T&�c���x[�>�๏�������ٔ7H���{��VX���x����UiBW�Z�u�Oqhv8�/�K֜1���hH��x[݁�ߎ����)[���`�����{�4�fC��2a��5����~-��Y�l{�>p������xc�̯)��3�����)�X�?���/���?q�EQ��4F.�4��8d�mŰ�g��3���rE?��V�u�L^�dO�o�#s�B���!h�ؗ�����Ⱦd����9NG��|�P�eu��@�&�98���1+Բ�E�KTH;��' ���_o5*^��`Lw�a(��|��S7Sx�t����xr����X�`5���xQ�=�r�t���Z}R��� VI������ɱp����el�*~����R�@�K�B)�e"A<.��+�����3B��A{�ꠎȸ�XJA�9&=��DB����m�߲�f����'԰#��	��n}e�Ȳ��3�1
&���)��yK�CWj�C���Vd:c��&��)^�K�(?�E-��GR1��8��Q���˧ܣSBù
'^3�I8ϣ^���U+�_�?��f��_����v�9G��Ҷ��{�y�hb�5�a`C��1̒�*�U9���$�1�ۣ��!�(�wR�Ό�����d����"-Gu����T�w���}����tlvz�?���(�B���F���	vڡ�!���q�^yJ�\�����=q��o�%{�qݱ��������`�����G��"�[M1�$b��3����,��w���Θ+8�����~�������U�|���ls�~g���/y"q�+1ck��`xy^]�=�VDt�	#�������@C-y�ѿYx�P2��P�!{4Ph�\�D����@���O�P~_ZT��'��9�wr�0FlV�Y�=�i��!j��٦7���@`F/��
��9��})[@6l��� ��Mŀ+�@����v}����O���o�k��v&��{%]gW}l��WMp�yW6~�i=v_{Y	M��(h�RE�xY?��bPIN6񋅂��Cg���ta�C �,�Ucmq�@>�\_��cX�;�3�!����ʝ?���<�V�a~=�g�fx�S��fn��6�Y���0�}.l�=ߪϔl�t~�;_2��a")'�R	����G���A�;����̦�b���9[�b�<�|�7z�(�K�ǂ^�F�4��lY�+�.T�To�i��ht�N6����b��c�0��n̯O�
��P�N�^b�����V���'�e�x*�U�#aA�&H	������{U9������D�������Z.5��5� ?�_�z���T<	�Ea&H~�E]z�p�!J�5G�����s�Izʿq��,=d�#+�T�I�ߵ�/����	K&/�[��"E8���	���i�ȼ��7�,��v ����b�c�M��2�������UKct�q4n
$2�v�+�)k電l��
��7����#[�_0�
�;L�L���y	���o�r댇c����T=�&F���ҐN�)�A7�>���k� l�� ��N����ae7;2CY�����gƗX7���?��"�-ȖA�xa��c����f^�Ѯz�'?[���5�ӱQu�wjH�X��u%���XƺFPSQ�/���wb�c�֑���y	_�`�W��E��F���[Rո W��/��Bg�*�TC7�L�[a���[�M@tk?􋆝3�=����
xx�dv[�޳�	_e3�Kנ����R�ⲛ�b���jJL�4WH�(���v�_&z�LQ��������s �ff�:�Z!mښ?X�68��q��Ay�2�e��O���M<�le�˴!�����|�[��ƿ��r"��+�$�=g�����/Y�U��"_���x}f��Ǻ{�?������=.�ޥV;q���hC�t�`�	Q����{�>$���5�����]�9��ֹ6TiU��lzfY��3�i�����'�\��E��� t�&�z��P{l���F?�	5�!������U!��rJ~x"LL~���8Y��Gg���&}����9�K.0N��TށM�R꟣mw�$	�v �U��܏D�#I;�Q8�͖�T�ȥYB�]��Q��c+h��jǏ\�,�J�)c��L�D/�@)�� ̂	p���b6�F݆Y��E��1
n�ʡ��ća��k�l�X�3�]:4K^<(�H��VH����_�ؕ�s��T�*��Qr��g����C��WX�����ܢuwSݟF H�{��Y)]��.�鮵����E�j���.K��4B�]P}�b�U�B��>aεl��i�mPB܊:w5��^>j$�9;�����&N����G*��7�os��)]G���"��b����}�S,$�[H��+��8o��N��rJ�5ƟE͡�KM{Bu��3)B$=��	3��
7}ߓwv�*�?�%ҟ6(G�S��b�f�϶6W_��9t/M|Ya�M�7�����ݥG��:H����t�n�r�W��aM2��e�l2�������Q�Ws}نa!��Zd�zW��¯�X�K��YIt  �7���Gk���|]CP��HoA*p6T]J�@��x���^$a{s2�h�aaw:7��E�9��ޕ�k�J[������U��ת�L4�����͒D����Ɂm�����n�?�*l"��E��Ll!D#�*��
��=�[y�?f��iS�i�1͇�p�����3����Y/����ǩ9��`��iej2~�X��l�i���;�v��7Fx<#��UU�jD�����I��L�~�$_l��-�{8opO�X��ϽH[����h@�m�����X�?ٖR^���E����N��� �3�=h���n����8��'�s�ۤdO֧S)q�U.#5�G���R�F��ɩ�P�'�6�� �<�Y�y 'jhA�$��/�|�M�'��H�$��] �X۹ɺ�^��
����?"������T|2&�d�˾��Q-
��K�����N�1�����w4bLBa��o���_��#U���~���$�N���[i���X:(`*�g`8��>�(p>���.MZٹ���]��u,���E�`|`NwB�+ �a�K2���ƤW�N�s��͆�<t��?�U�`v�Kd*���.��V�m������|	E��Fg�'��Sͦ�Җ-�X�R�_��aN�rҠ�%H�����G8*��+%�6��+B���:/x	����C��G�Jv)��	���q�m�k��� 񅫓�?��u�]V: ��c>ͽQ�/�;���_'�q�(��Zj� LR��S�{+(��q�F�g�����%�g����'����<�|Z�>�x@�=�o� �h�2�$��J�7)�P���cWH���t.�Ñ��>XN��]P��9gu��>ػ��CX�6)s�)�=��xj�|�0��U���O�;%&g9)��w����%����C40G���8?,��pVI�!�kMzm�Ts��{t8 ��!��ZU�h~��[�K�.�"�����X�3������2��_ʋ�E�|���3�U�^d�¦�T�C����%�R2nUƇ���dL ZL�ϩH�Ȥڄ�v��]�Z���B�w�;ߎ����$�3�D�[iDf�T�3���2P��@��m��(k5FZU�ʀ%9�zB���[e�db�t��/�����)�_�-f?\;.�,)lG;���H�w1Խ�8�	D��X�@�եϻ��P��	2�!0+a�0�\�ƻ#*4>i�۹�6���c
�߱ndభY\��G�����!T�����'pwB���%�&վG#��@�T ���b+}�ç����%��O+fj���#�R��q�Ϋ5��Û6�|���lG
y.8�x��$#'�K��}�/��q�\���i:V�dyHº�œ�rM�YQ�;=y����&�U�^|���ù)���t������fG-K }��'�@��.<���G󒹶$�@�'ض�gd���6.���Ym���Ǐ�LP�h��-f��4F,]���4�?�׭������C��E�	P��.�@Xꍅ��}̿
�F,��1D������>�X2O5�=ҡlտ.2�C��@Dg����N�A����+�BC�U�K�9���g���q4����[@\�L�x��f�!>ez�R ^} Nd� ������=�[��2��/l���45n�F�[JNx0���FA���u� ��8�ݱ�ڒ��\4�X�SްcF���$��/�_+#졯#�z�/o�0��"��/��
W�ϐr��!���X�����ǹ�P*ŞCnP��cLX�,J���>�Xl�7���%�~�K�����y���6�l�`F�hlm���̮ʹ�l� k�`�(y�	N��1y�7��1P�j��~DkYv��t��E�GT{�2𿋮� ��ɳ���Va܀���\���?�F�ֹ����ǲ����*� ���2m�Ҹ<�L�F�	���3-�ݔJ���!'��l���ݽ���hAʜ��{,>l۝o�r=�`��O�%���T�����X�Rҵ�k���ѭg�� T���K��@ 6��O\��l�?�ұ��_OI,SMQ<�ϒ ۋ{Y�\�x�����E����A�GO�x��S��d6�H3��V�P�e�-���ik^�9{q����p=|���ʵ���\��K�gۯ�_脼�}�CL�F�#���FTc�a-,�;�D�G[Y����]�'���*�q`[��M��r4�e��E������6CP@�R=��6��Hި͝��ڛ�*��r�T.����p�g2�h���S+}ug2CP`�^�����4T�4C��~&=w|����A�*9��<"�a�����6����[�I!����=B+9e*ƚ9.�0�ш��V7r����m�L�����4��c�Y_=.,���x)C�
�@1S�v���gT�A%����� hdec�"Ӕ�3�(U?S~�)�n�wb2��Ӧ����#ch�	������4HQ� ��b�A���iW� 6j��* ���<@
`~�
-� U�jTz��I}^���>���p���nO���s�u�Z� �L,�؝�0˃~��i����	�(l��e߾�8��}_�b���g#!����r,�.eY|k��L��yƳ`��_t�+/�\޸5 �;�Hg�g��I�rE΋�m�Z8`�>PA�����l�\�����~o��<�!XA9��ύ=���W�)A1�&��:�x���a����d�����Hg�͖ʹ߱M@���4�8�����uw2/�ph��&RѰ����c�̉�(V���R����C���!a9E���n��!�z�Z�g�k~���ʖ�b��JtA�\h���˫��2�C0��O���
b��"/&U�ס^��L���iB�q��q-����FlM*�;�N���9a�>RT4w&��+����P~�FP=�n����S�������A��U�@��5�"ay�Ê%4KK��T��:uؖKËo7�+���t���;=�c۱A	-��{G�-�T��_��
��B��$i���ݷ�N�F��g`E�e5��4�/s98�V��� {+G��\��>͞����%
CRZ��OWw��=�z�h���s��J��>��P�4r��%����ݩ�y������Z�q�-�_�Mr�G���3��~�ݣ`�M]��}��+@���&���H���>Pp����7B�!�.8�~SP��(+� �F�@�&�gݛ���� ���2�lC�mX�a��!H�	�Yw1��)"��4$P��.+����|Sz�jty����g�,)��m����C�a�Ʀ"0Y�f�l0o_������f����֢��i ?Iw���y_R $&_j���j�F��A=D�=
�F���.��Y4K$MU������\�ʱ�x�=n�bKGV���Q��A�*�Q������b�<��l��ITt�1u�i���g\kq�5ۙ��_{�yA\���s/ߖ�?0ٵq\̗R�X8��Q{�#�<��Z�D�<L�V~�\)Qs�t�<�c�����.�<�P���UOz�)-4РB���f��>�Mq�R�{����E�ѩm�D�����+;�v�<s�S�^����<�j�Z�s��E�֫k����K�e�2ʹ�h�Y@��~©k�#�7A�\@j��	��'v�X�xI����w\4�N~��
��w
%�&X��q���h�:�TY�6�jW�������Լթ9%���B+�һ �X��5#s>^�־y$/K�}��:nZ��b�C�o��o���  J=-ykH�|B?�э}q�>M^��:��)��k��!v�09w1cx���$h�u@m�.2AHC��NE�έ/,�f�����9W`�|���7E1�o`��
v��l�+�.�#�Ur�(,`�X�
���}��l��䋲����!�V��IKy�:�8vY��_�w.b/��-b�JX^F31~̝���F"�K��3�cB����qg�DNu��o�Ҋʇ��Kc����4��W<[|d��k�e�V���r'Y��mQ�E����;�*8	^�[6��T*�;ᵁ�Sf� b�^=�f#�k)���ɘb��2r����DE�������Ph(� 0��0@��$Ztx('���z���}��&���R����� ��Xv�+�F��~��7�y�p��S���p������H�>gb���
��1H.+k�4��Q���`�}=���0@v�]2�@���Xܦ���͊p��!�P.Y�up��l�["]�汚�n-	����ޙ
��Z��j��t{9��W�����"$=:��J�p�H�6��۷�t�����gc�0!k]6rs�غ�@�e@mOӽ��?Eo�+ٳ�IL�[�A(A3�l���dI.9�����{��E������]xIK����x�P�����v��Xb���dS|�'�o�C��KX��d:dr�6�L����'Jd�oH�Ǡ	)+&N�VT1���n2GG(:cC(߃��0JY�~ �As�h)PgWʑ�f8�~�'��jM�O��&�r"~���]�Ul��Wؐv�����(ܪ�ב�M������aM�B��\Ŕ��o��O��`������6lW2cB�s�O�+q�	����	����W�u�z�5�_J�vE1��.qT_ P&%�X�e�6���3�	F{*eA(8�����m`$�ob������9����-KFun��ں��
�pi��9k`��E��d���((?�I(i+�{L�JzEmZ������j�] ��=�G[�3��U�bQ(6T�.}C?Fj#�U�$�
W��޿���n@�7d��Bb���U�F��F��4���Y3񓠪<*�^��n�[�g��ag��Z�6�jTb���|X��<-G��?�.�q�w�@����AΪ���6}�\��q�`�qn�#�N
�G@$��c�Y�tbD�6ں�ѫ�7a������A��W%3B��P�	�\�˯�c���T�.�H������ ;�1R�ʊ�>[�g~�?�q�{��>�̓b����$Y�\�1�BqV˜�"�wI�����~��>�#O��酶'7/���Q��ւ0��q&0�Ç;�>y�:�#5X�Ƿ��`����x�e0]���e��3�?�ƕ�S�\��:L m0��R�Ih�.��?��� <��A��wS�D�8�����y�)�O=���B��0�]�K�^څ"g�����LE��&?7PJ�&G���@k���;���
ø1�)<�"̗�{"�)E_�/�hb�� ���F���:+S&��#��-���S�<QҤ:�ӧ����? 1����h���ČR�V�0HF-�x�����q��Q��&�d��ӹX@˗����T���y��bST�K��M!�&Ҝ��Ƚu��� jK\�w�5ݺ�I��{��ɭ4�sXi��&:HU�hQ;�>�С>g�Q���0����Q�T��@lT����Z";��r�E�K*���Y说� �[t;��Z��%�?8s�b���X� Y�w�t�_;;S�����������L�Ұ;h���kl��2�VU�HJ����O�g"*��D�!��B�m���>��G�K4}㔹̈k%�뵀/��:����>cs�H#Jh��������)��� )~`�
	��%�D�s̾����R/Q�2��FA���FLΩ!Ҏ&:Ww2C�fj����WTS�aDt+��4S���Y�|���i�O�9�g�o1�9)�`�N玟j�1(9��'�Ʉs�Dn-.
<8=_�Xj&�٠���)5R��ړ}�C����x�LMh��o��G�9�{��������9�q���?�� �5�;��� k4d�d��I�1%6�S,f9���-�������8,bNXuՒH�M�؉p�z!k�ZW���s����mm��k7�_B$-�$�!❛.����W�Z�ݶ֮3�.�����3!(��8y�'�zA�3��C@@����ݳ�7e���{is3�Ug��.��d�
�`��=�W��;�����ÍS�wA�;E���#��5�L?�k:�M���fM:1�Pkej�@���p@�:������3(��zk����9�G_��6��`��.��}��3��Zɯ�Q.��( ��q
O�+v�2)#P�]m�:�R"�bbKs�:��!�pG�%��Hܘt�&F��5n�-M.A��@+����D��!�UDy}�>�`��2����>B��g��r84�4��ԏ���t�P��_�K�ʕk���`����pθ�p�'D�H_.�p�y^5������em'N0��t�@��+g�?�Rr��͆�}�y �5��M�3i�7�AH��sjX��.]@_v;4C��m��N��̿ZMH~p(<V<�mv+�$��n�����a��<�c�ٵWn��bzKQ��v]+@2�ZNŅ�5�J���z޾B�+O<F����s�,9�0�F
�!�{�C�7���Y¸N�)���O�ʌ���o���������|C
�ya�H���s.ȳ�R�륏2+A����Q��~�� E��C���`��J ���pu���`D۱�L>���PQ����²��c�\�`k�c��?i�]�茡o���訦�B��Vu�ƌ�P	��Ls&�8��	���N!Llv��eu\�3�F�N&Nf'Kt�݌��k��RkHˬ�y�L��m���,�S3Ϛ}�߷��.�U����Y�P"��'{����e>���P��a��AB�aa| 97U�l���nZ��jwMy�#qN���C_��]ZU�7������-�(i]�qo�N�1�L�O%�<@�}}n�O�~dB�Xd�m���ꬾhR첰7J�A�XF�4�Z�b9��3ı(�0��3V�c̡�?���<*�;n�U���ðB��TL$�č�]C�1FYd�{=�0ny��'d$m��X<��U�$�쳱%ǚ膲�2���O�B0�E�a��!4F���M����f�j�A���`���k^ni#�Ϊ_���XoW}\���<����S*�[�1m?�x)�A�ow����ݷAZ�"1����������IC�d�!�J�s�_��'J�}������U��P�������*�Rۄ�Umy��������ja]����{�;���Qچ�o��H�V�A  �9Kd~C��?�-
Vx���f^�M2:�]����s�ۜ�<,vt��`��T� �b^�F(��6��=�����H
M� >��H�+Y̓�p�E��pGx=��{̘j[�e��(��/�qE����x�rE�����#�E1��I���c~Ȁ��g���&E�4?��e�E�W�p�{zT�����в�x$Ԏ���
�
\y̒g�XE�79�в�wwzt65}��v�=�eM�8�U��Q9��f��e�}��g��	��D����4�b�����Y���Z�PKMXv����_�x��^�'��W@�#�2@�Z����Z����&I.��x��GW u��oN7��xR��,��*D��x<���c��;5c����݅V�f�kH�����po�T�?��Է��`�Q���!yk�Z��9���	�L�d�a�PF.�Mr�F��=�M���40Bwx��)�.��k�|�jcj�f�e�q��7�;���jO]$�*j�~��y�K��F��t��[�0f*��K�պ�S���ttM"r�30*<h��Ŭ21�ZA���J�6�\���m<e$܆����[ϡE�
~����
��oQ��B�̽L*%�[r���������,Yh3�Xp&�6v�!ϯl:2u��h�Qkmn��|وf꽞ϿǮ��=�Z��s���|FEA*��`)G^x�8"&!�D�,�t�l9���J\^�_b��`�i�i/^N�>0��kN��v�N%BǯGT�6|S�HU9��t�Ü�i ��i����Cރ�.ܛ�X�ᚉ�ft��UUr���p'�%�͓C��t� E�#�\�3N5����lh"�j�Ɩ��,]�Z�G���!G��(��VAR�f#9�մ��c��)�3-��w�D~˺�F�V&2��fS����2������+�A1�{C�g��f��'6�6ٔͶ֬W)@��EH�m�U���=�D$,"�����O8Oo-��<��#/�\w��4mP�c��̅4�b����D>�C�ue�toƵ¸fm����{�r�l�GP����}�k&vq�+�5~�񡌗�ǅig�n��WşMɀP��V\�^��1���%�6�C��l��b�I���N�&_�h gD��cv]1uA�5�.4�Q�@<s���7}�/s� ���{><�7gh�L���ل�:�֮��eFWK��#:>1�+��a&�JK+':lA8���c�"X<��\FQ�֍�N��k�oó:�����<����vs)�J�����23<aωS��)���9�
T�Y��s�� s�Uc�.��� ��`�=�d���:��j}�D>��ω�	 F�S�
�������.��o�?�
��!�{X̐��=@��L��̚�WP�5�;����ץ@��n]�ЉK<��Q��W3Ϝ=A��|�m,��Z�����{R�FL������E�1ld��$r������3��=kW��X�rt���)C~w������ҙ�*h�����kQ帰�9[1Fb=�\�mD��6���`K�x���D�<�;�;��6���G8�r��O�2\�"e���� %7��S��{�ߎ�_"|�a�(�Cs{�'��owb���D��ɚ�Թ�����Yy�@��RY��q1D�eg�Hm�Z��b^B��缣i5j�Yr<��L+��M����E�
]y.r�KΉ�$�զ@8��l"Ґ8���}l=q(LJ[9���nC�ť�ǎQ�bc�>0F��a�u�z`��х���ȁ��4b
I��&]1�U��vv������w�b?v�]��_�V�g+r�BTR��S>���-��P�Ijg��X�c��G~���_W<P�bY�u�,��#�1����l[��^G��!u�0Ȭ$2��puؽ�,l,ܹ,�i'�"�T��(E�7W�Gd��pm�K.,�Ţ��f��mB���v@SK?Ԩ�`�^��d��8X�g���$<�[~�;n,N�����|c�<[& ��a];��ݘ���~�8~<7
�E����܆���9��@<f�$msz8��~~5�<�e�U�����e1ڟ��՜`]H�]8rx.��Ǯs]������!͟<�q��p�.ܳ� �������g=@
����l�k=y��" ��86��X4Fסr��3||P��w�u��::n�Z6l0���(a<$�5 �^q��q&�E���5�v��H�U����ʩ��?�O�\�z���3�h�a�p3WX�I�׷��t*�<�pj
�ە����H��?8ׯ��6G�H$+��ۯu]�l��:�={Bu(�V� �FϾk@0�EJ��̛�s.(��İ�!�0��� ���g �)���d,uoc�j��]��0AΉCN����)a�PK��[��PV���l QQ��5�F0rE캆;�P�$�D�`a�ɵo^�9u����j�HD+4��PW"'���+��P/@Z ��`��I�֚� �^*�C�g~{���"�]����2�y7�����%e�j���ޛcS���?�af�X+7_�;U������	'�6Z�8��>ɚ�k6�Fx/Y�97G��5f�g��Bk��1o#�1�������yi�,"���8��]�c���Sy��iT.E�����kQ�xud�񬿧���QT��.߹T�F�oQ�*4i\�6H��0��ڹ��E�}&�Fu���$��KT� h�#�*����ұ{\M*�v����Pa��|K:,����#����}-CN�/"5��C4�:�T&��G*�P�M��pfSĩ�$����ڰs�z�bd�����˭��V��MY:g��b�"/�5�H��N���z�.��a�[��EM�����"��v�g������>���;¬0�q<�4��M����l���fn7o@�Km�t�HB7��F�'��;���o7@�
�2���#�jR�O�v�e,���Ld1�.#O(���o��1�[��{6�vloL�v#J��Qy~�z����<���9Q�a�[�ӥ�J�	A�4�-EG�<�V\��047�f���]���^y�x�M'v�H���WƳP�o���s��P�-���$����
J��'Q�� 2���ڈ)Y�?-⩆��'T�n�d��RD������$���/� 	�U�{/��m�w���&�_E�Ǳ����|AR�g�޹{����;�j�/%c����m�VC�9t�{f� ���-b��~����s5���2�5p[��Y�PQ#�q@�&���e��X>D{Ew�t�Ϟ�t^�)M�lXv\R����9���^��PQ:xL��[�.��U�XJS����[o�4Q���^�;pS�~�.H�>=G����uv�A]��c!c���n��J������z!5Қ����#���f�}�L��^��p����r��:�Qn.�t�<���0�x�e2�w��c(�?ޮ�-���l q��a��7E��i0 {�s�N�@t�qBY�ל��ũ�R9�c�Qc��wG�{������0���N�;Qj�tNN�'��7X�� �'L)�(G�]vdO�R%���i�L�4�nv�V�&y�h�8E��pQO�{�'�����-��C'�k�%6iE�暁"�c,V��4�Q��ׇ��0
��0�B����}���~ȟ6���^sj��
j�c&;;�?ba1�����f~o77�m��\���3��~�[��re�CLL�m���w܄<'S4e�L*�|=6Db��r���V���K׬�M8ʶo������!y/E�r�Q#!I'�k�C�zmIWg;��oiRozc�W�S�6��%��E�s�a\(-�+2�FL�X�ySuא���b��L�#�K1�k�����n2Q�T�@(P�䄛"��`�����F��<���RI��AE���5#�c`�/��`��A��w�bN4$B�|���,I��Ui��P%o>�ط�EBτ�Ni��4c@1�v���^SF�P:6r�k�A@&d�Y�u�����3i'��0�4�
`���/9�r쯧-[C���=��6*V��&7�C'��i��Tc��Θ����ߎ�
4^�#��EF�� 0�*�80�oYY`|#b}
x��'EԾ�ry�UW��L�D֎���T�;�i��W?�Q����NJİ�1i�d�Qr�V�{��������s�L��Մ���\g�xs��v��+I��̤�իD�*�/;U��@4z��O��*Wo� m��Y��^i��貌�k�5a���b����2[��Moҩ�HL�|�7e��/�1�����\r����qL0D��?g+�BRVdi������WLx~m*G�oI�f	�?�h����&����$i�$uZP`��3lc�L���2�<�,���6�)]��H2e��W14�l���z_�ӭ%�Y�>���,v�f����9��_��(Y����:�(��i�zA��q+��L��Lc{��3�U|�f��������M!�����Y�Z~��`�f��5<�X�<�'�PO������R��x�f׎�6{���/�m!���t�D�����kI��S�EP5퓷�fӈkS߲c��B�ޏ�ǣ�3��y=u�����igF�nXz���w��L�F�gf���:��51o�MH��(����ቼi�3���Z��?�o#���	�����D<5���i�����k�p���o��ӄ�<�mEP6���]�t
"��֎��O��x�^�����&�����9��o�#�o+ڍ���X������ڠ�BѾ��\�ˮ6�m?�N+_�Vx�k�ʐદ�$�&�#)�^~�V����濥��X�8��_F��h��i�ibV/:vMi9Q��	�-*A#�y�i���=	!���E �/�/!�&-c���55�-_LYv�@Sa����������\���{�!^i��d&zB��\�p݀�=���ͪZT�8q�<~H���v#4�8�gx�T�I�>�T�x�⍓��Du��(�bZ~)�Xv9�<E5%�7��َbr"m��B�s��ef�=�+�ͺ�|s��:>���RyUDUΧ��X�+FII�����Q�|�6�R�yCԢ�j��'.��Q�i����k���l*I����4vғ�X�r�^˃�r3"g/�A�X��V�M�GK���d0w8q?H���0|�����$�-<C�d���g��Xƅ�,�AoH��񤞮;؛i:�*�'��vd;xi�d�ݿR�v
�	l�m�,hc�Gu��(8�d��d日mw�=��*:mhB�AEB�Z�}~%R�Q���]^���͇��f���Cm�䘊�����e�K��])	!� (xC�^�:	q���[�V���鏫�g`�����H�@G�a����Y�4o�}Z���(H�su����.�4/B˗R3<�4i	=�Է@�T>������ {�[�zǠ!*�jA��q�[�]3Ց�>_9'�|�����1��� $�ߠ�F
��OÃh]�4�o�3��5�5�_���̖�hD��|`�����+H^��!ຼ�BBhF��sd I/��2À�	�A#9nQrZe � ����3�_������e���K��r,�����3rΖɹJ�����g�}�S�1@9�jfm��_'|���Lt_��B����pw�~��#;�dT��|�F���L��4��^���J) ��)�9r종��K���R�Ք�����h�8MF�y�:!�LS�~w�0]N�E�=�r�qxު��A��9T�)z��S*��b������������q-�Pir�x$8,ͭ����J���H_p��g�_h����r��1L���n����O�p�o�gm��u�}�Wb��n&���) Y׺�9����?���q�=ˉ�	���#E�bu�B&��{�����vؒ�G��� _�����`8\��)�6���r�~rR��sT�:�0n4M��e����˧����t�Epœ=���(�֫a���Qv���R�KLB��'�	"���R�D�3��q)(��퓀�9�@�q��WAX���1y���(��_�l+˿��!���!<-q[ӯg(�ƫ嘄L\sQ�V�O(��"������� s	VJD(�*i���ROX @B�5g=����T�_�v��#����B�!U�ؘ�6J���+ �qF0�M�5?'G�R��Z�ig����ظZ�H�2����_@f�����#0�����(ׯ�WO�|�RQ��
�ܰIF#�H]��2��D\mC덡2z��:�n�Q��)�(�ּ�)�-�-��\��i�	u����T3q:�,��s�/h����A�
������Bo����>i^�TLa�1{L*iXI��r��,��j^�i�����`���wס��(��o��F��,]�_L�Q�Z�̹����>DTq�J�s3Zc�?�~l�yΏஏ�����qJ�3�¤�繲TݍB/r��R�yI@����b<�������tRQ��i��i
���)��ʚ�t�F��d�u��M�-�ɳ�I|��E�3�;�=�Sj+�>����}��Q	�ƻ����Z����$z(�� ���5�d
>���S�z�&y>��<���Z���Wb�3}Ą�Q��-@��D���i���(�@W����ܘ�b��kWXcqC%29��e��6R��r�C��ao@K��3a𛯣������z`ahB�,��fݷ7�W0 �_�������cO�� �>cn�\��a�\!��gA��:RMX��H��y9���ɂO�=uW�D�D�w��T�(�}��C0����u��$>�^�a���˓�Qh`�qqpr� G�z��׬��A^�l����&w5�-{���,�K�N�|`?�5p���J�"н=�8�N}xuf%wz����J�#,���:���4�e߳�n~�gŉ���J��g`fv�+�����ŋpw�]�˻D�r=z� ��R���>LB;, �$0a���Nx),L�X�D����?o�So��rȽ����F��R�tL�J�aǬ/ܙ����y�`��R�e��:��>&Sn��!A05d����Zs�F;�Iӎ�|_V���	˷,� Y�0j�"�<ر(�Xx�&jP�4����5�ӊr���%�2'�w?#k�e���]�TR^�4Ué6#]�����[ :�-�λ�ep�f��Q�����������B�"ŧa�|| �8zˊ��P��3kxqN�d��5�4���1GR)?��5ř��J�*��5��M����GD���^t�v�� RG
��z��i�@yr@��~ѷhz���9�Xɖ�YkϼʏA�9:t�s)�=q1�L�o���i��h;�G�#4��w}{%S�j_5�q�ߐ�3_��;��;����A��4��*A,&�|J�޽��֚�^��P^�<6�3�;񖎯>��	�m3��'���-�;ƺ,xS �����2c��ge	C��2K)i!��,b����+6��t~=)6�W�}Y9�`��{�ܾ�'�x?@��=#������#��}� �\��ErQ�Yo\t�un�mFA��2��=�!5p�q��%�Y�rN��H��N�oDJo8`��2��Lv�-���c���Ո:i�#�`�;ԫ�F]K����Wv��/.{�t��<Q��7�T�}̤�_>�i���i������bs���9��A^�<5r��/�/<%�֙S?��Z���.��Sl )�X�*l����LUǕO�☟SR�)2�?v��vsT���I�k==�?!^��t$�I�B������f���p�i�}��k�W��}wNd�oֵ�%e,�˚k{�!���M嬤qX��k��F�5�H��y�+7Ky�]�"���"]s❋������>Vj�]�#y-H�9"'��:q�i�O�׌�tf��S1��x�@ʌ�%���aKw�N�jK���7�	������f��o���Γ���bak�;W6ڈ�f�.F�r_������{y��}��Ms}٠s?���@1VK@Z�����fػ�o��������0>���[��\K��]����׭�k��0"g��na׹]����v���3�J�]	u�Z-}����M�ƒo�;|�^}���5�`�h���Cf6�# G�	у������ߊ��g���㷏M��z@��4S���I�ZNaS4Ų�*��͜�c��}O�_�O�l��ja�2�d-�e��A���&A=�_coq�_E9C�,B�&�*��q3|v��~�O�J񑷰� k�bʔ^����ʈ�c+��?t&0e��F==���%f�X�w"���v�>�Y�J|�3��h�Q(�.�_(6��D��qInx����{{_��54Ȏ�&���D$�q>B9�zI�y$���^SÐ]�[ۉ̭s�d�g�"���	*�,��[]q=����ӈ��,L���*��5�ą)=�����Qa�����x����(Q	���G앨�k���eX�.�"�xO������]��>�l�y�(`;[�Wo"��W%s>E-��3A�'�E�pk�_�����)P�Z�"�QD�����|�'��UbX�E%;��j�.�M;'��1�uք�	�R�J/
� <&��4E��41h&�֪Y��������ܸFʅ8��6q8R'��c7�|z��'��DФ�@{6�hX����{�#զT�'m
 �٠h�xЛ�W��G�!Yո$q����HH��#��V��t]�e�a̜Z|�8�i��BϏ�y�|n�/��*�����Ӕ����J>��[Pu����ɟg� ���3��d7{d]��q�����)L	���(��ﲘӈ����g�	�ήץe��l
��ղ�F�#D䥿e�p1.ʛ�<�q��=�N�V'Z�IN��e����"K���R�70i<o�*[���0>�@�x�Y�ވ�y_b���x�5Pg��q֣��IDsT���7Yr���I!�T�IE�z]D�]����		����G�����}��-=�]���r˰<���7@���D����O�����(���G���ˁg�n�!?1^-S��>���'�|�-�~̃fBUGR�r=%�T봡��'Z$��@8�����Y�O��D�+)zD3��@��]���}���li����>�'�MK�����1꫰7�ci��0u�HC�k�K�m���ʨ�|������K�����<ך)d=<̃S�>��8T	��c5(f�ˣK���q��{v�����Rh��yE�{�b��۬]ųO����̸C���vts���ة]4�g�%��*��L�8y��O8-;$��=���a����Nu��K�d��� �� гJ���e-�Y�s{W�}f�8���w��I�����
>�j  ���u�Am0yfu 3Zlb]AQpz�`��H���#�-���SXBvxLeJt�r�P�7}�-��)7ջl���F��Y�:kTr3a:=�)
8˱���B1��d#��I�z�ԍX��7{�Yݸ�@���#PD@���{ڑ�|�'h.\4>M���a�N��6H͊֟{�FȒ�+����;M�nz1L���2 ��&��?B��OS�8��?㦳0��R��+�4XIQ1!�:��t�� q�-q�g5���*C:T�)�~�>��nʃS�� *�y�/�a��	p��~�q؈�S٩�ی��T �6d���Flh"�Zӭ�cW����gl��ҿ^R9�B�`�^�y
�2�K�b�F�y�GQ� ��F�)�Ρ�3�[��F����Ɖ�P�ͳ�ST/��)��d���69H��R+�E�97ݶa���w9%dOs�u~�P�Ÿ�G�jjR��M�"04��?�A��d���b]�L��eG�/+^[d�ݖ�Q �/I�,̧�́'Ӵ������bK$p?K��?Qg?L(9��F�3ۭ%�ٲ ��k��-S�����򠁲�"�]ܪ����jI/u��4k��l~�~,؅�N ��god�k�{!�F�t�7������{/ed�>E�3o6�u4�ɊsG"�:�[���R��"k�E��b��R������8������뚪.�ɾ���-l� 3n!j�J M:y����=/��<3�X�:�W�,�M�\�`�:L�o�T�a
4����^J@�6��-��=�)}⠤M��7��ᘊT���D��TS����|����,j��f��u�\�<���7�1d<����64��*���r�5��E!�q��ݖ��y	�PG�-�#o-�!@�VK^���=��ԉ�?r0�&�j������J�8:b��*_���_r��O�
Π�,�E*�y^�����b�=���Z"b~�3?!��d�������� t4�A�Ѭ$p��u����B���x#�i���N9s�rʌ*��|��!|�J��_^��/ֶp�vgX*��+���{��X�$���<sF��8��RP��覴������w��8~�;P�s�t#U��R���߲���tr��%�S;ؾ������������h���.�a��2Cpa �"��<�x�#��^��v~*��a��Ο���4��Pђ�-�x���d�6>n� �kz�uTB���8-�'X~*��nԷp�fX$���|V,jd���$O�|$��⽼�Ǩ|��3�@}�I�01�Q����۞ʵ^���I?�l8įN�r0�����]hCY!!g{������m�����֧��}.ْR�u��6Ǥ�Z0@�ё��z�j#���Vƒ�q�7�ts�>�Tʣ
٬�(�*�P%P�."�A*J���'��b��^. ]��_ZDA{'|�+Y���e ��t�|":�$��>Vq[3?���w�j᫨0#ҋ�w�σ��A�E1I[L3&�w�_�w� a��A���b�~?(�dD��S:��Tt��Iz�22��ln������A���?
��ic#8�?F��N0�|E�Q��K~�\?�9A^��[틻D��u�ߪ��4�^�_����q����X��ɪ��*e����TI8�7��5Y*����Rֵ���(c���N�R��eY~i�Խ�ov��>�dAje�a �bE��K�H?��T�����{x@ǩ����*.����#��E�����tX��-k��k��n��$�/6�p�l�V��@�`�2�81|�T�K���s� �2���.Uҳ�A��2�e���B��yE�~K���w���UUC��d��Q��Oo�ޖ��GZ�&�N;NDIW�rV�v���p	�/�����%N�dA���C,�	�aW��n�b�ĵ�W5s-� W��TڠI/l�ig�W�MR~�����n��>:9���=k
ڔ�M��;��m	�!��)�T��p&�$Ay_�b��>�T�eN�~�Rl��]�M��̣p>1LZ�tl���A��p������S	_훚�NK��F�&�q��zl�Z̽X����UJhJo4�ۍ�h';"�g�<U�Ӆ���L���1�L�ɝ���G��ڹ貣j��-$��Μ� �ᱡ 8��Y�L��OF��!�$�d~v?�0)�1?0$���E¹�J��X�_/����$��n.K�!_����J��{�Y�qlv"�S�K=D��J@���rf����.C������qP���|TS*������z/2��s$Y
�4p�xmY�2h���݈��J�Jqz1�;�zΖr�<\"=����d�n�{����K�����W�l3P�769VW�Uy
K�X��/��M�� ��z1�j��l�o\9�?��̀;>:��b�� lz��zW����S� �����D}�Δf*wbN�b���E���f-w�<�nU2���]�wY�3��~��&4xj��!�+(@b?�Oץ�i/���V�B�p$��CT���p�h���3ţ>�j��8-b����G\R�����$B��Fɩ�r���)D3�|ES�'��LF��FA��\�5JhQ$�V�6�B�ͤz�P��pD�bǾ�SHh�Zќ �Io�+ai�Y�h��dNw�W�\l�t���hb$��M��s+a$�P����RaV�:a� ��8�lljg0���E��@,����;�8嵟nն��?�E\���[�#���Q���M/l/zw�@�q N�W9��	P�{*�e�������c��f/��s[Pl�����f�v�p\��X/jw0�6ò�
��ʽ�Z݄q��{�����l�E�zQk���zKBw�Ƌ�3�_|�OQ���x�&�澸9ew���2gwːn�ǈa�>}�+���I"��TU�j최h����̓ȏ*��t)��fƍt���+>�c�>��0��5��FhR����[�f>V�d{�l)$��7�,�c��~�l��El�v����}�}��Ӗ�y��y���q�ը���ܦԉc���D͍��)�N'�:�n��y��܂!�L�5CS0eޑ�A�(����?5��������2 ��x�u�](�V�3٘��K���B5�G ���~�ݡ�n6G�H�2��0�k ������Q�"mc�"#�歖ެU|�}��3�קmoS�>J�Oq���u���[�8�)8E(�W���m��6�7lHt?��/M��G$I���R�bX�es倅�;� �ֆ^�!�f#2�<�<`ԭ�����q�h+�im=#$	�k ο�_qZM ���%� ��������Nҏ��=��/���D(�9	�~`��/����K)��Mu�;Ƃ���u|S�MP_�n�FѺƛ�-�
R�R7�.��Q�mx_�0B��������Q��w��tP5��Ni	K�Û
����<]3��DJ^*��R@$��J[���D����_,�a��-w���IA�����׍�s����7�����b���e�#��ۍ����5�¹ubO�kB��.�Q�]�X�v�����i�{ԡ8%z�`��{��蔛�oϨ���ʔU�7h �y�S��۔?)p\]%�D?�x�F�����ψ]��e1y�����&e,�1��~�u�X�����xV"�o�<������ �3�I!�<yc�!���� E+��vG�m�5	�(����C��֋�?�-f,��u1�C�P��\�������x�q���6��/�<?eN[��i>�9�3��D��:����tM>A�Nl�����u0Z�2�3Y'��m�4��
�MS�)�Z������;k^� �pA~����T!x�C*=4F�j����A��ze����A[!Z���t�l5V�@���@[�uo����O:�g��������I�{��%�c��oם�m���B�WwzK�z��b�E���l��0�TNj���kND��-ފ��>V�kTM���k�����5�."Ě,����[Oek8h��Xz>FL>�p+	��$TXͬ���Yٯ�{�o�qF	*g�9�H�p��/d�N��.�bx��ő���Q�BBi���$J1��7D�tĪ���F-�_�zːS��� N��7D�0t����J 
;T~۶I����������4�o@�sMFX!j5�>��hS�]�~@a��NS����ںӘ��᧝Hu"������"��YwF~v^�3Kf��Jj�\= ?����B�����������~/a�G�-p`�Ҵ@���&LC�ϵh@l�K��я�4�,�缰 M��V����p�@�Tc�x+� ��ͩb�V�:�	��=Z�W焝rC�;q�!�9��H�9B������fQݛc9 '�U�%�d�5�oH�ٞ�w��v�y(���͞���R]�"�]&��uNb��a�+	�n�D�MOo�F���Q��G"/��Ҋ�1���]B��NA��<�J��WC�[�_q���X�߁�5"��	��cԿ�TU�Srɰ��R�cEBI���X=�w
/�	q�3'���J8�\4�-�Ƣ���sҬ&
k�:_��+�9�C^s����J�)�4Ф���s���l(�P���G,#mZ@ `��5$&Y����配�9�`Ia7����=��l]W��R�vͽ0�A�QS^���tⷐJ�����r��k\y_B\�^Y��P�,��<@�GPNA��g}�\���6�N���5B�Y�)n��ln�����[�O@��d��"�qI��*r
j�4@Ed����y�&̔-k73��gW�m��j-�o3�7\[��|`�P��/N�򛵹�8�Ã�`�<�nn>��<�F��ņl�$��0��_F����{�2xE�}����jD�mV��g��� F4�J<́B�.Wh�iɰc�JD�5'���L����^�R/�W��#P/��@�Q=���;�!�Ʒ��g��`���Q�L���i�أD��I�^��mb��(��G7��%�b��@�z��fZ�꧟b�a��ǘ\��u�����'v���/,V�|5�#δ����䰍oMSf#�]�ˉ��zֱ��c?�ܤ�W��wd�S�h���f  fN#�I�{��Cfc �Z4�q���RTk�[�G��E�Yqj[t)�c*o���F� �kP�×�>2���V�����9X�I����@J�{�h�^��� L�ݏ��=_��*pp�@R�{?5w-��fU'(�E�=˩LS��<����q^�Z_�ǂ�Y�b��9��wѬtO������}M�w�lh�e�%��q ���߂y5�"�Чc�)ҿ���F����:wx|�k�S�.�7�ՁPs�E�_�>�/@m�O'HEO��i�v�A>�t	���X[�a�&����&�:И�/-�Ǣ���?zd����5R�X�����?�KY��z$�BV���L��z�a��p}��X��zB�7!��?6������E�M.���+7�`�(>���5�2Ld��s�y�R9�#-Ia��]�S����*�5f��拻�@c�]�}Ww��Z�����u鷑�3� ���z��tnOȜ���XUp2CgTJrY �uxd&햌W��\@.�k��EL�h��ڰaO�U��g`�a�U6��1 Bo��
�|sN�b�>�X��>.���Ah����d�O��r��W�ܳO�=&�/���~�6Mh{!0���A�����]�3M�s6~�<�7��[��_8�d�yKI�ǟZ��~fr��ؼH>�f���W�������PE��O�}�k��K�����!��pT�Ǽ"�^�#����8��҃&M�'��;�2L/�)i�K$g��T��}�`���h�,ز�p
C9��AK,\XY�	ʲ@�r�����7Ֆ�#��PSM/SJ�=4T�*�H.$����u|@�K$\�A�?%ʂ���%���B�լ_���)�ߑ���N�94���V4N�8��f2DM b�U-� ��=z����)� �;��C��(��~���|���OQ|Z��ێ�p�M�S5�����Q�S����|0��H2�\�B��o�@Ϣ��å��˿%�!���s����	a4RHUoB�پ���8 -g�(���W��ZTMֈt�˗J�m[��E,���F�M��JĨ
Q�U"r����(D�����7�]˶�(�Ts��f��3&�ک�a�;���Jݔ��bICμ�}�p�#տu�aW�+Oi�������������y�d��z��n�����Ȧϒr݁C_".7�2.U�e�F�/�����2Z���8b�U��l������h�p�_5��G�e>�g�_Wkd��,���&$H�B̧�h8"���׈8�vn�D�1):x+��2H�N���t�M��@K!��r|�[]�bhh$ʇa4m	��l�5k#����01tg"�e�c�!��-�]cGJ��ЪH�[)���mh�W���sY���*�D:ɶuGA�Y�E���A�8��ܘ�ҧ�����䀬�s��Qi;1����'Ȱ����$��B�8��YѣRJ�P+�X���~��D� q��%_� 6�Q�֫��k	��m|�/��K�gq��w'����^5״Rf^�؃Q����)шv�"���][G�g�ж�Q�B��񎪢ᮯ+W�0���S��2��#�le�!u��)�ԙn����;��N������������ʞ�>��IN��Ȩ�q���jgA�2XJ��.�^m	��6D�9ho�a�֣iJ���7�uV���Oz(�8�4�o��$�v� ���y���Zٷ�N���sGܶI�?c!�+�	|��֋�I�:~7.I��.���mDA\۝o��kʺ�����f����b-�<n�G��!�N���a>~u0�y�[����r=�i� SD�������>F<�y.=a�g���H�"oA!�m���[�!E��X�|o�lB(�7&��`�b�5�oM��NXH�ޕ����׉�Oj(Y�ed���&O�ͻ��ƮC��?�F^kE�81�K/fg��b���C�i�`-%uv^��E�Ε~��X��i��W
��A�c��qᏨ)�;��˶�M�c��q@n2q#fї�c��-�k�M-�g:}߈^�[����ovW�]�ϩ~���:��ї��j����p���5�[����b�c`��c^0w��\�]e�G��ן̫r�e�8���o5,D�H��u������BZ��*�:+�q�6*s���U�'(�8)*��=��ii�2���̋;�m�2�(&m���^l[+�j<�kN�<��򑡶Nw/1s������E�y�0>�3��-3�O������S0T�x�J��N��m�&�ɟ�|V��UfF5�	i�\=歱<����E7����x���^��#�q�3��:�S�̫~��0Lu�K� �^Y�yCk�@~�2!xN�^�A��u
H���9l���`W�ٌ�%ܛ[E(�XQ��y �/�}�ꭈ��I�iUhmTQl�&U��2!����
q�&�?���g*��Fy�*e�x�{6�ѭ6F\����3d�*�E����[�\�udM�h������0�Zdt�C^��J��nP#����
u�/g���N�d{�P�k�6� v�QJQxID!��*J��^ȾCA�xo\t:sQ� +/+�B�Q���9�w���!�:7�׍ Q�Ë�Ng��Gd ���*�:ɋ�xV;���IG���},�7�g�b��<�.�襰zK���DQ��䅨�KԯƯH����8����(�������;��H�4ѣ��-6I�j�AR��c*Cs��5ᰭ/s:�D?�E����t�Ψن�a.�/�c*x�7Z�m��
�K;��*��!�֨�6r�����P�M�]{�i���Z-���E-�:|������՜#���4ΪX<C��q�^ů8�٢�J��4�������=� H���&O��0[���� $��  Y�=�(�uS:y}z��v����u�5+�#��u���C��_D�\�
���Ȑ+s�`C��6���$-|�f��5�E<�K��
s��0� <�2	.���(l�B��Kp����H0��Q(�W��:�:I��ӭێ!�3�J�{a�x��˚#�IȂ4����:�ç�`-S>l!Y��\�ABڒ��<��ȇ��q���]W��`SC���a�r���Lgi�w&�!Eޝ$ov��
�9[%7k��v~�'Zd��d`3zʍF��>T��9�H�qVd�$��׹�M�l3��\��P+ax��E�+��	m22�m�i8W��K����Y�U�ry��	C�����y�G�vg)���cy�F�Pz%��H9g��2W*���[8�9���@-���Y��Hb�!1��T�C�zk�ǉ�f ��V�����8�J�me�t�h*&`|����z��7dռ��Ľ��j�b ���?Er���ԅ�K�6!Ewg�#����9N�a����9=dۏ-�/����[�4���|j�2f5ƥ��I���)0��k'z&2�fA.��v����r���R���m3+�~L̫x'+�'�t=����}�O��˗n�5E��@m��0;k��O�����8�,}��ER���d�'�k<2\e�/��^|���=�:�C
��d�������S$M�Oamo)��`��sT(S^5���5,<��' �WUg�+��%߮OYO��Q�ݎo�u�<)}�?��W�s�6P{V<��4�O^SyV^¨��I����SB�#N8��w������QP]-�t{�B��������p`����H������3���/T�aB��/^��R��'� ��gL
�]HS��ipy�Ru�:����A������|W�y`�h0�H:�/z�7��sgoDq�H5,/�(���jM ޖk��ﺲ2��$m����12|�1K]2�3��x�+�N_��$����,,ª]���҆P�4�o�Ҹ�q�/�q%^�f�n�Eq�4�n���10նm��jX���$�����h�w��gKW��һ�ʕz�.w����Q-C2¨�P���v�@$��'5)*�WNgG���%�H�˹j��6ʪ��li!�W�M��� &(�->�V�*C����9¬��֏析X��Ѽ���lN8�Hb\�{w�6�,�|/��,&��z�[Í���ρ�b��S���6Y�r���)�_��JL�FP9hC�<n�^Wٞ�����ئ 
�x^��'�,3p"8,Z�R��H*/�`�(��s~���y�f���}���fl���/9���&m`8U��%η�T|�%�i�� ���BҼ�V�L#�[=�!����F7���puq���[pg$����?&��P�,�<:���/V����ZI�CV$��(m���R���������2���ؓlӅ�*�MD��zOދ���[� �93z�� I"���ATxS���s���H	ȘR�j<�-��dS�s1�����A��Y!_�� �Un5!�fH9f'h�f�f~z|�J����}O*)n�
� S<V��<o�p\*��Z�FÛ������*���:��� ���D.�|�Y�*s[�������՗�DM�-��?H���<8���fb����'M9����^Y�(�t�f~o�+��t�rb
xtj���~��5b�=)
�u���'�1p� �I^�X��⇱�1�6�����6��|B1��}fV+��f�^����]ӡ���ܹ�Wi^�I����k��!�1#��2�ύxB���Yʺv�K�b��!� ����Wh��u~�lgy�d��p��1߹(���/���?�W��5��d��B\�2iKU�z�3������0�[��MV��\�z!�õ_�����q�����"�����X�'f�%����
Ru�C�_�6�~XA����^�̅� ��������T珏/4X>�0j�i�ۓs���r��;1Cg"���+s�PgB1˟q٣��)9�J+�M�k�k�~֣���� ����)��*�Xrkų9���<�>��#���
���}HB�6X��ۃ����~��\�!y̍�+@�����x9�[+�,�:!��c&�Uli�Z+�m��ڪ���Ks���	��(���s#�J/I�z���43�
��颃�0ކ�LJN�,*}�����Ϋ�!i;�m�9�GB;�g_|=j8D��_�{���\����wd���b���	�1���IH�۳X[ݰ�Q�H���]~.�?���s:�B9�15�Zx��F=S���O�"���m%Dh�@b���b�ꕶ٩B����t-9��-_��7|46<�"'�t����,8��=�[z9KМX�w��r^d�^W�V��6L+�����K����B&�6�y=])���ne��I!#��ڣЩ	�~
ȝ���Oɛ�V��ԕ��K>kQz�&�X����8�09������P-��U��e�9�� Q��ϻ���43_�JuZ��)! ����f9?/��*�l<M;���W���Ovʞ�~ݍ�:Y��
:�Ķbǻc%!�D+�P���ҹ�&j�����<eEN�=��u.F�A=�z/=���kt��:���>�^�'�ڞ�|��O��wn�h�(ʍ7Z
�=?;G�g�]�F�#Z�$83��e6�#�n��x���R�i!�1U�_�3��uB�����@F�R⪨6��_�����#�xՉ0i�;�& ^�q��J�K�F����jR�N�H#������ύK��P�Ӳ��cu���Q����r��|��M�Ua}�Q�sO,a�ɖ�B#��^�U�F$=���@L�WC��[�P�k)����f���x���i��&��^˟�P��{=9NDX�b ����)R��qh&�T����**��n=�W�#�Di�ۼ�@�_��*u���P����a}�Ǡ����%���0`r���<ds�BD�i��An�G'����;�f�k�����G[��-':6�l���P��q��ۊ%�9�1�ȫ��\�^�(�A��JyQ4��(q[�.��{��h���ܩm��2�6��Ps[�x��]�OD}O��(��m6m*�R�h2�w�M��^�
�dh��������~,JY��{w�^Dw�A�{@�0X1\�P'�� 5IH(���������l��k�T���%��3��Bfa�U����RT�m����LHz���K�[J��Ugd� ����}�Hڑ3�|��ߏ}IWf�z"�������%e����8��bT��j�^YVF��p��7�dQ��/X�NS<��1E�Ȍ��[��"�
��~�Ԁ�P�݀Kaz�JK2b�j���xr�?�s.y\�f�o?_+bOl��m���x�J�_F	U�=/�Oxm	8?Y3C��|�61������`�s'=��~��K�j�?�i��z��|7) 1���xO��Ħ�!Q_��3�1ݏů� zG���O� �b�]���[��6_���0~w�&й&4��)~����5+Tx��Փǖ8�h<���G�woT�?#iM�J~QV�UU�-����^4�~��j�%�f~�K���8�ͼ�/[��*rNIu�ؿ���A	��Էm�?��J%�3�2���^��?�,�H��������x\�͠�PoҨ��H%e�[_���t;�<ߡ�d0Mp��)�6��������o�Eq�~kWB
���k���7���0�v)�{|�� ���]8<p��jN2;~ŀ�|܄^��"VȟMZ�3'F3l�UC!Up���,Y��`���
8U"zM0ò/C��*�/�Nxc�N�R(��}��W�2lK��FqQ�
��v��Ѳ��$����U�|>"1şہ-S-���m�g.���S�nq��(mo��%S�=���폪��H2�6vi�}�2���U'����5l@�g��Wqv�{�m�4�/f$p[��pu��H�ᬯ~ƛDh����Q��P��T�ȫ�1�5�Z��2 ]8$�f����f��pWB�A�tT�	�F�t`��t>*����8S���3Q }���Wu&P5l�����S*.;�D$�F���=Q��Y��!G���~xz�ª�7��?�(��}S�!��
l>�K/o�A����ܕ�H� ��\���&�'z���>��-d��nlH?,��R�������iU� �5���8�Sd, $~�r3���9}�-�:.l�S�L���fY�MK�H)k���#_ T���:�g�s9�1�(�R��?�\��^'�⎤����e��3Lr|�1�I	�￁51X3��u���.��5�I2mcp��	9L",��n�#ǉ&�c:���"̉,6�q#��nSժw�j��K���2�oV���Y�����)�`\�O�Z���6�>�j�T��X����q=��O�qʭ��2���<eS�����G�][��_�*�Z�}�D�\�D5���MhG N;�JL�U3V_����E�����t5��g舷=�M�o����p�DŲA� m�g:��g6l�j�����P�m�8DqL���)w"Bz�Zx7����^s�hL�H�oͷ�(Y�{��P�5�(��̈́���WŐ!��5�E�i��/ʼ��`�ceK�U#�Tڒ��C�'�)�O����	j3�����F�A�˛R�!~6�����>m}��W��Tl�+b;<��>������/A�c�w6�
��Lw��vK]4�Ob; �ޡ<��ַ����ٱ*�.m78J�f�1�x*�%/��z~/G�z�0z�E¶�`k�(�]��@�B�9<��[��+��͵A)�S+$�%�k��Ms:��/�y��C��h��)&���I�55��|TS�a`�-�w��%�+�]6j��Y������I�loB��n,[*ѹ8���g[8�j��{��e( dPQCJ/@9'�8�U�u��]J�$��\u�s��t|CT�y��'+�,S���̦��5�u����9F��6,A7�˻�g�'�����m	���k��?3Zz�x�3ñ#�DU�tYA�g���Ny�"�U����Q-�������[;,��:~����7 �f����Y�8��1`r�܅k��T@*�*�|��v˘_�����)���"��V�:m�q��6�+�E�sw��gV��3օ#^sm_2����2*ҿ�����Gk>�4��߫����D�����-�!�]@y٨�����;ג6\_���h2<R<�"
wr���$����7s���Q���d�D8��f������k�v&$����D��w��U�{lv[��*"�K��ls��EP�H������,
K��X4(��t�\ڂ��{g2yé�p9Q�m�����^����oFLI|�����S�T���{z�5�;�Ϯ�$��u��󭮸Bϧ=�8��:N���T��������W5}�;0������Q-Y�>�9S�M�y�c�;0��/s�;Ĳ
�F?>��/�\^x����;��g����\�� ��gV�J&���ǆ�*������ܢb��h(Z��O��ɞ��D�l��Ǖ���L~���r��ȵ3hQş{�hĈxx�2���0��� ���_�6�����T*�������q��G $9N�T�������y�X7� d��S�d�oT�h THA��)�Nf�2���vW+
7\oy�����3 �<8�h�1��뿇p3{i%�>)�8@�1LL��b�x���H�<N���RT )7$9#Z��G:i����ŀ��WO�{��|���2�Q��/c�����nc�.��r�q5�+��e����������v+R�!�+`�ހσ�A��Eۓq��l�	��q
H�{�!��dN^����:�mK��Vb�	u�vI���ц���>U��G��)��x����$��Gy�ԍ+D�nh�c�SCt�Z��Q���n���}�]�H�:�ȱZ��?n��,�`b:���a��~`F��sC1���T8ќ5�^뢱yN�A�.޻Ý�r㿘ʷ]��~�G����3�3w�ΔDZ�T$ׅ`���0�DgAg#U�7�+��m�e��t�I�(����3��u7&�$���Z�;/o(�������7�K����O"�K������$<GV?��W�@�9:�G��
� [ N��R��S���G_�Q}��7^�Tc�����݄7!ҏJ��_�Z2�:5oF@y���x�t��R߬�h�h/j_*�k��t�y),����ܘں����4y����X[����ͷ;���y�
=M��7�eyg��xg�&��^#c����N��~*����
�*���*9�F��7$(�8���#�,9�zp�}E��43�E�$J	�S��TЎVn�AE�O�k>�W�EY�cV>)�����ȇn�D��j�s�OlkR�E�;�γ�`����\r-?.�^B�n����4��I+�.g��	���߾�d#��
E���g���WE[���z��kv����-(ȋh8 ���V�c�?��2�]�3^�J�@�.u���Z�sS=�=�@&�f�A� �o�n�u�2TJ}��I�/�_��f���;����:K�jK�P	����p��ɰ�y���]Q��� �������M��ҫa���7<��*�j" a] p�?4�����P)~��'l�>��^3�j�^���iA������`��W,e�B_X�x( �Wf���لk�&/q2QI)D�T!��Њ�u������)��l�B�y�����N��^��fz"�(���l@K�UI�F/у1#�<�2Q0D�ѧ?�B�b�z�ى�\�n�m�7[�-�&b����M��+�*���2J�Xf��h�0S��a���3�Wl3��B|�Y��z�`���+���j�ַ����I\�苙�q�F��Zr6�jBT�[(�	�˱2б�w��&�Z6�"^)%��bX��%��'�ie��7����Z�S��S����=�vo����@*f�w#��> ���M�B@BdQ�q��&:-���}�]�\Nx%�k�YEs���i{V*�?�g�l�|��Z+T����xH]��8]��+�kx~ɗ�l}r���R=�<��=L���PP�aU����Nk&L��w�-�Ҳ'yn�[K&��|�+��0d���6¹���d/��ʪ��Jo'wk�k��q�ˊv�}i�Sת��|����5?'Ym�+�N��[�{.�^�Lp�nk�N�����@�0���l��<�~x`� �wY϶��� ��lBTV��4�u9GZ������,%�%pGzP�1�[h�ix� �.W��	�E��$Z�Bt����\E(~��#��
�ui7Er�MWlRP3��������fX��,�����GGxb�v��`WUa)̩9��T�_a���8��O��;6�V�xE�z�ݼ��W���By�y�B����i��:6�')�b��GD���+OK9��a<�Ї�5����l�Z<+���2��ಂ����E{~`Z��	�ՆC�x���*uo��x"e?%d�7��P���h#
J&}<�7���7g��T@��uڝ��H8�xE�ۙ,�����h���.MՅ7" R&~�y2OU �vo��
��Fo0�z�Z@_�^="�i}ѹ��tЉ��#�� �����M9��	8ǀ��& 2����O�KE
)���GY��w��%���).i�}J�aZ�Wu��pU`��Fsǩ�]N��~����C�"��43�Y����޽V[���zp�,B:��[s�Kb�T�!�V�O�U-�wh�|�.%$�ŤH�֥��2t���,0�H�h��x"�L��\�U,�T&|�m�+����zZ�e�:/��lfL��[�X��YG�}�WK�7�K6s��������s�0�	F�J�n. ��KƁ��Y?��Sy���Ca���fhP�8FePV�1��~7����c�z�2�-u�hE]�l��EH�m@�Ȕ�Ф�Q&3�E�� �గfH���^E~f��'1�bHG���t�R�Px7 �&�����RK��k�؃���#��2�����M
|L��)ϝܒ�LY�֎*w���wOV�:!����&N8?[��fn������r�uW�z�k����8U�y����'?EW��!��ӓ�V8�V�#��D/�W���6ޤ���D.w`�٢�>nW���k�h2g�8�,_�ôv}�a�F"�� /}��̢�&i�|�P0:A��ae�p{Ԗ�ʼA��m	s�ma�v��c��������IL������G�N��ت��ɸ�P���>�=PC�X��C!��_]�	�o4���m�������P��1�b/���=C��htx�4�ք]�=�m7�e�1�Z��&mI�����8�o?�!�j|������l'��T����<
~N�>�Ή�7V+��$�	������E�k��?^�#��HpyT�r����l�1��8v��>���K:h���j*����Y�d/��~�ف��R��;�m#_.Bvn��� �����bʙ(2�T�0Q)s1{FA�pR�6W�-q# SW����$X?zUT:��Ӓ(��Ԡ`D^�����!�C\�dbv���}ʄ���V�e�-���k���_��c�@l.?���[�|-�@U���5��@�F����_3�ҩ�۴η�E{���s�?%��৚����w�E*�������3��Qb[�b�A7k�5����.�S���#7��c�umeY�����i/g�E����z��E�F�:^�=�p��56�M¿lrYʼ���+�y���u(�5�hW�{���'Qfu�f�'��v�%����2$�͏�'o~���g�Č��{ㆣ���7{�^��$��x�<4��58
�J������#�;ά�����.}t�n�
�mo�Ԛ�ޜ�6`D�0��e7Vv��=�ӂ��Gʦ^������թ�D+���P�M�bc�L���[k���Y�ԝ;%\>�9s6�D3E��Q2���h�n�~���L�+��
�=y�������+o�}~mO5��v��f"2jZJ���ң�t�v�wl�8ΏPSկ��8�� |~���IC�G�i���IDr��B�&e����$�D_���Fg)�����¸&
jT�K{�>�����O�
3��S��saI�|wG���ǐO��J^��K>��(��`߈��}S#�Xce��/���_Y���YO�Y�"��
���e�Ɉ�����-��J�s���:5��԰�f�^���i\NT�6��Z�b�(���x�����L��FPʴn4ڰ�A�Q�8����%�m:)�����ه�:L_үb���.���#bwBx"Tp��K>�WW�*<�P��$+���T>hH8�'f��x�t��Dh�C=\dE���}*a3�����]�R#�y�!��3����)'Ai%$~l�xv�Q��B꾲v�.�..1r�Q�@pԀ���ѝ�V��/T˧�l2�ҡC��s�3ABM��A����]S¸6P�O�a��X����.U�E��YN*LaL�%2\̩�Oe�φ@D����Ƌ�u]��T�F�*�f0P� rM�bȍӰ�|�NP����j��6���Wc=+4��]Ԙ��~@��5�$��wmg�I(��yGu�c�4}�_��E�5��v���q�U^�ݵ:��2��#DR��!A��v�g��[T|B�SA�j�Rp�?:*cړ>w�R'�6��*J�"W�QI����97�Ǐ<�X��dx�����M^���;� ��6}�B�Y&�4�	�4
�@!HW�﷘щ��x��R��2{�����x��:\"\i�Qn}
3T�y�{V���.��b��jL�L7�r�����P��*ai�: ���٩�F���)D塕����Iy�����}#�J	^�ћ{u8:�45���^ ��H��=) d�F<�,��0VH7Ϯ% O
??a���&��J����nO�A{��0�?����߲	�4=D��]y�����wg,�gO��^�G֊0�9� �q�Y�h�����/ʓ���-:@�K%)��rܞ�A�;P���1�/Ұ,�z�k�y�C�*�flܒ��mG�i�j��A��4���!jv��0r��.�Y�_�k/k;��7(��Z�
8�]<Ȟc����l���go���^�0t=ϛ���<��.� `��a�Z�Lq��u�4&u�S��+TUVGgK��n�\jC�奸Us ���)�����қ��pG���d�GgVdHh�O(wj
"�~�;1�8���y��r�f� jG��F*�4����?��?�����ue�I��B��^�h��6k�7I����N����]�i�]S޵%�v�{��#s�7'܂��gʢ�m"5����Ϙ
�hK��{ą �>6p���Y]��p�09�N(�:�1�X�@a�/����o��[���X���aqr�����%	�wG�A�l�dY߷9���N��y�Os�����y'����_U�0C��$6"a��Sz��J�N�H
�`�nP���vm~|(��/��U!�h���Db@�S��߷�pSx�BMa�?3|
�-�F����SSsQ��*)�qhTX3�[��#�hs�)
,m��P���*p���b�pw����d`�M�x�>6���e�����% ����o�D�V�<l�{�_��jj8�%l����� ���N�y�~^�k���bM�<�w#O7����\�)��7@��b�$;����3�2v�ݮ�s�Ο���ۍM{������~(r2�6�>�LjI�)�п҃Gx�v�c>�(eJ�I�6�)zb\?nQ��5�ԯ~�K�D�Eb<�v�)���f
1�E�ZV���q���ho7�l5�;�2,J~�|'W��e�̲��B?'��"����H�[��
���������x���O1�q��E((�_y��5Zd0��g8�{	.�N��
s��ܫ��o�j�<o}��},5[��&v�ʒ�hi:�	�n�4A��`�ߴ���vi��(�a�YChh���a�]ݸ6�����|�3������B���9���B%�b��Y��uU�3���Ή�/{d�&���WGïsxe��d�Jh�l2O��M�|#T\-؈!�P�WǊ�}%>��h�AaM�B���-�iM�m�Cސ���dOH��v��`e��en�WW<U����bdc`�6��D:K���F��X��43y�@�ӚOrcoO��Ps7,�uxX�ջ�n�D(N!W�7WHLX$���u+����M��ڌ%���Mo��SPzc8��B���ԁzQ����^-�	�)��4����L�rFX'�0����4)���{�߰�p��R:�(7�U� �&�p8�3��і��G�X*��v`&z�m��7�4 o]�����`49�w��#'*��Y��
��1�q�j��,���gsS�i�4:��^���?	���ŧ��������ӽ�edwP;E���Di@n��Y?�_�'Ĕ_�nц�Y�A���4*b�>̤AŦ
[l�;dm_��V9J[G�ݓ�uIEh��cM]�=ə�û/z���KD^z�^I9�����V�k4"��S\�� ��>�����z���ו	۸���41���:�s�1iP�|�6���~���C4��Х���G5�q���7-Mr�a�8D��h5�ۼS��B��'��J�d���&v��,w�D@�͔�Ylt|��%ۓ�S��3j�N5���N�M)�as���^��3ѧ{ J��ws�}I8ma[��}���C�'𲝭sB�Da�K���+d�k?�r����^�FA�ە�J��RgE�<�Y��h�w�E�h��r�sb���*�y�kO�<���v/am��� �ө�j��lH�c^"�_��ԬvxL���s&���-�5fY�8��a�u\��~�)��犯×��e��ɧ�+�5�y>$1��s���h&��Ŷ`�yw
�vϚ_l^�ۊJ�1-�SԌJKBi/X*�~�/�.��+�M׷@z�E2$����]���<0Ӫ& DK��ҳA�&
��M�h4	r���?F'�(c33�����[#2:�y����?wE����_�	x��|N���Q{�0�m����~^�I@)"���%mU���R�����o���p�>5���x��~���oI�Jq!e���=��BH����T[������K� srPN�g5t3�٭�{J��o(rO����&)���P���UoOO�$�p!b��'�\���y�-w�����ҦWT�O���l�Wߤ�b���Ts("ޙ*k�UbZ~��sC>�2��
R�B����2��#��*��(h�&�r���T��7dq)�R߷�Δ}h9s �E���n�ո�ٷo��X�Z�[1�U��q�ظ왴.'t)�~�8��KԾ�{L~�djM���*v�}3�\~�F0E�D�0�+&$����{��L��Y#���n��C<�҃�3�M����g��A�3���\���l��"�%gt#&c����Aɗ�3��0-o@�Eܶs7i�9Z"����L_�7�����
H�MD���1�j'e��9i�:�mҰ͜��ρƦ�� ���?�g���,�	����
ٴ��T����B�v��v� �Q���v�`�!_�$a���\�Q��?���,k�,��Z
&"%���*�����!��!���	���ޖ�A�B��FT��:V�L��Ry򪸓+C�Y�w��
����F��-��в8��籀ћ(�fU�^5�i��[�V��/j)#�N������w�q���e+�e�^j�F�5ȦY�E�&M@؉�K�-�tu��H���u⦋�z̧e_��FF"��1:^R �!�j'�D��o�ب?����W���;Y���{�9�%��:�z����6�!��$'p�����v�s Yb�xD�.pl� x�[��K�,d7��C�iXj0���+�?XIT-��#%?������#�?,+�N�?<��նcb�2�8�F��5ŵ�v��-�~&U(���t)���r|$�׻�;�k�w���\mQ�8��fcH$���
d]��No;�Q;vx0ք��ǩ�DL#�|؊+Y�ǿ�(�㭬Dp���m@d������y��gJ��!r$�N�F��aI2h!j���+{>:[���o����<X}�D��y8+���P�D�l��z�R\�pB�n���RW���T��{g2�;$���^�2�����L�;���CUA�(j�a��E��j��gb�G"&Q�5�ڔ��@�l�1�6�&$�#uɮIL)J��"0�ƚ�P�0-i{P�h�@�{��-��@b	S�&7����;rM^��5�Cƥ��L�B�/��h48�j�XPy��Ô	(2��W8#��1����d9�@`�?��Z&�%������	v����db�U=��J �g��Џ匉:�[ӡ6COw{�� +j�&�D�s,A�k߰-f7u�7��q�ң	���~nĕ���oY!W�.."^�ነ� ��X��-2�)����َ���/f+t���X��
O�o .����g�.�V�0�'��=:v2�Ҧ�:��@ l��3�+gV�J�J�QH�O�xU`領�	�sp���S�S�+������&.��M�c�>(�w+%�G��&���ij�����~�IeVd��4{zo�{�C�[�^��������Xg�����'Y�\�sʑOîr��L�>��[3����1 '���c��ށ���.k�G�:=��q�M.2E1����曲6��q'�`�v"�Q������R���[�a��
oo�2�K�v���	6���֋�����0��Χt��+.O7��<���"�"ʬ�<^��$�"�c.�=�($��qM좓�ya�;����c�����������언ː]U�v���f�e�Պ���O���6�&S #�8��;Um�E�������Às�	K������O���q�m-����Y��4:��G���=�EjH�n[E�Ҟ~�̔S!����Ⱥ�5���Ԧ�D���BѮӶ�#��_��T��%{j����NY���^όa�,Gt`"���P�v�atI�*�(�����(��^nև|���ד`�vh�%���5T�OT���Xc7��N
q�ܝ�U4뷩k(y��e0�d���%�?��n�rnGh��u�QŒ_6��:�P�s�D@�����?���j�>>S�K���"�V(�ם�_>2�9�N��q�
������Kh��DlCg|�Kk�r#��R���C���.;g�PaF'0��t��3���p�\�a����{\���9��n�!m�� C�>Ad�Lvh���<��'�Q.@H�c�UvG�=���wPH���T�M���N�c�FwA�U�^�u��o���/�"�H ���0��2N ���$Ζ,��nb�ge�t+;i(�?>��c�u!FO�:n��9�u1S�eu�b�jN֪5d��U���#@�L��ᇬx�+��6���np�*8���o���#��# �J���p:��#��.*M��Ec�:�h˱����af�%u�����Jm����F�_�(���W�zM�I��)��dDg�ݯ���G���%�׳}\��ي��Lf~'��d���9:ق�b)HH=��#����^Em��|���b�'��7r'(8���f5�}�֣��Z�+J[B�7 �/〃:������GùQ�v!�8A�r�o��OM�k"��k�Y�����rr��B��I6�]��#�ä�j`�#Q�n_Ɵm�ʒ�\�.`�8PW?�*��/���� c�
Q�!'�<<����)mmV�,7��}�x(��!����~� ������O	WƜ�Y�L0G6����bo��ol��J\B�оc�u��6|�����;��H��=Zߔ��)��k�8�rS�ɮ�)����-e����6"(t����6X�A���
P��-�($<�gL��ص����������Y��1�$|�w�*6K��ԿMB�?$,D\��
��^E+f8�(�H�4��W��@��U*?�4Z��}���M'H����»���J�|�����|wV9N����X:�]])r�/ӌ��gA��7�j�����a�P�[��a#��m������������b.�J���ܻ�������b��L�W�p0�r��.h�參�&��n�Pu/q.Th��+|�![�΀���T6�P�`��<��,��(?^�{����l����V!�G�mn	����P��I8`
�ru"3�ߧ���Av��s����	~/=���I+���r�I����67bƼ�޵���qL�s��%�*���Bo�{��L��]&z(՟*O4,�N�6Mw_��`�M�l1�g�2~ØH�RDF@Zٟ�b���rE������B��Nlto-ć9���ڕ!��`_:l<wܞSƐ����^��]�8u��+����s{{�/MfQ)\>k-�?ϯ�RC��k��m8g�u<�"P���Zڒ�q��7!VG�p����q�LW�yzS�
/5�63� �[v�NŰ{��r���(���� Y�w�����x����60�?F[Y ��X�,�^cζ�n����rԜ�}��Czí�l+�lp�.���w#c�c5�L	�I�����Ŕ[$ԋ�h �����|�+��I���1��j���(ƹ��lNՊ�|q��[�L�"�j'�\��������̃�5�ʄ.t�R�7ex&�b�E@��W��G�p�]%�bp&N���)C|[�yA�V-*�oH5q��;kiqV�\tK�d������C�Ya�� �>�tta��7L��0c��Α�{:!�ׂj�l�6P�@�d���b��
Oj�����o罳nspc��Hꅖv���)��I�I��UGE|xM��WbP6t���]`zo6D���␎{���#q���Э�i\���9avD�r�W��b�޶��]^@�8�g`;в��Y��,e��	�?�;���]��=���W���B��P jܸ�QZl�;[>���0�]Ac�]A�ױT	ؚ�T�û�/�8�le�M�o����ߥ���Rtq�0O|�L�԰��ϯW���~]J��6A���a]��VӒ�oL:g��!]_���b�����5��2��:������=�t�s-VX����"�(v�V�Bg=X�@��$[�s�gDJ�p���D�����i��&Ui��� �6^ Cp��:?jF���Ɖe��Gp]	J$s�O0�Ŵ�Z�>J2�ez�	��_@>����2��*#�2�[K>�5v� ����E����t9m�Di}0W��}d�,�)�G�L�D}��*��]#(�'MǱGY���.��֯��)#�yr�o��|��>�d�D���\*��A,���[xn���W>a2}�X�$+��T9M8-cB�ke�i��"�|�$���^��JT���3P�@K���}�B����N���>�W�_ʲh���L�"\�5�Ei�<�(��z��7(�DwN��Y�n�݊t|��< I��X:����.��[���Ӥ��)��HÑ�`��Խ�H0���q���#{�\�@u͘e3<6�X��6)!���=)06H�0�{k��0��y��_~�=��/�i���o��ur\+��Z'���X����:�:=���]}���ɝ-y�萗�ZP��a봨=�����f����Iw�bn�c��;E��Q�hPZ�@�m�J��������$��TD)&9�)�(
+ϋ*=���s>5�����<x[�o������ZK�"|�n~��ؓc����פ��@�vVY&� @}�3ҫ����︪J�w�NX�izK�ܪҚ?�ɚ���5v�e�5_9�b������2ꁲ����ۀ6��w�l�{�|� v�W�g���3�ܶƊ����TF�^h#�(��4���F���	��ŘP��q�����S++ښ��d��9��PX�4��Y@��k<'���tنC���J<-6�_����y[T�P����l��'�K�����5��/A&v-v_s���J$��!�@��\R$�h����`�W�qF.Ax}l��α�0WpǼo�8�����"�S:���a���i<���-��z�����T�#�(B|o�<!��,6S�~#��wgxrה�$��ߔ�!ЭXG-��y�fr9�a_��9�6I��#�c^Z����oE����c}$�|��d6��V���]�<=M��0oh�6y[�9�\�*�e�՞w���m"t���=��6��"�@ؒ�J9�/,i��cWm.��p�3UH��O�ǿL����Q�� j��ct��FZ�N`(T��k��S�eS���~�Ӌ��j�8Tđ+�G�}�:�`��Y���"��.�#��w�����[{4�TU��~�y\>�p��w��A��އ�����bݠ�;��K��z�#�!ƅ|8� I�>H�t׏�K�Q�`ɼ�-��mv�]'�%ʵR����z� �kßT�B��S��
�����e�Hb���_A���A|
V��_�Ɗ�
��!f��w�B/��,w(ͻዀ֥?�G\��G���f�?��5�rU�g�Hφ4Z�;��l'e&_�.N}M��*��@�I0t4r���`oO����������pr���N1�Gt�[tQ��@�Ů� ��˽6XIM��/�ԕ�g�{�9k%�����%�܈,8��P65U�Q�|��HD:$G�o�#w�����z ��:���6���2F<���q�5Fjc�~���u�Cչ��p(!��Tl���B�)�	��ɭ�<'������$����yw����<*`�:� o/%���4EY||Ey�c�`���o֒�f�q����rF���fM��Q���M4�dҨ��;E�+�)�2h�Y�R��2�r�e>r�V���g[�Ce)�ѷ6��0��Й�/_�7w���x/�:��y������j�kMH�l*���1`k\��;�	�r{8(�PB�(��}TR��'��;�;�L�Hٻ_��QNMr���
7@���Җ@&U�nڼ|O�*�A&x�����7�Kug��et���H�Rk���
�֫TO_	�\ұ�i�¼A]�T�,����[ǻ$`>Sa�z�L�����O�����(�n�P{�*�'�V���`��u�QG����O'YI� ��d�ڣ~�����5r鋮ȳ~5x�ިv�?1K��ԳQ�zl(�5$�t/�`_�?�r?�K��L�+<���'�D4��YU+"ɅI � D�����Ev+)(YVotZT2Y�ƣ���������.X�&�gĎ43!����m]mBX�~��m�!;{��,lY~�Z���"�5�d��7A{�šo��I��,��r/! ��.N8�̂���1�PȾJ���f��Q�H���y�>	�љ
�(�0|�� ���?�a
�F%za�k����Y@�����IPy|���T��=�hI�!c+|2�����"^&#c�*i��+�OYUj(�=_e��#��S�ϑw�nS�����Z[ X�"v�}���\ o{ ��*sV	�pn���:V+*є�kc�G��޻RƓ����/.�&��z�6lNsn|`�v��r0��*?���H+MJӳ����gb��"�hɔ+�����fO
1�yqi%B_7�̵�DA���A6� 'FoS�ZVJW
(�b���qJ���x$���弰\��Ꟶ
�:~���2{���t{�M�<��x^��������e+���7э���j/&��@���e|fЃ����
��X�H�s�l����/\{;:$�Z���$��2��Ug2�%��8��ȟ"�!E��Fپ	�F]�n2P�1�f�=�e��*�h�ga����`��+>n�}`��V������7Nv���'[{=�O�v'�ѺI�Ma��8�%�("��N�<p�饜Gs�Y���J���8�� R>��V��8@��]�����%+����{]:\ym�	�G��$<�iإh�uB����l7���d�T�=�1��*)����O�%�����?x�o��r�Vڒ��9Um��^C��~{3I��
J���%a̶�?B��Ez����� u���Ge��yE"[#��N/�*�Lt��r�^��Z�dV�1,F��boG���@�Ǝ��.f-�<�=<s4�,�]�٠g���zB�7@ �FH�DW�:��� ۃ{T��/��z�����uj�>��l1 �"֞/��(��IB��+jL�4g��hu���?�'�OSZ��a�X���T��ӹ���bc��,�"�E��6���';B�t�N@��L�~v&��`{�����y~̴���P�B��s��L�:���V����b�`��[����}~�e��}4R�iƱ?a��[)�o6��¸���'��KrN����l�L/L�D������u<cj� �/����&qjr'_x���*�����T*��ۦչ�m�MC\��+YDI��'U~jUH�Kl{�� e1�3�_U s�v�z]��'�M��� ,8�F0�ԟd5��VjBzS	��I���T����'�G��ې����D;I��5R��O��L^1- 6��)���VϕY����"�f+����d(� ~Y�|��m ��L-K?[V�踃Ƅ�N�XX�m�"]��հ��|�߆��I��tېK�X���v�A�Ml����QL��#a�_��vL	��g6|��g�4��7K�C��x@˨��b�������L��(!
�h�xq��
_Z�8�<r��(�q�=xk?�G3U'���/j��x�P����_���e��6�|ߡ�T�����=<\%�^�^Rhy���ӝ]���w
���L�<:D5���rF�Ü����+�Wi��[�#gU�S���}#%�ȧ0g65�I��$��yY	�������.��I�J/FI�.��&��W���<�^lZ��`�J���'cyŅ|$m��3V��hn,>�7���ŽM�`�J�=R֖���K
-~�e�i�Aޮ`�Z��Ѝ@8 <�Ǟ<��\T8���c����ʊ�^r�p�~�=��\�o��Y��\�~O�jF��"��N��h9r�Z�vT�+��n�����Ǽ�6����]�Xf���[��n���&�ee���Ng��9[r�wy�W7�d�溒��-$�="��T/�<��1H����B�"��#Ԋ�h�9'kӁ��½{B�ބw0�����C��ŀT�	B�i�z���`��x	�pd6i-������6�Cm���!Ԁ�y��y����J:��(�7[�d�?o�d�4Z>�����1�[W9/�:��� 
�N�{5T�p��i�R����\��[��+-��ORP?.���]��3�=����w|�ow9[�k�]L������<`5�+�j�����|}r�n�s�����L��R����	U���M�U4���(�C����.�;b�W��~�'�d��bk`�h���ַ��j[{�վ�pϗ�}���b��ß¶PEĲ>�E��Uw`�ʸ�0U���Z;���=Q4P|B�êDD#�eINH�?����,�cht��U@��4�0Ђ��}7��F%Ù�2�tJg�)pr�hVP^k���&��|��a2.�J��_\l���X�-j�P��C7�^���U?��mbT��kO�o��*��yu��\�nH�9_zL�e#��Ӧ�Ѳ'�x,��Cյ��u�=:�����Ь�ea|2�)&�J�)Ɲ�E������Ҿ�5�e:��F����nV�4����������!�O�;������W��wd����5�0 "/�1��b>����w\K7���:�E��W�u7o��W��5?����(!�+6S@���z_�y8� ,�T㾚R}��͘M6���Db���� :�k1J����)�̧�]�C�9��͉F7�ݸ�}��!�X�ܮ�Lq(o��h��� �]��}�abׇ��l<v/��_�{ �'2��7 ?Za U��-�2��H6���ӎa����1Ց'OM��`i�(a��O�V#�/�H�^�"��(+��J`7}�(o�aM8�P $�v8?t��h\�9��h����g������.��w�X=VS�G��s�`������fhtt �C�P�ϡ�o%�<e�5�oI�}��E���ҵ����ol2�!�o'/q��4�v&��x0�k��Vrc�#;+8�/��fy5�j��*�1��o"�y�:�Q�~W��w��rہ�#�*�]1W��fi
���;�����OE�O��(qH�U�C��O>�^X���o�R��� �RR<�!�E�@�;į-�^�MD�������&\��6��[u��� u���I˂�;����UEA銛 b����s�� ��������nQRi��7U�q|��Z=�]���	Ɂ�I4����N�y���f�uJ>���Җ�z�ș��F��v/f<7e4�*�t�̀5�)4�AW�� ����G��Ee�y�iA��^�-=8ܧ7�'��! �o�DwjB�����4f\�٤^M�Ϯ~�a��l8ξ���Ol�ol 2nWY}W��3=�6��A',�����ji���N�ӎ�΄��qd���ᖯ��>�	���E�!�r�Q[�M4o��P��Eu6-r�U���Ԁ��c���?���l&�%�=$f����D�� �ݭ5��d���F�&�_�ۊ��b� �&��z���ng$��.��:������P�*@��<#�TA`�*,9�i檰��n���G&��帴�{�D�֑j�*:HK��\���F
KlCHrX�3�߭:CE��6q�Ǡ�v�q�ap`"PǗ꒎-F�	�B�l��m$�.[�~���p)��*y��R��T�:���Ae�ȗ�{\�'�O�ۻ�)#աѽޘ���ⱸ�ʐ�
��3�#���Hc�.@";Ҵ�g�t�`4o�v
M�0bʯ���R��^lԅ����M�����W�c�`�ʹ��ӌ8�ĥ�>9l.�4������'�ty����{�,	B
��R�(-[��21�j�V��ث��f'��v�rD^5a����~��j�~"��i��%Ô5�3��y�o��I&��W�p+=�Y�%zI�����1��Ii�A�4�������wy��v0p��S��O{��Gv��"	E7���h�KV�i a�Az{=�P�@��[w�yp�.���z)��p�u�y�ƞ�����M��iϮ��#<㔂4�������������ԓ�􇱺E�r
�b����c�eV�'8�:�*��+UL��EBS�)�T�ۆ��"#����݉�"xy�sa����EL��Mշ��13]c�� g��75��)f��.�y��Rj�fEn��E	��+{T�`�ID�W�FF�iO ���gH ��u�d�L�~���.��#+)^�J��,��D���wp~�`0jx��8�L��4�^������<�m���s��f+B�0���Z{k���^%jl��î�����z�6ӟ[�
өG]�]�~&�Z|M�n����KG�J0��:,���Kl���3^�����O�n��D9Zi�:p��b�˧�Y��ιqhP3���a� [7�\0V�Y��_J�u�D��ˢf��:R	�zm�8�Ĕz� �7܇H�:�,by �v+�n��$|"8䴬����1�D(���L@�J6��@z�ƹX`d�C��c�Xh'p��g������yOȶ����)�&�=b���Z��p\�1���H6m�T��z?���o0)��I��������;� �������ɦ��O'���-�իG.?E@4mXά@Z�r^f;&�����5�-����-P�P�dFVp�Vݕ��Ox��v/�OB͝~m����'���о�b&�>�5N��9D;(v��B���:��UgU\B�4wO%�P��Ӻ�2,K��w^��ǎ|l q�����Tg��luwF��j�ʞ�1�j�1�K�B��˲�H�l �)ąF�2$������ U���O�g��Z�V����@�[�5�!� ���f��%7�C�������Ŗ`�Q�3*�}�k��dek���l�ğ�t4՛�m�c/#��UĻ�\?{�A�f���\�%�1oe��� |���o�G��*���6�����d��Q����)��7��}�̂>�%+���l�����J	y�7��?�
�O�?h�!�CGI��=]�lۖU������Y��_��4�xa&T��kӔ[RfdN`�J���I��$��N_�F�k0FS椄j�-�c�l3t��i��3����m��K*n,Z`������w�{B8}�
]�L��6�W���U?��4����4�2�*2}_ ���Qk>³���*	KGİ��ɴg��|h�A�b�䁵x��;��K���uH�����Q�ꑢ�֚G��n�L� s��}�;3Zv����.T��*٦��C,�t��^�����D�
A ��F�i�Y	�I"�E[��KH���C俣��d�e	xY!�[��o ,�#`�ˠ�^eR����6Z� ?bɲ�Ӎ�[0�	a����mWL��4Ro�K9g�)�sN\U�H���k<��m��4�>�7bK8��`�l��H}�����lh�8���H�-�m�� �LW��7����2|��鞀3����M��7�ܷ�LuX_*鵤xœe<�n�b�pp���ܮ��{��疴��Ŵ;��QI��xu��ҭl��!*��Eofj�ej��l¨��:� ��P�2�^/�қ���I�����a���1,�ѻ]�����;����p������$Vq.���@�3�2T���/N����zF��z7w36�fEa^'/���І����ȿ���0a���6��-!ӓ�qO;K	��UPٕ �1��Vؖ��[|�-=�S��&'�bH�tu���fB������_�JCS	o,6{nnV�=�z�=nȋ̃F�����Y�"�!-0f��Xjb�J�<�޽BK[��lOZ�����V҂.;CA�$�C�@©��Z�V�s�4b��
�`i�.D��gR��
�O��?�Pu*��W\�)�<��k��p��ߢ)C�K�vt�@�����鶏�Q��M<�.ɀ�S�ڟ>��TU�Ag��E��R�J�sR�"x)�%�Sd�W��B?]{7�\�
�@"^���ojllEf� �$����R�ÉU�89�V�Ddt��äy��#w�k���t�W�����-�G��6�WɊ_�G3���SK(G�Q�.��:��� ^�>~ �6ي��I/��/޼���F�M�2��q�����=Z
�4N�N�	�����]�)�/���uT\�k�M��˳��񖚐D�9kTbK���������DK>��~�?$�7�H�'��*�s�����qT8��N\驚2�_S�-�R��[�Q(���_E�7m����VΜ2w�]`�]:!�mvͤcr��6̀}=I�XRໜ?�0���=QԆ��Å�j2�o����K�M8����h�����M�6�B�Z~c����Y�M��q�M���w��q�,�/呎�wW�=U��%|��`[�FQ472�>Q�����zRFъ��S��)5�l�={k���-��:|'}8��i&XA��$��B�C~��)���<ra�4�W���!
A�k�(����͓��Lل�B��i�*Y����j*��Y�@	�xknM_� �u�� L����R�m�r�Xʕ֡�ed�8O��=��F����kJ�Zf�4c�֚�������`%rne&@X��e���ĸ+O��>� ��T�[�昳s���#��'U�5��Z&ȧ��,�-���K���x]uc�?A���?�jynvAV��1��)�;9�@NlS���7�GEN��)s3y��c�ޤ���Y���df��%g���,�6캇������ՙW��	eVŵ�RA�&A��Th����D���$˥g�E��N�(����@��\D)Xl��uXppMRѡK��͙��t`���*��y�$D@k��ġ��R-���l�2ʞ
΃��& ���n��q$X�Nc4���Y��wR�KJ�k�
���jORE����{���77Ab��ټ>{�[Ŵ�-�4RZ�n'�� �>�?/�Ȏ�	J��d2;�s�PϏz�5<��k�ᦈ�>�u:�J��)�w�wwΊ(��B��Bo t(f�W̗g{A�S���E��,̣c�-��9gA(���IXL�dBr�l1[�����hͷ���=sE�GJ}e1#���X�`=�SDB3�F�^Pl����'�o�(<)R��/�M����{Ԍ�5��عmӠ���D
��ʺ��%Ds]s�qX8�$b��BKB&V���y��"�Ht7�0�l�� �If��`�>:�l!O�@�mi�f�8Ō�M Y��8
���@}��g�v1��9�P���!E���#a%7]x�VzskP7R+��{��ʪ���5�9'~.�;O�orw��y�VP;%wJ*�����E�f�]ߌ �:IP�R|rg{D�;T� Åe�?9	ҒJ��T8���^�0Ul��~�d5:M��nR�������2�"�H?��>2�*`�0,!D�?�p�&�Qh��\Ii��(r��h�Ea<!��q��2;���Nޞ_J~{����������X	��E�h>LKI���X9*�۔*b��Z:����{���'_��5�����a�0+������豵Z,X�ԁ���쐝0�(W��g�M�c��&�#ۧ�55I�X uʦ�/�QS���Dd+Zhx�;��ÔUU�8���X�#:(S��O�;Pg�[T�w?�����T�����I����������UnZUO-?�{�q����o�_�ۏ�a
r[�z����n��*�T��(.���x �I���O!�W���'V8$xS��Oyi�	��U����̂%�~
Op2��.$�Xg�,O��AG-��^�|�<���"�y�W�����x���������+]B7�b@t�3e/1��
�I�
?1���ؘ���~���rE�S0���L�/UsN�Vs l@�X�bd~�����U&��Y}F��pL5��T�v3�4Sٔ���gf����ڧ���$ $��:�U��G#d���|`��̐=N�\�؛���)s�� �a�����g ����k��[�}�RU� j@�����g���x����*l
���~��3�[P�X/-=FD�U2ڷ�~�$��A�`h�	��+������֪Hk���ě{���Y)���0�����ח)����0$oI�
Ҡ��v����{���3Z�*lC�f3���ӳ:TO�#}ғ>�\Wn�~2�
ʃ��+AY��
[CyN�zz�\�Z!'��=�cP�6K]5�gB|�h��ؽ�3R{	2�O���(���8X�����Q|�hL�se��!7�mX[��ą�~,�ԌK:�\�匈oQl�}X�����*� J�"�����@���}�N��\ۜ�U�L��!K��7�?���]��LOE��H����]<��r9����i�=�mj�@;Z�`,�P��k�#&*P���O$S�a~�e�v����Ɖ�	��r��N��w���	�)��-.#t"�����/uc`���w����^:��UvHC]�!ĸH�>{m�ֶ�f�Q&�$r6:M���,�~�T��U^�/���r�Lm����]pG,�.Bl�'��D�����M�����%VzTqLH�6b��&�&��;8$֞bC�������㓣�
,B�m=�-����f������������e�1�_.���U�P�φ��U�eS�і���GGC�%v�k�A��FN�Ga��8��®�b��5;2WЂ���tn�}���k�YzE��ɺH��H8���^�,[=��lv�6�7��/�!anG�O�2�Q��re�EZ��YZiJ�)e���gZ�A�< Tΰ�^bne,���5�ka��b_v��d�V���0 �X����F���)S'���n�c��<>O�J�Q�+6����6�q��I8@���VaZ�iET��J(7�5\	!R���l����hs��7�3��w���a$�C���^��5~�o��Ʃp�Y�tT%Λ$n�V��{����������<p�����)���n�j�TOQ	N�U!�-F�뻃�F�&Zf�gw�fo��K���p	U�4=H�t��y�����fZ�{�Iqw�#"��d�X��אָ�1��n>�gi��ʭz�<���jZA�k>���j�S��_Aϣ
Iͽ�����p!�Gn����N�d��*#xIno�|��~fJ�ڿ�P`���LX���1���{戼cX��v<�$$n���CՓ�yͶC:L��K�[�-i���"�Dl����ᐽ����'�M� ����x/��ߡm�H�y/X�F�_8�i���O���Lv5k�jA�ǐ�")B�O�s�����c�G]�៓U� 7��?S��3s�
��ҽwPE`Ƴ��z|B���N��]3�����^nBFZM\uB�h�9�p��lZz�5 ��}���4yDq�f=6G����eǱ��	��~�ݏl����5�-2'V��@C�r�c[�����ЙiO4ꈂ��o���J�V�Nַ�=e(Y2R�{5�3E��f���Q���{�""v���j�K%��:\BG�s4���yN:�>�E�� ��l�Eb^f 5�R��V՝�b��9<ko8.�5%e8:�*�z<ϴI�w�HKo�[�#��(����1�Y�~%�MXM��b	�Q�_�ީԡ�uR�XVז^hI�=�"7)'M-tYd�����5�q�Ԕ��`|�xF7z&Xh.��Y2X������m�`v�!�����10S$��(���|����A���}J�cb&��{��P4��&KO�:ս&���a�
� �.�Ok���ȯF��I*U.��x����vD�W��i��}��g]Y ~����_��[
_��Z4�]6��"/��嫧L�&|ɐ:i]L���̭HQ��о���"�����0�M�̓��Ā{+s�"�9>�^��¯��Y���+\��:�#�Z�p1��zS���&M�.τכ�a��P���2�cIE뺖�U��7����0p��U�q�c���!�����Ye�����h�}N[�'�Q}v�*,��PTo�4͛g��k~��Hb����@fj槁��Ļ�|]x8j2�snrV+c�ˠ�\B-�IE��Mu ��"!kc�2����<�ڝfmA��������p�獴��(��Ur	��VO*S����v�����<��������+���	�#��f=������&�3���w�c�������ܵ�T˱aiG�4StH̼������t���s�P3�~�샧�������^'[V��,�|UB��]F�#�*�n���������q�pU�z�i��IK,̓\��$e���'�ܞ�-�ŭ{�eZR����p�A�0��?锇�S�0�n�;��P�Y���N�?gq����Q���巗Z��(m	|����!���#����[�h��Ԉ����\���	/ޜ������Mo�`l�*:4�-95;�ͯ$�$)�D��Ohaz�ḷ{e����z7q;��2�"���l��y��@v�gi��2.Y�)�-@�=�03�DJ�����з�����s��Z�婯�Ǩ�΍������K�u�+	اe]Vgx��o���~��9E �p�ߏy�~�y��4&ă�Z�X�t�9�]9�8#�E�/0-�@ 0��	  �"� ��A`��ԥ��
O-~e��;�zI¨�b�f��2����i��6��P-N2J ����C#��ݲ8�{@��4w @Ȓ�N�g���W�O1dt�ef�����i���1��JX��25�����ʣ��7p�{�2�lr.(�ϻ�JCJX�a]�ἴF�P����?��T��H��m�$i��2F����;�KS�0�ҷ�V�����4�"�q���#��L�{�j��P6]�-���׉��A�W���J��<d�Λ���t��0�
�H��!{������V���_r�ޏG��0�ߛ�Q �h�1�/�A��~�N�yk*���Yj_���
ٕX�n���K�`�XX���._S��"c*��L!�:��,F����=���C���=t�3*dUb�BAxb��L㒋A(8�Ϫ<�c"`9*^&���/�sƜ>*���l��3�H*�V�[�ډh�
��`�kM�V�����,H�
�EN��C���
�	����q!�s)1��8���'�Q��8�Ta�]�( "�2a#�6ur7BS%B��L(�\m{j��qO��+��m��0����T�����)�QR`e�h|Px.��%��G	�D ���).Geމ?��O�n��S��*���Ѣ�0@�<�v�]C���B��n�虧p�#A��E'p���:�e6� 3�Z���4���U���3(֏â��7v�WV���JE��X��8�b�`��uN�I�2��WO��Q����b��=��j��_����^��i��C��1��%��'9�!�T�t�n^]���1N{^��b�ʵV$��q���%��wp9�A�R���˹��um.(�)���0�P�{��$���>��@����>W�N�a�j�����B8��}p��p����D��]b҅���#������Y�$E�lŕ�+v���;8B��
��3��O���A����`��2��=�H4������Y����u�j�r��7�=;�9:�huh�J����Gz&Z:��m�8Y1�QD%�+��;�Q'���%��c��,�M8����n����(�3>=�U��Křv�ѻ}I�Wo.��q�%!�
�df�_OݿU�!�T�%\��Z�T��]B�1a�a�Pًh�%�����T1ZT��kÖ1Y���3���1���w�jM��^��Jg��[����O��Ɨ�&�!NN"���|>��V5'Y��S��Lf@b��=��&�Hz�O����A$7�Û.M��3bȈz,C�
����z�9�+��Ծ�_���h�7,r3D�̟��D[�?e��>����t���x�����`���5�
4���i0��E�,ĸ�l�Ô���A���軫��?=i�wT��ߑ�l����餞���e��i�j�X��Ag�lF4VtRLE��Z��)ܷS:	/��*���\�=R4^�`Lv����yo������ǯ"%�|�k
���U�Xr%`=�C����[����$>)ϲ���r��+]w��r�B?�,�b*y�/�s�k?Aʈ����T�����"xE�Xk���uw?������U�zPPť��8�'��_���;��l��R���,��tT��v�
�s����g�k%5n���kWd4���"��rӒ�B8%�%.'*��6�"r�%Pvw��p¨ɾ+�mMN�f~�Y�so@��+�Q�3����t��jqDՊ�P������w��G_�C��^�ÝW��ss��dW�����
�i��VwZ�E���y���V��w������P�ه���C���^��
�xő���fP]���dU�_r��`��&�|�@����Ttx�'g�G��?	?�{M{N�E	>�M��o�(2�ǂ�j�?��wB/jS�#!s\ٳ�9�L��1B��ӵi�,�ϒ�D`i�E�?34v/�U�5����?n�\�yIH����O�q�!�Q#r�I�%ި�(_NI#b�q��<t�e��lx��H�lS}���Xİ�m1�>����Uo��h���D��CB`�qL��+Y �R2��
{�S���~�VK��BzjE����\�o�#1���rS$��t�ӱ�%tk��3sw��>�>3�V�5�+���_ݙ �w�9q $D1#�H���َ$fk4íV������GL���^��h��(»���,v��}%��Bh�J�*�ۡ]:����h�KI�d>�FH���(�T�\��x�)I�H� ��� a\�IY���-+��d)�<ꋀ��A���m��j��c� IXѴu�^�(����"����A`�ԁ�s�VoD�Q��Ke[�D�V�|��k7q�N�3��+ �C�àv6�Y��ր����@N��x��u��I)�ed�ޏ�V����g&��ߒ!Z�-�$��Wj_���5������O@���TB�/� %q��\��I�0|N�sd�5]��S�W+�3�Rӈ|��aY��쩱"H� ����2ԉm&xk��Mu>�ֶ�~j� C��sQ��t���;)�jn?t2���&����i��LV��w�QS.�Kv9pFh��s۪�;����� ����`Z��*�}6�Wm��!�Τ���(_����Z�˨���}ޥ��ZH_�ƣ㓅瓺�w��W�AzO�y>�rF�zZrY����Σ��_�j4�{�),�@qy�S��|A�g�������7������6��@���:^�?�&��yi��C�V�i�.�<���K�S�$l�o�ÿ�ξ���pI&�Us<FSWx��O�K]���O�%��j�a�'=����s��勃�U�{���'��x��
b����LS`P�֊�3����4�
��zG�0_|��gL���i�Ԛ�xXԐ���y��g�zEa�c��S�*�����;�+a\���D{�uհ��5$��S/����I���[�qB���f�\����P��ɨ�D�VE&�x��M���^���4��(��H�>�9�jo�n�ʀ\ET�Ƀ8���]�D��S�̣�ќ#E�'�{�7q�?}���7ܑW��W��)��@��э�99���!~����c�#a¢��m6�E�~2oJ^�Ty.��I�Ér߿D)�fXs?��5u@�����&�� j6n3S�Ѥ����2c1}(�M�\O�i�m���k�x�c�C�k�y����fR�mE�/��W�p\�5���V��0ل(I��(l�e_� ���Dhry�p�R��_iK�s�?�P��T��Of����֡)}�GP[p{D��0�FR-��E�6��n��,���(�pe>|!t���}���1O�~
E �$����y��x�1G�8��Px.P[^Ƨ"L������ؐ�8,�����$~Y\���=\��mp�-Y��lt�W���0c������O�\�-\ٝ��*+apV�3Sad'�ƚM�G��d98HfG�Š�AЛStu�|��$�����|J�h���
^������[q!�@��pY}�5�o#�4�]�2��2�nq�ؽYV�mE��ʊ�+'5�q� ���d���4���X�U-���k�X��b������q��r���3�W��}�$V���+ _E��}?S]U"�E���m�)��2X���M�@�z�O��B��{�/�;(V�ss�n���?�� ����mC��M���.lʄt��� �GQ�U1]�a����ԡ��X3�`�p-9%��M���P�0��{��kq�=g2%�~?a��dR���~���ik?�RU�.D������&r"��3k<�z��L��F����_�wT
R�oнy��VW�4��^����ͭ#�`�
|��`�n�RK@�(��~#�[�b៼R�XD�A�#�b7��Zx{/Z��k��[W�o�I���[�L�K�@�lSN���� ������CQh�H�D��l�`Wj.2J�_,���yh��`��)c��rq�5����N�)���j:<�L��(��>�\���4�:0����fU6���?ė�eh"�F��L��A���1+��E	r�8��t�06��;�N%V���+~l���@c���E$����lP
��Hҏ�<�,��\�<yC{ʳL@:M7�.O��u��р����CX�n�q�C�<�'m9���;���t�G)����T�������^�0���C2�:�\U�%��֝��cr3B"�n����7�ю�����>��f��CA�ࠒb �	����Rܖ���p����/h8�Bx4���U���1�^�=��2�aBw-(BP?�ZHZ�w��s�*�Pw�m`8��ͫmB�U��l_�sA�Kl&�z�����ry������[g����ު�~U��D֥��U<<����njY���et��f+z`��+iT�A"�l3c6��_�Ì�*�����4#s8}���>Bs�ɬBg$��<�3>���ם��Dt��%~
%����I_��@��7����Y���֓�����5d&(q:���C��������nDˮF����""�eq����C�����`�=�?�?nP�@���l�N"A��o�%���5�1�A�(0�44i{�T!6&4���~���"�+$u�`��$tX��N�/��V *`�Df�o�C��SLNae��V]���	��%1s�1��Dr���[�*��ͦ �G��ޏش/��!I�DL��V]�����Qd|�Ty"����d�t1ؔ��x%b�M���ɤ
�M�Y�!��k��=�[���l"�&lܮ����s�.��KR.�M��m�U8W"vl�
������ٳ����V��[mA�+d�FjO{�������3�3vd0��~�*n��D��C!�����-��l�q"JPn�Rt�D����V���F�ֲ��#�;�|��U�G��a�bɕ��	�~;&'@yp�\�ߧ��CQTC�lFe�m��=�XH�RﺹniS��oв�_m��6�׎D|������P�Gx����E�XvO@�ځ���a���Ր�;��N3��{��R�>s[āt�5����k��3`�-�V��Zd���љ�c�a_��0�F��.#\��Q�2�Q/�������p���<W��W�l�G&���ې�>��&6	z���uC�˃�eG B����0\q�]t~�:f�̹���n�Y��զCځ��۪� (���5���{V,�x�q�C/yr�#��5� J7r�hD"����*� nz7�0i�hHA�r�����jH��
��!YζW��e��n�=]��>�e��X�~�YԠe�������Wp�e9����1>|G:ǳ���q��1��냏"�E����㻁��ĥ��RR� z���hu�ɾS"c��F���B�f�4��W�����%j���it�^�4�J򓁬-�������?83T�(e`��瘧r�2Q��P[V5�2�[]���,zQ�LE�E�M��v¾�<����>��7А8�&����ȣ�oLH�/�� ��{�{s�:iL�f�#%��<���h�D0����R�|�����=GC��{�:�$�7ȿ�e�=�}�di���Żi�S�X�pG�����P���;E�1���|� �g.*))�|*��A<kÀ�� �Q6s$X��Q���*�q|T u�y�D��y���B=���ը(-�VN\�J�2�P}|a��>jm�:�Ƴ�l���IYi��
�ȭ�@��^�_'�ݛxޫ�|���pY�����mr�+l�ӆaHӍ%�� )ߘ>G�c(�L�d������~<�Y'��SW���M1R�݆���#��B��x��:���e/bѬB�}����}h*��8�JH�M�}G۸�@M~JBB�����l48��ۺl�˲b�i��m�!W[���*
-��_UZQ���'����rY������;c��UD<55�$7��`�7pJ����Q7� Iн�EP��g�X����m�{�:�S�t��"�ͩ���tp\����Ut�T�s��o�Sx3�0���Nz7u��2ҵ<"��q{�-��D��zI ��{�Q����F=ڋ:�j�!b<Ä��7Vp}��΍N;��j������J�6�ʄ#V��2�ja�B? ���J_����eͲ��D���e1�+�h�����X�I�d��|��v!���p浧�wR�i�wP���_��-q$�o�F�]���k6��~��lG�Ǝ`Q���pn�v%�ENߑ��	I9f���@WL��x�U�=����d5��{h\���'r���D�߈l�P�uu�z��k��c���-����B��Q�2�O�gI@�������g�KF{�q�f�N��NZ���OL��9	�]&0�.�ۇ������ra�[��
`�A����P��@aa����L�2m?�m�ֶ����6)k �t��J���6	bVs���h�﯐�yЋ�g�Xq�tI4��������3�#��j�3�g�ؾ�E%�L�ԛ��U���f��M �����S���d�iq�o�:�&7�RiؖRp��'�=t���j��z8$� �A�#��%>��ѓC\L�n,},��}c�n� ��h�r$d�n��9���yF%/�%�v�G�t6e]S�s�F�KG��3AM��(ө #X�g�7�<tl��/T`���iDX4y�ős:ߑ���w�ߢ�!����k�M��J�Z����XՐ�?��ۃc�D��rQ��J�;n�KH�,��j���%�����|�cqp�Wȝ+E���N�)]����C��QWA�ǋ7V��]����,$�S 5�T��tݳ?�}�O�̊ӵ�1�Ùೌ�}5Ү�w6���c8�*�c7�}α����~``o!r��UWG#�и�L<@_��e2i�8����Ac�HM��2��i%޲�u\{�"_v�H0vc��U8�Y!:t	��܉��{����b52�Ͽq�1�i1��ۨ��/��HR%�܎_�B�S���a��$�hB��OΩ�t�fQ�_{�W�ǲ�e<��~ǘ�.��L�n�%��������=�����1�v蚱��'M�y$X�jn�lC���K	�U�$>2c��5�2�QYM$�PR�^!���,�/k�2�:��tNn#��`�b��J��a��d>��g�X9}��(�����_�`U�^e��"[��n�;���YMӅ�˜���_W�YjI�\�N��};f�n�w�����j/8�Sx����ٕ	 �
ʐe�6�{<����{��-X�,Τۯ�5u����at1
8�`�ιF���lP6����wE�R;�}����L�֢��Rй3�D�j.
$���9�H�8�-0�{5VV��|
�1cj���	��ǚ�^�h���<�?'�֮��omtR�.a4���eba	Og���ކǒd����觳E@����t�Q�-s�j�6�.��c�����ٔ��b��V�v'2��i�𹀝���F8�#%��+_U�����^�p��|_:�M.��'�3F��d��>M�7�Z�ǯz2�3 \���|�E�g㰩��ػS6X�O0��!��O���n�۞�z�Qr���D�p��&V8�T�Z;vS�}4zj�8����[�"TL�y?$Sj��I�����X��_�U�{�o��d^��]�]v6.v���ڋ�2#p�,:j}�v
�.|Nzfi�}�:�P����֧�|�cﶕ���:�{�(�'�2�gF�Y�=�@�F��}g�PFfZ�:�וN'��lK��Y���6�pjQ]@>9�孬����`a� �E��������c�)7���Yt�<2(H�@+��gx s�yҮ�@2�"b���z 7��Ȥ	1݁�)Бw�"�`�77�Ǥ�q�(������a=!N�)��	��,;M'iG��@'g�M�E�BB�~3T�,\u�eFb���ad?��R����T�!�j�V1lR�y �S�h�W�*�V���h]|e�`��D$�+�>��:��Fi5�r>@];������h.���̯�|�h/����WCj9�}�?�U_珏�.���M`��d��'�1��X}sk63&��`��q�ૈ�	���tkUF���G$z]�����ӕ��C-O�ۛ����m%�E��T�015������Kw� ����FF�o�K�kh:��^��Bߗ�e伅���ssz�&C�'3�c�)�(���n^��>x}�t��H�֜T�m�t��W�S���{b{�);b��xIqC\~�H{�#J]D����|���;:u��=2�e�N7�IȤ|���7�",�G�gg\N�k��� �f�5>K�,\0C��B�]�	\�llH|83h��0�q�l<	�M�VR�X���Zms���0"�Փ7U��>H�-�i�I���Ц(Xo�RK��^��������2��Xz��	w�`�E�.����\28}h�<�5�:!���~lA�`߅P�H�hbG�5�ֽ�A�7C��ǁUr-H����`��ㄒ(n�k���ȫ�F����@I�]�fy?5�?��O�I�G�g�%#/����^���t�k(]�iIO�9��7��xS6�T��hfz�b��Q[�Jނ��#�S3�8
�^���cyr~�6��:��ה����D�����%���0
5�\S^��sQ���i..u �_b�aVv�Z�T� g�.�L����ճW
��2�qof�m���Zg+�H��h�������� q��q7|�=�1���v8bP�d+.]��!vm!x�`ƒ;7ߪ�7l-Gg2�=6/�� %h�����0��C��2&#W�xV�V�CK�ji��TE5��l's�N�A���r7q���,/�䜍5��	����|[���pu���� �}�����f�O��x�P0x �!^�ƦE��Y�p�B�P ����.�ˢa��ݩ�M�^��1v��)��gK��ǿ.�T�Q�D�KbF|�R����\��VuIn�Ba ��Ő�X�]�u����Ϯ�.�XS��YE��,��VO�vׁ}Ҿ�FT�"^a�y�J���G�׊+�©�1;�+G��ۙq�Av��X�r^Ef��*,����6�Y%�_���V��.ow켡{k�@ /jLH:�h�C'Ѱ��X�m��o���BCᆎ~	k'�E�H�V��#��0��\ffrNYu3�Oq!��� j@�C�K�Qd��a0/��y_3�tr>���cY���tỔ\�4��ȳ8�h�7��t�G.��޼���k�/������J�=₋,T�`�&ҵZ���i�E=���a�rm���$���6���/��y�]+�mzs��:N	8�����&t�a��舳c@��P.R�����MNDdT�=u�|ٴ�-pּ��e� �E#���v��D�[U2��D�!R�uЄJ&�u���l��`��	<�D/�"��\m��鲐x��1�:xO1��퍳T�!�+Vr4y] �D�� 1H"������iQ�HR���5!����I��s�AҾR�U��Թ�aV�;��V�z4j~�ayq�Lh_�� ��P�am��Íy"ҏNJ��[��ں���2��=_1�>i��q�fu�N�<�:�m��������x��7���Y ʨ���u����j�n����׋ǌ>��i�>2Gt����L��������S�/m�J�-s���k�xG^�h;�}�e/���y�I�Uk��D�^D�H~z�jGZ����&���sㅐ���i8��y�;�N���cCX�K�����{�?��OV�ä��#o
@U��O���گ�aL��Oƻ�ᵮYxQ�EHPwnSU���[/��������T��o�C��4��X�|�r�t��t�^q�2�{W<��1p{VQ?��,��ȁR��{-Ϛ�'�J��-s;��;eEx��`to���`�3�=�m]���v����PYxwwM�lz'ԝ#3�%�Z�?�w������_���ܼh�9��f�[�R��ཌྷ�b�G�E�/�@�b�}��I�1���{��~T�����)�|�<Hh�Ojɴ{h�=3�t���>�����r[�~]?R���dHy=0�8\!�'3���8�^�&�E7�W��;����l4�ߢs�R6��^b�gE���G-N%�%vqh;� 냹���#�'8�i�L�6D4to+�W�@CM _��"(��p &^f+�1��J���Kp�3:K��&@y��s���|F`W\/K���cu�����վ2�-�PRfa�H��V��Y��J���S�Ϣ��3Q���a�u�]�����Xu������	�i��$ �5��ޝ�9��B��S�F,@w��L�������WdǴ}"Bt�U��a�Nr�:d#P?�?����;����'(.�:�ۉ�<���7�$1��(��x���tm��@������n>����������jU�q�?C�Y2��u軗VW��E+����p~3
�[��>��A����U@.�N8����d���?Y���x&�:rɇ��E�Z'ݱ��ΜP�l>gs���ObE*RXn\�=�+#)ь�e�}qΩ5��n��eEOp���k^�4e6���dfc[ĥh�Ia	Cy}e�G�
Ņ���L}����������Q-����H�����8L�:��O&߄�E�fn�i�3F�z#��}�©x����~�(��Ūs)�ܾ5>�������`u� �l�I�q<�v�����Ȃa������W_lʙV�dk��0��G;�<�	h8#BFӦ�?S/�B�m�^��!ߢ�)>$��lJ�����}�P,�d�E��$_�D��.��`x"�es��iT>����n�zD�ה�0�j�/%��)�:FL�E��K�������5�IL~	��-Rѫ�H�I�Έ�H"�.��)1���I���I�R��Z�("�ʍ�>6�9�c� ml�j^b(U�B��F� ��X���te����Cv����qԂ߮���m'���h�~�/4��b�Mu{�����q�vDq�˨��a�L����'U�(�G�!t!��n?]v	:R��
����䷡��!_�&�]WS�n΢D��g�1�n�Ɨe]�**!�v��=��a���PF�Jm�!@,z;(jD�<.�hm<�Kh@b~��\��M�,���Pv	:�I�O+\�����a�����b�����F�u�&tIxͩ%7�z�H��� ��?�?��������(\S!�C�H� �+�F�3�E��p��wl��9��Ι,]|b��Ŋ��0��w�����o��{�D!A~�`�F�E0y&]�ʊ�|g�A!�_|�p;qL�|��jUs�qp�_�{A!}��6?���_$0K�)F��KE�q��{C�}�3�sߛ�x,�Y�(�c��Y`8�H2,�;�T��|�k��QC
x�Y�z������{7Ș����H�ph�)��1w���h�ڐ�K`a�����z��|��s!�bܤr9c8�l�$Y$���7���N0��v�)��M��OC�y��Dw�s���4�}-�`ɮ'��t�D����75ؔc���V�����������f��J��/�%����I<�T�Y��nI<V�;��!x�YMgy�3ϣ����:�AcN1f�[ ��Aߧ��%��^4~��^KI�QJ��Ai)����i�F
���o0,�� �C2��-%aO�Ǉ �`�t��
�M��u�34���� ���������O����{�>���&r)���y��m�o#�=���?��w�N�Y����*����s����Clk�s%�R[������j�R�"��B�hx�6�Ulp0="H)��d� ��(B��K������������|XsHq��8v�^� ���[���z7�ĕ��VqZBDzS�;m-��m�zL��h�m�����a���^<;�|&$�s��!eԵfx���3[���7j�ҥ��7��l�m6f��X��Xy1`/%�`�5(i�C���Cm�0ڒ�0��چZǺ7�3O�^�5�/K��]9��A���x*ϲ�e�����������O�VI�,���X�!u<�HP��\À��&�ۖ۰����̛�%U���R�rEu�̺�rZ��\����?69��C�3�i玊��t����cq�'G
�8��ܢ�lb�o3�x�ޒ����i�����S]9����(ɤ��	^��$��[k�k�s�.��(�f�}  �?w�Q��JiM�A��|g�<E*���� ��S��� l%!���J;48x`c��*@��1�1@����M�+�o��p�U��xϟŨt*h������<GYXl��(=��*A0��Ӫs�~����C�]�eG�>��C+��C�8c��뷲P؛綳M#{���L���k�:ͣ;l/��z3���c����k��.���R�MrM>Ğ^�Ň��[��?
��o�=k$C�Dl~���N�#�/k�ǯL
�4ʻ&�]���� ����?(VG�rU���8�eҧ{�@��-��6�,X\��G���i��TP	�|�$�1�ͥ���T���`p�۠���BɄ��k��F4�4 ��d����X5��I
�����.���w��.R��1�̜�hQ4�|�*1i�%��`]2��mvX|��R;���\���^�1���"�{����Y����t���������v�q��;50�z&u&�IL��E�hv�7_l���#xiy�������`\IX�i�M�y��MD��G��2S|f�j+^�p����uoa_��l( �U?͢+L���뜊��;���~��F�G��\��F��z���k�v���$��A4xe@������q~4��B���Ȍ	�7T�d-�f9�ىPX�`��[��xު��a�l�5�\By���Zcǫp�m��H�����#e�W�����V��i���yѭ]����f�.sv�KOx�~a�J< �&�9L��ʫU �����ڷ蚺���ʇ(b9�^:4�sI��N�~smvlFd�<L��D�A^8��ʘ���{�_�7��i4��tz��60҈�"?��遑Ԭ�����@�C�-@�#);w����P�i#���$S����ӆ�;|��
���JW�``p��N3�}��qn��2��p)y�+��6�Ԗ44����f�0I$%�������H�2Nj�PC�}��Z�d�N�LA�	�2�aQ0�����o��(�D�aIn��Uv`���Ç/�Q`Z=�� u>�{_����y�I3P:w�&
jG�P�3�H��Ti���
@ڄ������zi��>[�҄+_��1O��:��ls��:$�K�E3���_�f��?g�C��$<c�k{�/�P�qˆ+�*�SHq����4���g��OD;dY	��ͨ��o* ��]9j`�a�GT�Q\���*Ì���!��Qy푅��r�n��	wZ�]"3op��Ǯڣh���I�r�V��7!ܫ��PtKד�tH{_½�G���H݊y�'��#�m�����ݩ�s �\�h� ]��>&�'�����冹#�֢����g�>���0��r�"�~�/�I,&�-7����~&����F�2��f��@�n��)x�ߔ��/�h��
�yb�Z�ߪ68>�2=�O�U\[���2#��%��ξ��r��v1O��@qk�P*䶺�K�k��o�S�Wm3S��I
Vh�@����jm�O40�3{�S�@HЍSa$~<�'0������Z�C�ć����4�`g�Y��P�����[�`�ƚ1�H�_$^&�I�'$��6{����lC�d��L�����?�9İ�W�P����ZP��Y�1ܥ�S[�-�(�m�](�1u{�u���`�<��$"��*��DyƮ���"i):6��n��ֲ�g�XY�0���mD�`2��&�~���k��5$����v���N'U��[�[y!��fݟ�W[5�5"'���ɽq�䡫"���K�A��N���8���-��+HX,~����OS���S�=���|��Mx��N�.�'r5�����/,b�5�O�S������v7�A�e~뉢����:Y�������+��I��iP�8c6�d{�m��R�?F��|aeI��@�Ai�W�{�]6�А��>#YG����,+�n��S!ΠKE���z_X�A3�U��S������	+̷˞�o����^�c�FJ처�
E�Nz;,4�{<s�^�]_=��g����~����9����Ǝ��)�6�.��`!��.���r�v��]]C��.��c�R�*Fo���\�(]K��$Stzz�@���["<���o\T�4���� �2w1��K-������ܕ#���qɿ\��G8@n㋸�g�1������1!��WW� E�ͤڽ"�C/U�;�����ȧ<�!��a��[�b�;yL7}p��.[�$*m!��O`��%��ȯ`9�l,�AYTׅf�H?��xaO���e�{Z���h�#���"���;9�#ѿP�(�u�EtR��� ��SZ����e��@��D��(c�g�:-Y	C�M���uq��b�S�3��?.�`ii���SC���	{'�./B\]����ƠtV�s�����,�8��x��pM����K>ӽJ޴1�ߺS��G�m5��ol���oۆ�gݵ=����=�� ����f4����� R�(�`�@�}�� �b��ݣ3�5�6����2���R;�*��`�!Ļ��Se	5Y��pv��E�.[CV��!r׹�کH�Ka:!����"�8�����&"q
�U�
�&K<���|��1I�z�Ͽ�*M:�\��sGi#4���b9� ��4:�[X �,\3�L��+P�Z��`���Y5��备c�lN������4;Q�	�i&�c1���.t�#6ةep��(�I��L���y$A�X��'��0L߆�/�c��mK^�A��@�P��C=Ή������]"����ˎ���rc���h�7���Uܵ��_wp�Yh%�J">����*.�,�?�Ԁb+?L��nq��Q�������7��������ݘ����3�Ӥ>:λC\_�GD5����z�T bܔ�R���59Y�S���XD�J�ܝ�:��L�gmK�T����&@�߼q�7���)}�[�\�L��������K�H�k�# �11J���K	�z�k��hJ4/ ���IVQ%��v-U��֩�1���5�I:��x��^��ԓ*�c"[��M�'	jx���}�'����+��W��O�(��cߨ�تM�3Ѵx���d2+�҉���"�(��D~J3b�܀�u�y`�[ǩA�K�O�P�0��A���e���ާ���RS�Z�ii��d�$��D�����+oJ�$��M������($fu����o�����X�{'�>*�u^���RW�:`"!vqf�>&ֺs�����k�k��S0���v��<I�d
��vkQ/�����C�=�J��F&u�줛wn+�~��紐�*S�D?/>�t��`T�ڛQ����9l�o�(D��N
���^���-1HI����ƷFgq~�Na�H��þPf�C�lc�3T�������Φ��ě]	.7wJ��T�)�1R�*Q��������uԯ|/�$;�x��R���9OQN,�y���O��D:�#�g��^�tE�E�;�gD��n�u��#i2��m�:o��R^~X����3��{w�Q1%�1��p�K�Kj�#)�����Lv�n��9����O=�c�󤦯��̚���B���)����z����u���A������!Pc�I�~���9���@��� xp�^eo;�����+�ە�5_���*-�������Zy�ME��<g^��K�|'�3z�0o-���ǰ�|����C�B3���)Y�$������n)�T��~1��p�-��KE蜱�����Y�/�V��7[����<�=F�n��3��7�����y�&�:�
|���P�-�M��B:tO���f�x�:k���Ȑ8���3��p�ֱ�����nn/2�4�J5�d��܈���9����A��7u4��و�sX�ŀ�j�Pe,VL���Z8�v���Y�R,�#����v?�@�S�	 ���.��3�tw��</Յм�0�F�m�[[R���8M�����_��C�V7i`e�]^;&��B�xz�M��c����t�@��T0Ѯ��LK�P��L����S�@��K��v�1)VL�I�Q�%g��b�RT8I�7�2g����VF'�Ik�0%2J,�܄�CƢ�T
����[��V�G��W	n����rB�V���1c<�ym�.xl�W��6�>�CIr���SQ?��"�C����\P�/f�⢡D��l���A�R/�ꐈ�����9�4ܑ��a�w¥�xS�P�,��.����� �-T��0[�G��! 'Dց(����zD3�y>�Rf)!���$�<���~�7��N"�L=$OI#kz��]��)؂�,)���1[�G�G��9�Md����S�Tt��u�ܷ��y�_b�9�������=��Zb�ͻxIk�딐K�����ǜ��V��V�w��/c3�Nh�oh6����^�z�S����"T�R�2(���5�1~�(���CC%�&�����[)���!y��J��y�m�'����5�������"��Gq�O͠y�\�F1~��V9jj����3�˅�e��~�����]�}F�v�R�y|��0c��~j�m�.��q�L˜��H�Ҵ�<0}=9�~Ίs�����P�QLC�R��e��/��`$��=�Um^���A��L�_�v�A~^щ[֪�mVN� �x���l&UmU�{�X��
j��=��"�@�\77𫛿%�|�C���F ���
2�P�&�K�F򰂼�"��ݟ\�e�4�l����Ǆ����$nXc��S��)�0�?�
_����>��tE�D�v��z?��(�$�s�!��Im��� 1�.z(�f�gx#���O$&m�s��/��T��W��O����-&��8t ���	<ڰe)w�G�X�.$g�#��\.2����ʔjS��~��1�h�[eYP����H�����C���QK��eRs�;V��J���+L���I!�MK韦xE{�d�~�v�DU!
�6sȤT��R���ڕT�%����߄l���l]l4��e]�C2y��A�q�cῬ��r5�̢�vԋr�8k��%�`�w{I6yi_�3�Fm���U�hg����XS��&��fc�����jخ_>b���iְ��wM��1𼖎$<�f�/&�����	�{Y"�*:�w��=5F���у9L�R�g�Ƙ��R��*Vq��{8���pW1�:v��`� ��̴: ���M�?�`_]*��� �N>R�=<��<st��]n���yϣk���RP�8��'Kb�G��9��^�Ik��?sM���Y�~��O�yp�����X������Q�^�
Τ'�D�)\l*���[j	Oz' ȑ��wg"u�L�׺��|����H����;S��&ª/]�l�w��m�Ӗ�s��֬�#�6��`�`�+�-q�:7ǉ��3c�_�.���.�����3f���=�B�Et��k�ޙ��בB���!Pe]k�����a����	�`*v|����e�`s�����_X�0�a�-:p���i+�/��EY_�8��[FY�!���V�$�x��ך��|;�
�JB�T��ښ�]re�R�[�r��ZE��<?k�k*d��Z�,vT�s'Ϯ��{6�b��T��IӅ�̻�j���yt��& k}y��J�7
�DF�@�^f��/�w��I�Iӷ���+;hd����9A���=�,�1v�Ec{�a��D�B�$��p�dYbB�C(��<���,.������i���H�q�#�/�k�Sr��I��u�'B�&?FN�S�����@۽j��iP2VW�'��{< q4�8H�p`�ppG���)�)yifKW5����Yfg�qk=�n�Xչ�s�����L�n�
�2�����]ؙ�������B�����f+����)��C(�I�>[ ��(j��G�[��ro�'��j�1�'O�8Y�N�Y}���H��']t��g�#�$���1k�h&�p�u�b��2�s����|T��Y�������;�G����5����
&�a�Ie�VyE��,u%}���ə��n �!�e�D�݉�	j�:]��g�O^��T?���I�y�]���8���eW�u�#�q���6p��5'����j���(�S)�u�&��'�'���l9_q����8�=o����p��0�+Ut��6���K�M�pW�&,l��Q��^��Z������T,��<���W{��rrMt{�ža�t�-{# ���UҌ���߹
�s����%��!O��_V�$@>�_�8�vu[���N�Q�'Q^y�_�����񱤷�
�1y��!��@v������H�Y*N��;��]���-��4󈮕�u��6,coCq}��5�gQrW]�4�5��I8򂦷���'���������-��D��e:���GFF�ʲ��3Gp1[u��'m�i�~���8����mE��~�}`fJ�29�:�������{�咤����.��O	�?A1�7R^�DJ\��*Fv�ͅ�0JI�QI��m�M��A�r�j�ejIR�d���G�`�?';�Ş3.~� �.c�8������;R� m�/4<�ƩB��~f�hф"��kd��*.+�i�1&"Lg�1T�I�sF����j�B�&�"��Z�dV����Y	.�.@&[���]Ϯ�^X{��4��R�n^�v�"S�݆x��} "Y�Mﾱ�M�i�u6�/�Ƚ��LGԒF��#���1N�b��~���|Z(��h��%��	c-6
��s0qE�"Y��j0�%��Z.�zml�����P���,��>w5]i(�qN+�_!.��[�Qsq�r�*3�G�}BeX���%�Ŧ"���\�� �%UOȂ��ޚ0�U�4|/L`?��;��4Ѯbu9*g��^�M}V���sq&���{9cc]:����6b���V":�f-�Z`�=|���LȰ����3.\*���M_B:␐�}��+�9I4r=4hy,�<��,��V1c�F&��J�V��䞂�L$Z�q��_o�<ѣhU0��s޿�{,v�)�L�DyVC��?q�^w��['6�VV��O�AV/���)�2qC5 \��(���>�M!�(�ݯ�3�w�:�lKgI�\i
�lʔl�QRs:�0����"���z-=���`*?ô�}�#KM�S�A��fV@Xč%���֐l�p��W�;Ĵ�u��q�i�ڀ�#qX����֍���7W�%��K���"�v4y�zz�Pe��d��JW���?gv8���R�����f��P��W�A�0�
�K��:����ɜ5�]H|K�&q�c\���j�/��r��'Q�7��q�OÍ<d��;��S�ֵ˝w~ze��]��sm�W����o>��\#�ᄝGv4Z�J����1t��[�b��׏MB\�rr���:�;���K��M��pA�W�!�5_`칓�'�����J�Xb�8�萈��	N��n,u���jMzR���q�N} Ơ�l�pA�<�9-=�,=kR	���1�?�4s�N3u|��Z�)� rY���t-*�����F��YG�;� שgu롹S5]�m�G)ad����T]Uhȣl���ibo)�6T�v���<&Ӽ�;�V-=]�\��r?��Q�u��!}>��mr���}�j�a��x�����w�,-u���Qn���=*Z���yq,��*�[�#�C��DL�-- �Hu)�GP8����݀K��{�(T�_?�흱�d.M���k��Y�6����Ю����f�."�U7�)E��J~;U),��5��M�ĸ�����{ES�Щ���/�����S���R�^ ��0�����0�n����{K�qS��w��Y��zL��=u-]��e�N��1	��IN����yH����k��?����b�o['��?���9�JfV���\.Sѿ]�Ȍ���DS���x�<�?���$[54��w��0�b娢��ú�ʐ�U���&�;�>� /ݏ�fS.F3@����М����q8{�d��%U��G��)�0��)���U.�����.(��9\�3JU��Kl���x���;Q�B��$�����]�k�����ĉ��<�7��Ϭ|����ė��~\��h�Ը
{�7�g/$n	����I�M�Nt��Vӆ�����T��6J A�L��<��OHqr����n����r����%8�nj���S�g�(_��#*\7�8��7�par���V:xrˮ��V��Κgƀv-�R_�y�dx�T��v84��Tr7#^�x����p9�v�ЅIi�oz����u@��G�������W��h�c���7w���D�����pы􎘺�Iy-U�75w��: �1��G���p���)CH���X�5Ը��=oy�\�UeB��^��+��v�%G:�dF�PRA���7�ct:7�?��,*�����J.�qjN1�YlC\{m�˞��Lp5�ڭ5P���2��o�	i�T@l�Rk��K������sÚ๱qH��d��ߡ��U�
�bD���\޹"C^z�٧��ue	E}�	�Ř\9�8�m�$q��o�%���j�MX�Ҝ��1ޜ��r�wA�S�۾ә�FQ<�+���w�.�{��Fr���<c.��$�z���'傖�4!y�^�٥��� ��h�v1�K�ô�!��x�n!5�wu63ԦFd���ԇu����%�S��5���k�N�޼�M����p2�xL���#���������K[8�[�Ծj�ۨ����Ȣ�/�!��
�!0�޶��O��G�B�s�I�~�H:oK"��|�Qd�8��ۅb�2H2�J;���=��aD�--��h���ܨNz���$���-B���i}�&Ν8,����8���%��ගK���X�>�/���v�6hGr��C]	��d<����z�~�:�{(W��)aSW�P �ړK��.��j���a�����L�<�Bn���:�

&���t�~��!5L/�抐���d�Dg4�|REB� O�Pj���k�E��v�b��M���"{eڶf�j���9_N����J/jU��k��G�kkkD��^.}�^WA�kyK����*��䅽ZC�0��pQ��)�gt��B�Ə�*�z�O<�tiK�Ȳ��%�v���e�_�������<�*k~lc-ܼ��ٶW���P�7�\\n7�s ������LcX�l�{��@�FL�ء5�I]WVb�d�/���<5�Ġ$�^�¶T齺���m�=*�Z�� ��e��DKi�Ә�w�d�\H��,�j_r����
վ�Ζ<&��t���C��
Oʱ���J������Ȥx����N�!r����\J�<���Mnz]X�X��K��^0�_)Yw�m�e��:q�/���2�fȨ	�G/����ȾL�|��| �00�,�Y،('���Y������6D.���J=F
l}��{7�[8��sY�a3�D��xs5��R��pyR���l���GUWA �"��?(�@��+�	����P�?���8�iı��_����p��玑&[�M�+z��6�8?�,
����t���!�b`�0}�@�p�/����Q�>���M.�w#�;��xU 
p�C>"��D����g_��j��7����Ȧ����hE��O�\2�T���<�A��}LJ����R_V�jR�bc|ǈM��P&�E����P��޾�
2�!̃�����m0FD[�E2���� ?P���n�8cԜN�Ģ"z���D��}���n"���C\aXn�۸�,?+	�A����`����1FF�,FnG%��R�F.--�i�R��&����
�ꞵ	L���w��@(d��5h캃�ԧ� �n��ͤBy����*$�p�����r]�k�\�;>���w-����kPoݶ���<�}}k�f��J>��R�}���m9^�u�����a�����b+�NeשӅT>�24@E�:�GU9
�%eE�1�`.�p����,�Y�t�S ��^��r-�x쇭w��e�^�Ʋ�0�ǘ'������ XAUh���c�ϙ�P��^ة�sI�cyA�N7��SA+�p���U��?;��x��R�n�E�� ��*�i�1��ƅO�2#MhW����ɖ+'0AeJ�1����L�WNԕ�뾈G3=�ߙ?���UHC1/����Wn	5��y���Z�&'|�+ac���}T�_�a��ch��yb�ր��Rvi������p�i�<�[���X��C��������PXVn6���D�zvZ���B˫����P��B
��� !<�9n�~�/0 �Y�>H4���aF��.Wr�E�y@�9$ t���e�G�ϗoF��9.�� ,Q��c�dE��`ݴ��?�zs2~!_+��8Ɍ<�5#O�?2���n�j�nj�=��C=�t"~Z���n�������K�&;�A�T���a��r��k�4�& Ǵ�s2i�پ�C�-����;1�2�P�c8I'��ᢔ)���@�Y�ɳOye��Yy���UandfT:'il{�3��C����7��֢��1�;Oa�Ƕ�ܬV�=MS�̋���q���Ku��<t��zѹ0�ly~�E{5���9g3�v��mp���)j,����Um�f��������R@�cH�AE�0���ێB�Ra�� ���{����z��� w���9�y�L���r� Q�1[ �Gfϼa��0X�r�x�pJ{J`e��9,���{7�rXqx�=D��Ҷ�h*Ԓ�7�ecc�x\p�P�W���6�ҙ^��L�,Q��."�É�<�v@)�Z�Q#F��oU�M7�2�����h����<�S���g�~T�(>"�E���@o}��ʏn��H�L�kω�����$�11z����1F�������C���
՞�]`��  �����=����s��m}w��XT�S����y�����.8X���Z�|N����c�3���~�b�~P�a���[�ʔ��I���'�5Yca��&RǑF%�ڙ����0yf�5�Bc.�m�s�z���<N>�K�4�	FO�^wq�r3F+9S����J�d\��.�k��YOZ՛;`��S�&��"h�Ӳ����B��U?���*t�Y�B�Ɠ��[�RD����9b��������0=�5�7e强��:�q���+&��~��K� �g�n~\\®t�S��iǮ����i@���4�nv#B��#��`�	��;������V�K���L1���`�Ӈ�΁�I�?���Z ���F��h~��md�G��^%"9"@��d�ξla���ͼ��=�ę��V�:/�^��e�e6{���ԛ�u��G����pR�4�UFP|6R��OvC�������6�i���-ֽku5K�*�V����uJXZ�5���X/�]:[�4�o�}C��ߜ��5�=����<��81L���GȂi.J(��Z��x��%��!Dme�w�IB1�z�w���s7e���*�d�{��y�﹍}N���� ���	�-�<nO7�!�:��2]ZZ�sY�o��޷����t����ܦ��n��d�����"�u�}���K1�#��U�3h�|�i�a{��ڤ�"�~O+k�l��w����^�$Y�h�mA���ho"D��!I�4��_܁��p�Kci?��Nhh�p=X�)�Y��pI�..G}���Q 
1����hA>rȞ1��~6O�;�,emY5*U�A,�H9��]&���[�%��C^��⻟�w9W����D�u�s�e�����cZ�t��'���5��p������F������r��7R5ܥ�+�i�e�\�)�EGDR�Б+�j������x8H�t�����!�I�N ��a�ݱ��D�'�V:�i�=�7y�w�A*>�a�f�D����vL��n��ː��s�Lu���d,��B���x@E��q$�M�m��pN�[�&���X�p�b��;����008")�L2³�Īb����ts��i�3Rļ�<���.��#n�=څ�b��ŉIa��؏���$W���3��kn"�sx�>��� @�jRYv�6L��?s�6Av�����홦�J>�������&K3��|��Wg�D����AU��w�5��:��P/շ�60�+�@ ����?����)��%m3&�x��w����(�s	��n�H� 8�Z�y�ޒ�?���ߵ���1�gk�����ՙ��z�ۈ�d�
�����HI9�(<1�G0C i�F0R^�RvM���RME�u��k�#�,�DFlY��<���x��/�{R�KQ� k�K��"��?q?{�\��Ѳ�wW�Oz�����F<�6z�7;��6�H{�����GlO"�5 #� ��N@y��@qO�� �R/�y�~����H+��и\�Jt��:)��y4Vˢ��YA�ӲH[E��J���l�@�j�ێ/q���P>w82����7�lT�k���	�˳�S�mˇ;�H}��*��x���	��yF�3Չ��R���Z�z�f��i���J�`5!M���1���M�s����A���t��<J�� `ʓ�n�6�5|yv?MT�F1et| U�;CK�=a_�8e����Dz�Q~ �.L�����({x]lN-���g�9Er�k����ysV�"�}�~"y*�=�M	�H�oHx4<�A�:";-0!�'�gK��n�^B���٢��K�:p]Uˋ҉���&إ�|�.C��圷�ʽ���i�n��?ks-��ڷz�z�YC�.�[(��֋t��:d%_�h]Q6?A�o?��:�_{8FW��V��h '
C
�10�/r�9٥�\�>W"�hnPj�5b�jSͰ���T+g�T$�u��$�40�ʦ�ܝ?Ԉ�H����п�@~���31�]�[U�)l@-�1s���`X(� �[���uZóC/�dID�_��`N�m≪��W�Y�h��sy*CrcE��?'w���be�����e��m��~��h�r6���k�vxm��s�:�ܔ�s5�d(GV{(VA�W�tl�;�m�c�0dDE� �#��\��ш+���5S�p�h
M����֖��2F��V��8�1|��i0��+:����E9f��~�t"�IH��P0lZ�_�FMt;��ٳ`�V�j�̔�k��+�6�P�]9wqv�������T�*�7�A���q�8}{�-�'�����=��Ye�<�C�V�\Ī�}�=|(���&Ф��V1j��Tf�a�Ȑفq�o_Ũ4R��yD O�@�i�p���W�-đD-��a'�DH}���f �ߩ:EC���5R�[��ZKz����rt��^33߭�/����:Ϝ*-�BI�����1�7�F�P��n��C��������]_���]6n��[��Ej�Ƞ_�P��\5�e�*�4O�K;���.����ud�H�	1@bX�L�k� 9�B?��Z���*M��XE_�e�#S^gqۭ4R�q�i�LN2A�U4j��Z:M��+�Yت¼&ꡙȼ����?�/�D���tw�C����Ĕ
?�hE3��.:X0F��������d���J���O��:�$���R���^�����B��C�������ֵ7w��w���5#��F+"+�5Mf�U���{��6�sUV��9��Sz}n7&kCr��Q���¡��߂��b/�=;���Jo�������}^i�1�tC��|�߂5�&"ƁF����� �(1��[Ls�	�Kcm��խ 7LYՒ���v�����f�K�*�������4>k۵�IJ\��[8�Ԥ`溱=A���Ab��S�7ߘ������)B��{�~��:�ҍKⱟ�hn�@,\eL�붰�:,a6ii�M��-	�cH��,���LkB2	�j&���f5�����u�
tީ��$�W�q|y���,ӆsA���H�7��B������M���f�k�ҏ&�r���4��be]}Dcm��u )/�D���wj�m��u����X��4F3�RH�T+JS��;�\��o���Bɤȡ����#�M{PZ'Q�p�˿���\�L�o��x�Rz�[h{@u?:$�E
����M#���av�g\8,˩�'���3�,f���Ec�5���2G�}r��6��p�}���B��N�B���*�7�;�r&M��(o^�v�y��Ź��n����r$)�O?w6�&f6�d�Z3�ܫ������I[˰&�C1�E(R�k7�!�_X�Z%L@�hSJ�נ:%Ι�^����38`�.�Zx��j��p�a� e]�nE�ņ��v=A�\��O��NL�yB�c�x�p^o�Ԩ{SVA�Å���x�{�x4M��oW���Vd�~���c��П�hC��I�ɏ}޴Ec�Ǘ
��p$�3���ZI�`F0UB�ؗ����x��:���|Fj�1ȁic�����!C M�S3�����V<ա���,a-:΋
�;�'KOq/�4nb�bw�������&`���N: �j���Ĉ�ϿX��fw�u��Q���!S��t����j8��4��Ċ�'�D hA�#�,0%!3r�6N8F�Ѝո�@~玲�x�e�%�PS_�<i)�{��aC3Kg�̘�,u�	$��?e=KM�����t��C��o6�����VAb �$\�YT?�5�!��M�W���yޗ��~�jo��	���~4�Xя�2%�O�3�[(��3ό�M"��si8�Ǻ�,�D���u�3_M�d�L`���"3B�F���^��fD�#V�k�n�M�Y��@A�W�X�-�m���*���Ļ��e�ퟅ{�K};�ɜ�帧�
EZb/�&�:��������GSm��].g���α^�?f�:�µ�`ə2g���:��U��`��#?߰55ɧ���$��?)������6@�Ȝ��ۗ$��9B�������!�jt���f������-��h< >P}�a|��<�0���-��^�"Fq�]�5)BWS���in�D�Ntj�mx/������8���u��V�o)���2���o#-tm��y� ��B���	�&�������S�ݔ-T�U��[;aTS�7���dYkj��UFƗO�o�|sV��s�zT��5����4FS�w�N���+���)F}g�.U���"(��dŜ��~$]� <вa���J)V]�@C�\�pj��� l�L(�[�	g��`lf�z,��e��zt\s��b�����qB�w�W�<bHex�EKa
�6�)#��
0�)���߫/&1�24mx�浓n��ޛ����d?JZ/5�P�ӽ�"�C��KYݨ�xD����Y*���#I��m�Y�J	e�q�I���V'G�o��!��eU`�T�*�i�.5w�����3���L�ҵ���inO�[F2i�Ru�Q��@'�N�^��6�^N����B5��m˳��Z�J��D�9R��%	�-� �ۢ��L�Y_w-7@j�2��H8A�`��5f�~���ed�Ys�n��ۧs�gib��+7�ߴ��} �l���e~� �]�N��!�Bs��7��]��F�j�cLz�Y-�aʇ��΄O�����m�fH�ޝ#��1�co��� ]�%O�S2!	�x�O9�aF�t�5&Wg�YU��iKӃg�dTnc �7��ī�{������Y{���G0.&7���t����:z��%)�Y�A�y��;Nk�x���9_�5��R�)���ɫdr���2ڮ��,C/�g+�+�1��!���YL?7��P:��󙶩��2&t＊`vZ}�=�^?A�l�zH��V��t�&\��*�,Boxc�ù��CZ�	&t�3p_��$�[R�0���t��T�A�A�ĭ@S:����}1�� O;����������+Hhs�2�w޻`zp��:�[����JQL��%^���t?E,�D��*/��M�n(zf�b�R�Tb�a���˘��@��+��1�b����^�Dm�A�Z���χ�<��(�U�͕(���hKh�����������MS?ǟQ���-��w��w�;y��3̮�.�<8%G�zW�d���
���ݠChohN4�csGv������Ł�@�������8���xI$`�`��KD|'�4 ^?��N�-�Hגo�ȩ/ђ�s�gy�<v�4�x�o�nuK�㨤��!Iʏ���)�۔mD��è[5d�3)�),�؇I��"�z#�9��f	���D��'Ŏ���8R_ԥ��-䋳�.E��?�5��:H��q����q�>�+6���ڋ`��d�f�(~]���oQ���jy�0��x�(X�ѕK�����e9V��>����1���������[�Ι�g�dM3#
;bz�����Jxu�)����쭪7+>?�cQ񌐄������1i����:���0Y�VMC��~�^L��qb_���wt/9�x�3hi�`�e2�L�U� 7n���k�ꀓ]c���Y�I���i��F)*����ωف�����+�`+�Q/[p7���͒�*F�m�/����L�aԞR��}1�AjD�D��~\2� �0���GJ���36_T�`�x�j������ϊ�Wp��� ���,`5p1��2�B�+'�?x�.;۽��iF���$*_�N������vO��Z��}�����j4h�nIV�dYŲn�5]���$����ߟ�m�d�S�����_g$�g0��AV��BK����B�3������z�X���:�P���+��R��_�D3�����w�����4};�	�m����욇e�h̔��S}n�)�;z�g��������{
���⪆���sr2��v#���K CP
DU#��\'j�Y��_���n�7M�pde{|#���R����(Wt�������T��K�X��3Pd�܁E�B������"�`CGkǧ�h�q�oE�S1o!�T+�{�7;���y�>5z,ak�l+��h�õ�(���W
����)�җ�؆�3I�_\�.�g�����b�ҭ��ɍ����U5��A���{�d"W��i�&n�y�Ж��n�U'�>�I�Gʺ Ծ%��#($ZMk�����1U��;L��]��Qs> �Z��ֱ_�q��s���j�d❑Ӫ�ٿ�'nq�����S��MpEo���&G6�R!�Sl�+�n`�<6��H[��Z������WX���2���x~�[tD0�5[�k���v9Z��QZ��0�l�S,�����^�I-��!P��l��.t���Lf������ѝ.�Q��b�Tn	�q�_�5�9h�v���5 ���\��l�%II��w�k(F=0���zա?���­W�{�����񜴧U9Q�������e=R�By�ˋ�_�zƛ�_Z�*��ܫ'�0�����	�՜ęvA���@��p^M�ʿ�Md�����x-r]��-_X�5��Z��
0�oN9$�!5T�AqS�9y���c ��<փA9�Π��0VZ+D�+O��>v��bv/�*9~=H�$�W���
pA�$�-z��Q:�B*�䝵���nȏU=��b��uH':섰���G� �Z��!��!��S��GIO��3��^	(���g+P�]�l�Wl�CX�DQv�:�w�6�`l��u=���Q�d�w���bo��*	�����`�����{7��Ot.�@]CȜ�����0(�-�o�n���-Cj ~&�.H���:�x���֐5-�UQ�|@�}��^wNE
�c+$�X{GT *��l��9/;6�9v�=��t- ��Z~!�J}�I75Ս}! ��Vp"|.i���g��=��Q��[L!o�^%2�ܚ��)���E��|�L.���Z�x?��}����Mh_�@Ϊ\!� {PՂ����310L+����<�0���q��M(eH
};3�}���>���m%m�mT�������@d0k]��F��W5��J*3{����.�n_�׀�d�~��s����rJW>�l�ҵ"��__3{C��)��ꖔ�O��v_�����) ]��a<���!��oJ�A�t�&*?��9z���g�����}��]�^�r]0}����!�Nb���^�'�W%jq����Xɷ<��+���K�u%Ν}�g����9Fr�{7L����(��3��<9C����/��C+�:����?B;�@-�3�e��OI@�J��Xi�#��.��D�e͉�H7u.>8&�7o<bwg7%+�&X1+�F���o*mEyh��w����iv�f��#��	y)�sGK����~����o4J4��}��\>�c7�)�צ mi�c-�WQ>����K����ne�K�1l��(�px)Z��
��!g�	�`��xZ�݆/�a��j�I[�~l=���]t+�r�۫4M~x�-�����e|���.גq���S�^>�w�	�J���R2�����"#�	���/E���w9�S��Vm��zw��|4�c�����.7�q�P���jmV��*���G{ER6�ܖ\2s��D�����Z ��ө��; �u�/�0���Jt��/(�	���
���@�Tc[A �m�p�� b�Ņ?!������^�V�e�I-tF�;�ǣ��E#�t]����r�Y/��ʙ1c+��vBY����E`Q��A����#|��;��e
!a/d��ʦ����_�B�P���"R�p�Q��U�۲H����{��e��k�ȴ���ɑ߲���|�a�N������ή�Q�^�"q&�j9�S�*<�t��o��+�}l̸����E3�=�L�S�|���L� K�R�X�y��J8jҍ�"i�����{{��|�� *`u\ E�K��
�FL��S*~� ,I<�4S��U7s���9�K?T~�s�P�����I�j��J?%�7�6f���/L��>�ϊ$��>,B�M]Բ��'4��~XsK�F�Hg�p�����;��`Z��PO��/���n��������R��}r-}�L�A�8-�D1����Ļ��ݟ��h(�F,J�`v����O,��=>��&�Fk�r>~�jp�HY�=���k����w�z4��΅��'m����B��<7&��DK��Mp�\7ة���+_q+�Uk�#�.YK��2f��&���Em��Ϟ���1fEP2]+���'C��K~���d}��_���:�f�y������#����_w�EQ*g��z�7��'x��*8^��~��3\���9]�G��if!���?I�������b�C�9Y)�	�"�ʄԒ�n�h����Bc�XK�2�ñ1��?l�Ï�a�G8,F�ͷT	����Qd\+q&w�b��Ȼ�HVd��y�/�6�iM�;p8oTk�h~����XÝ-���ˉ��e%�^ZR�ɉ5��ʢ?\��G�k{L�_��F>�/��㸃w����sL�s��!`��㏀]������W��ߙ���N��X�w.O�n���<5�18*���P:V�G@_J�}q�Y*�ʁ5�n���c�FZ_
���(��KF�����d�R��+Z�+a����ȭ!a�J��VFZ��Y�}���K��#OZ{*&��������ϣ�^�t�㨫!;c��]��-��ӟp*�y��)��&�<����L̕t�Ԃf��l�P/�Yn`WT�Lܶ��&�Rh�?���0V� ���ZL�2a(>+��i�2���-�25�7����o+�bֱ���&Q�
�YU���<��nߊ
rv5��yx�3՞� s�,m�p��U��i�|�t/�[���y��bΊ\�����CZ4����Y�Յ�h���Q/n�����!u�����m���v�.��ם&�PR�T ����n�W�|8s6 �%�pɿ����q)����Eʈ[�d^˖��]��Ȼ6�gUt��k\@K��1B�T��7LBd�� ������Q���
{�����,�܊�m�,��IK�I�)��C̫�ɡvr�0e���߮�]�W7�DZ�c���-,�	��=�N%��� o=���YI�2����E� �e����d	~�Ư�s�+msV��k'�ܭ���e[j���5�=�%����K?,���L�C Ð�gK��iN�P~<��h�ܝ��V_q����AJ~�|`i�VK8B�7���&��1 �:���։�l"ظ����FQ�Wu@�@�����R����˨��\S���Eg�����Э=e�'���}��^4�att8J+;{�8Z���t �:�nv@#��4�-���2�:��h�o $����0��k�egn/ ���������Tzb���9�Ҹ��=E��ݰ<�#���^�B�rꇵ�"���r W���!7�>�yі_�V&֌�OC8^�a.�O ��������,�}<���{�DPq���H�؁�3H�-����
\�q=I1�&$��W�Z��6`���!�}��-��h���-�B�H`=w^��>#��1F�$���
.q5o��t|uH�wMa��|�Y]�/��y;��F9�*��Qv=0.{�8.�M�iX��Szq�h��l/!��|���ne.����_�ɫ�Q���Xݏ
VC}�eFP���V�ߦr�@NR�x�s.���a4���=�+�J�(2��V8Nr�~1�o�^���4<���A�X�A���{)S�u�;"�^�Yp�:�P�	cB���0�v�nm<=R�;+c����5ފ�Ū9,^��N��u�<6D�㯫��#PFW=in/����=auY�9Bk������glȾ��E�6��)�i�ډ��p���r��Xʒcm}fN��U���GC�T��#J�F�^<"pk:�H�d�Ŵ�iV*�Q��hEeD_i��2�LGJ�Z���u��_�M�r��W;YN��9�>B�KJ�!lp{�o'�'������`�� ��
��X�_��nw�ғ5�֖U�D�d�@��[P�;\_O�~����<���n6K��}C3a/���>��&4T�7Rf����}�Z�N��"�0L�6��hZ�B4�,�oS������V���Ɖ2�iR�K�5�R��e�!*����~*X�{a�������L�8��*��VS�ߠ��x\�����mLC�"�8h����]��������#�.?��3=��m`J�$���4�d� �(���?N����T좀?�j�p�A��,s~����V����Ce�)R�
c�{8uKx�KЌ��TV��;(�y8����(X��>�l�{D��\���x{���X�\Qg��-����`�Q���Jy >���4��!�[�w�V��3���Y�EY��L�`W�|J,q���h %#���x����Y^ĲRnӐ�W>_�C��0!&(bM�Ooo�����������عg��J�Rm�(��1?�<��T��bv`"�Zz���49$S�:�]�vm���4M��lF'��~O�fr��gܶ[���~��C�WM�������g�xI�%���@p��v�4�����l��0/̞�=��A"�]�iz�C�����e�v?7Ae�����.k��?�'�K��o�K�J�?B*�le���!N���$��q{g�>�����޾��Ҹ����κC���ʌ�z�ݑ��٬<��9�dqP�}��O��!���δ��#\e/��J}�
Q�ֵ�w�'�*��h�{�0~	E�\E9��[�=�r��8N0 `Ʉ�I�'���W�6]����0f!�5�|/�/Γ�0�P/���ٔO]�X����v�M���.��o*���\�:J��:��Md����Xwy�<�]Y��?+�[�� ��.'��`��fV f>�Z�ekm��/�
�=��8����VZ��Mt6G�e����m��e��}�;M�r�����Jl��^o>��Q`��<ڏ0^ʁ\a���Ӯ�� ��=՟c�U"
7M�^����(�qC6�bE,�8J)De�ja��_��t�f��:+��n=���Rt��cVf�
��(Vl܍s��+�k�Wypq/�4v�E=���K����Ҳn�{�s�b�E]E�}@��\�FR�����3��a#�X��uÐkY�TY ��h����gϔ�p�_��Pk�Q��0����{�	dҳ���C�`mϐY��F�lk��c�:d��k���_���\����AF��h��#��C�����j4���bC	�����aLB��*��,�����!G� S�n"�񽍱>��A�eE��ˬ��hĬo<�lf8o�!g {���W��1�'�K�½9���X�l��g8���ͯrmS-�5ߑf�Ey<��V�o�&DDTm�/�Թ����Hc���[#Ȼ?I��%ڍ.���XGu	�!��������/�~� �uvo�nkx�¡@�h���ʈ�I65|�R�'z��Z�d���T��Z�����{R�F� ?�GHge	�JQр��d�/���U�PofB�+�>�_SS���t0|f��JWVZT����bK��KWfi�����u-���SW�7���֋��*#�_l�b{q^�n6��>�W�͊3�k��1,���֟ �~d���r@���u|q���-C���Th��VA�����E�����+ �}XԨήd��4��r�FL��Lo�Z�"�r;��[d�zȱ���C��{"u<�&9(,Yjt��W�;��l�Ԝ�3}
el���sb�r�(c>֬����\&�q�2\jq4��Q�a臶�-/�v����ମF1�+R}o����렛�l�g��
��o�e�c;^ �9
����\��3�}�׀�X��|X&�,0x�ێߴm0p�ε(�Sy��)y�|��2Jul�k �cҏ/<Ï7PO��>"��rE��w#��0�P�:wZ!~ѳ�^$�~=I*�ݒ�B)� IՀf�>��Y��%8!�����A@�4l�蔆*�b� �ӗ��畎��m2�`������Eɠ'��$5��X4�0�������=>����
�(����^��6�:����-�ȂBaU�6cw����R��#��ȷ�;�`笀�c��eU���r�
��4I�.�Ě�Y�Lq��d�4�a��<��a��?��m(���c�{�`c�А��b���'#��p�2�õqNc�pQ��d�*@%�������K����i��V̎���
V�*,Ž�������Di0t�9֖0�=yJ�3[�K\�����Z�-�dWλ&���J5!ۨ����D���l_��;�Q<3y&�!�l�r�|3�q�1�Z)X� �Ʃ��ї��C4�$E�J`$_,�$�&�</�ʱ������JC�AZ��^��].���J�+[;V_8�2���I�{d����:�|34� ���&O�{7�'����԰9PB�ȄƼlY����K�<�ꑜ��M'���%3�\��b�l�:b��L�#����9���>��N+7�T�6�(���к��8+�3 �s�^L����8��k���l�}��r�٨�C����SC+�4W�����H�nd�!\q�XǊ�Ƃ�IxY���&iOPj�SUU����Y�`��&��n��Ɇ��h�+lL�����pV����c�ZQ�WA�UuV#�+V	�9�I� ���.�e��fS���\�%���es����w*u*�r)��/�<�,9�8^��ܵw��S��yMk��3qj��
��E",V��<]e;;U#�ڤ�C2�/�.C�=�_����W`8���_�>Gkx�����%���}�3\]�ۥ/
�b�}�.a�s�_p�g��&�]�u���Kg	l��7�����,��Z��O)<��㧤�`Q0��iJ�
O��x�'��H�X�U/+�.�~q���K�w�� ���Bܛ�$m�T��q�|fD{(���'4Y�g��ks���)�K�T��]��.T�׋�{%wհ�kmfv5�x R��Z�g����3�島r����H�ĵ��gV�`�!�����@��:~~��k;@V���\���c���>���5tN�kZ�d_-C'}C��W�r�0`ⳆUA���+���8����6	�N�`T8O3HAlB��\~��'��Ӡ׬b'�^2�{���"�0i�bl�	�yS<m�&��!� �"H$Q<7h�����~�}=�)��ߘx76�,|�xm���z=����=bQ4s0��a��M�A��Uy4E)�˻&܏����H��wz�ily�j��Vx;����G�
�:�k��Ο�����-B�.#�dؚ�V�pXe�_st�뉻���T�I^5:��3�{a�����~���>-�t��~��#�{��Vudf% ?��#������T&�R�si�ݒͬ�v�U�E��goJvɟXTۿ�m�P&�C�oV������a��:;x���`�{�ᝯ5wC��T*;m��|�_F��Rj1�}/̈́ڬC\�;����eh6���x9+��iɢi%Z�%i�֕��\���k�P�Y���c�+-Ѓ�ֶǿ�!�:]u���G��q�/�'EZZٕ���.��㹂˜LD�`N�阙�c����g��&�~���ֈZ�Ө��9g�
�',���{�p��(�� ���E�7�c�z���"y?x&y�	.�68�9�=v���?	�ӓ����?��I4ś�1[?��W�1�"�}��~ur�����H�0��K�(*b{��6�8����������F�0��v�G�X ���Ú�Gކ�,�^����ʱ'Ҳ;iG����ܹH�ͪ���fV��87%6Ne\�Ox΍q�K�%��>\�\$�����8��>ox��N�zȝ���"��g8��POե�z{ȏ
wڎ�x,��@M��s7Cy�x����g�g�Χ�-u�GZ�@נ�0f�|�����x��-��d������`��:��	��Dx�ïv�n׶4�'�6��֐Zƾ͊��{��=0<e?f;��'��	9���e �D�&(�i.�JZ�Iܙ$����T�׺��~�=%c�����.O�� t�F���i�5,��7����1���g4��5�(>����.*X�Y!��5�,~�Rc�Bqs�e��	�F;x�{�4�x(˭~$ܞ�Vǵj�c7Y�����ȓ�����1�n{����*`E)J�v������T�.��P/��'��?��x�G�k�RM����y�� [���`v�ϱUg��)#����yY
�b� �� ��R���-kֈ&�@�`Ŀ��8R�#'�gJ�P> ��2��.�΃����ρz���W5�(��4���T���o,b�����![����)|2ym�Q���,�f+��gk!�o$�`�8V���1�u�}�����\���q�ɾE���:D ���"��)�i&F�/F�|'H��͓B{��+O���l���Ñ@m7Dp����٘p/�3���`���Y�"�"��m�
�
�1v��|"s�k���%"��4u܏x��p�
zCu�ܑ�.e�~�5�dE�@D[���V��m~.�O�xK�s�=ab/��ݿ9^�<�G���8A��P�"�Љ.��[�Q�x���!TW���9VHHJ�g6X(-�ktKb�S1jN�))CGE~�'W�.�Z�ܵ*���fSV�)�; ?���^�Ǜz]�}�p�R�QE!ai�h�~d�pR�(��f���Y�i1����/��
W������8�{D���pP5Dҵ�f����"æ�����F �9 ��|�����j>Dn�^�����
@���Z��(���wk���bG�?��@�W[ۯ�l��U
De�cZ1��Q�`�'Ū��Cc��I#���m7�P 8�b^;�Qb��JD|������?��J���ɖg�B<�fXZq��Iz;=ci��N@���o���VDQ�yɒ�C��.��麄�*��c���@�#4�7ف���a����@H�nBݏ�Loè�a�;w�2��
��(�}�@]Rd�J͆�˩u �Y~C��J�*��yiI��h��&^��$F�d$��υ�Q��X�s��a?eb�D��Z� �ol�ND������n�g3���I�MH�Q�����|��I��G�������iէy��C'�j�W�Q��XmW��ɑ�ۤ���<XXl�1�q_�x����T���A�!��-�37#����z��Gљ��;�a�k�QY_��9g��M59�9X$aq�h*�z�o���=_�;_��IZ{�o�[l�$�ᢛ���	^n���@����A���3�I/E��$��]�:%��[�*�D�?�:s����-�t��q����1��N���ҏ���\(�?W�/ʎ�P\�; ){Ԭ�~�kٲe�9; �aC�EQ�W�?�,�e���Bg�n5K%l����Q�]�����m-٧�3���`V��(ͿEJ���0�Oj�ψ�#mtr�P��N�ՆM�@f���aR� JA�u<�
�Sy�'O	k�:��:i��ˢ�WcI�_v�Jq�����X}��pV�O�HT)=�S��dg~aҪ&�55�c����)3P��XC�� �${��d'{��ǒ,#�EW�����0�RT���Q=5.it?�@X4b�ݺ������p�'�?g�ce#��vF)	ʒ�+5K#7��j��՚��W+@ZQ���{M���������a��Ƥ���Mc�f����3؈}���F<�s zc��q<?�
H8}+J���l6���$�|%��`!��Ռ�nn��Pw���^ ��Vg�x�Q�u�q�c�@3#�Y�8:Yo_I ����n "�\hL�E�#[9z2|Q��Uq)w���1�S��
�$Tq�@ʹ�����pcN�XV��03��V�P��Os������q��F��|;�<8��Hͳ�(��wmՓ�Q�]�mtyLth�kf!D�=~&���G�	����ߒk�2=Ў���7P1 b	�bL�R`xq�|����dW�Y�����-�?g�����ZC3�a�vU��_G�� U>���j8p]봸�VM��va$��N��dL:%L�P�(?@��5m�N��z�8�?Ql)�	/rCuC��d(�+J�]�Z->?��Y�8����b�Gl����|�m:���I�]XP�� �ئ��_���A@�śT�/icĜ`�Op�J��ˍ�,��q�1� 2�h�WHݼ�ah^��OU�x�t)L�O��v�����DQ{$�Z�hDܑ����ᯅP�?]�l3��
��Z�`0���a�:r�t�3��0�{T>&c-�%�,śbF���Y4�����p��F$�D��GB��/�������jY��r�+����A:+�B2����X�� P#8�ҋ��l+lǧr�rᬘ��n�[�f�5��S��X
!u�	�,��6�=�\٘ o��h�
�4��.�G�(�:x�b�w�~��{�]�~VP���\�A��.>����|[wf�=b�<%V�h@������#)qw����
�˨�SU	�E6~������[W�F��Q����'� w�,�s� ����p���u���M�jɲBP��$tGB�����z]��jA#����XN���<��SǼ]��C7�g�� ���Kx�eD�!h�3oW8��_���ƅ�A��OUTM���u��e�%�m�V�Lltm��{���^�����<�,>ߣ�}Y��>�(�:�x}q�T�ߵ��*�[2�o��2s��!��ʵlձ��H{����I�-X��<�ڭ�j͈>m��+>��C�z����'��\���i�v�F+�M�r̝�s?'zl�|��#f�b�g�N&���j�=���)b2��\����W+��E&m��r��i�<�O�$�9��E��l7hƩ$XV�`�o�(�;��B�\%�r�̉�G7L;�L�ݔHC�tK���ɑ��h��$>߶��Z�*۫�2�G	�b��b;��IAfTU��X �
�<O��2�ɚ�2�FZ}m�#�Y%D�`&7��a�Z�_�M�" s���B�4Nޒ�!��j88&>���{��y�� �4mB�u���j�IWG�u�ؚ?�bo}���K�Rz��Qj9'2tb����H/Wl�^��U�	�纀��k��ڎg���!�j����{C'���>I�Q���A�?d!���gs����Z���d����*�- n��}z�;K�ﵗC����
(��UGj�k�6�wwR�&S�X
eekI�����r�ҏG�D1mq��ٖ���u�go �½|n�������wS;큆��+�\<��ٽ��%=� W'�y)��fb�4AǬ{�V�B����g�e>����d��|L�����<��F��9��E�ZR�t8�e��V	k��lʊe�̓K*�{�.��Sx%KL
�f�̡���qǱ��`��;_s3�:��y,��1ؿ�1�Q$.9��x5q�&�St�*{2Ѽ���`bo�DcA��Ơ�%@�vq�����a07����a@����K
u6��Y��<��q����O`�iӂ�tA��ˤ
i��q�B������-�@���F>�R[�%�_�e��#�]&f�D���%��shԹȸ�3I��ӈ0ǁ.�b\�����'Y�mH��"`�Ǡo�C�vé�w!~T���]jMG)0͜BbM�*��`m�5��5���2����@��5���# �̝F�q���ߍ�f1��C��W%�C��znhlVN`�Z��<n����i&)m�d�>u�O��`�N�w_"���y�yNq�8�R���By
tU�$�H�e�9��
��jifq�4~4hv��Q֡o�S�!vb�|G��&�����f�0J�u��s��Q�uIQw�j���}��.�]XdJ�KdGv�g��Q^�7(������x����n��	O9�����A)mNv�s�[�S����Q��ڒ��_#-��6��Yʵ�pA�̹|5�s��wm���e�(4G���݌(�Uv�_�[������%d�H�b^��$����yhx�3#��>1�g5�l�Z��#+�6�~���Dɇcg��Ŭ)�t;
o	�F�87	����vp�ZA$��3Z���?j���e�t�@�ɭ��]���D Bi C��$�=J�Qv�� Ό?~
��^N���;y��iI���#)m-W<>?'��.Q�嗪��E�^����D6���JIƒ5xA� ��;�|E��b��7Ϡ�CZI�(�K B�	Vn�黵M(���H���*Ʒw��0�u��I�ذ��]!b���m/��� �O��Tx*
��΄�;,����C�4�FmCL�2�,���Q�7�S<��چ���bY���I1˞�}[����`�!�]�8��/U6���+<N�p����\L�k"^#��!m���e�H�d�����T�n�&�L"����<���'�/�O�1�Tx3�۪��-������fm�EO@@�ȥ�觊�&X��9���˧��4�X��%B�5q�� [�.R��zEx����*��r�����_
�9O�֪���͗�T��Ǌ���C��F%��쬬��Z�>(�D;~�L�����k#��.6-t;����w��v���� A�@��<<��,@�XQ:0�Z��)A7ߞ>M-� ��KO?�𲧹 �'�j�@1,�se��>�!��y�G핯��y�Ĭ�{��֋ǭs_
��a/�a|�CF��n/��v�K<����>#�{x�=�r6���(	v��Ր7_e9׋�3m�iK��JxYɓ�+��k3-!A-���؊]�'ߋP%/!�@��5��?ي;�
0#���M_{H�a��9���o`�4Iy�.�~��Z(b'�V��C<�`�S�����Tv�T�C��R6ì��ohw�dK��"7���n�^��H��>��8��ζ@3z�!,5~d61�"���>%)mcζ ��(0R�{CW^귐|�o�\�E����\Z"t��b�+IG+�")�Em�̈́��i�Ʒ��>�Td6�a�}Xv���l�6�j���Xͪ����.�~�6#L��ܻ�0��ej���f�`���'N�btu�n����vͺ!I�i'�4@��Vk�AU���zrުm"�[!�;`ˆRF�%�-\Q����O�_�3��^��\6W1wv�sq��xM�S�p�z�L�O�$�6�$/e䈡�A�x%�(�5N،�X������DJ�j��8�*XR�����RE�;�Bdg��,��S1_HÀI��6�E��ʽߚX�7T����8��Q�m3�Mu5ｉ�sd�f7+i�񛱐��ƅ�=z:��Xjk�,���
�LqԙI��H�j�B!\^ϫJ0�eo�<�dg�>ga�7|�
Z���x�<j,�f�PE�b�J�.�No� sc:��n���0��i��3ժ�K���W���}~L� ��5�n�c*��7|r����jb��Jџ��9
C�*I���0��Jl���=�2��ٕ"݅��� ��/P�|�5a@!�t����v�֌��+	�V�Yu��m~?�,��>\!i^�t�B]��Ɯxwzy�~n���§OpUBP@4�v�5�1�I��dJE[��mN�}Kg��w�sR�1xu�������8�{��K���<�ɸDR �0̬�ʓ�J�nf�����s��8�]L��cV��U,��jkʀ�/	���o2#�b�Zs����"�}<rk������"=���Q�F��/$�j�J�wP���L'�PBѠ�8��%��s�F�j��CAj޽�-Q[}[Fǉ�G�z��V·��}9$u�������r���*� �����M��6,����N4D�H�N��-s�HI՟��h�0�����T$s�>]��jG&�v�Q��������U��{:�a�!y}����|�D���_��Ŋ^�|0	��7�:՗����)����Yy�s�+� �:���$5�.ݖS�|�l�<Ka$���@g�x2�������y��^�K %Fo��c�ׁ+x�.�1z0���n�~��m�;��
Y�Ȧ@7s���O�
�����n�$*�#��!�g����0��nħQ�pl�	���Q�aG!�8���hMh���Lo��n��FY�g����R��7'q�q%�$��/���p�0E��uឮ6��2�C_I�W�+A d4: ܿA�h�gvźᝊ!r���	,�,Nj�x��\3�\�:�U�5�h��s�&bp���Sh�zy�p��+Q��Ic]3�"�#�K�������~��uA{q��2�A������˕�$#�H�D@P�>�	Rn,����t��]=���MЭ��6�݂���r�T��t��tgԩ�n6Þ<��5�Y�r+�c���#��f�',������uG��Ә<w0���� Ӿ����%��	)�
�]�"ܷga,�b�!C�cof���E�b%�J�#�-s8)�Ql�Ĉ�H9zW��@�O�
�T���Q��a��EE���8�i��RL�ܺ��ݑ���=W}G �1�|�#D�u�KX[��^_�Q+�%K���� m�p�3��^����V�B�g�s���n>)cS�à�g�#�+�1����B
>IV�E�㰦�o�6��9�%����QFO]����������ؓAM�󩒖nM>2�*�&B��jq�߂�z��l*�N�����f�FF�<Fk�'�Y.s��sr��c2���*�N`OT�M�xCD}��?��W;��&^:���e�RĆ��D��IC��\N�_��-�k������ć�x��s_�j䉮���NyI���-*�m��5NW@<�9��B�6�Pߠ��g{1�c����\=ꛯ/�)>��9Lۃ��tʫ�n���:������Ӽv6�;0	�i#�v3�&��������f�
آc��1j�;$AY�)Iu�i���P@m7#������6�m�9'�x,�v˙�@O�g��4�I��(�$���K�U���h�\�c�#�b�o����y�z�xb��㔀��=/(T<N�'s>�w�cL��߀����g��h�P����D�*�#;�|V�t�m��O���L�$G�IYtaK/��(�`��3�MF�ǦN��Kh��T�3�"n�Dp=��MǷQdC^s�>m��>#T�x�u��jε���koӮ�'���c�(Ù���"H�Pk�L��?� ��\)�V�u~�������.m#���F��,�, m���\K�0�69Hs�s�+L�降C��[AW�w+�\�O�����$��%�k��#[0R�j���8w���?�L�	���k	FdI
�l������	�CS������/��B��9��(���<;�x���W����u��� Juuƍ���o�dnxe.?X���v���U!l��7�����p:�NLڜ=>�7d����s��k�4�Sy���d��a2 GO+��
XjS��=E䪎^�G���[��vo�cH^�X��`|��8e�t�R�wU��i�X6s�����S:A��j�.e���2$��F�}jiam|�Ϳ%���*��ҁ�l�]�hL�-�hs6��9U��󷌪��W�9�v �Qh\?PJ�تe���Q���w'v�45�L��<��ǋvA�<��0�|F��Tjr��a�:�
I�ڈB�'Hjrb��[��#�<�����|g��o��ٳH8�ݶϨ<��B���ih�]>a�ۢkË'�v^���]�
%��j�3���E�[��R��	n��Uc��*�K�e�8��J�t��̙�5�g�$�/^C	�. ɘW	Q�jx6����<b0����?H����2��߳6�EC������w<���E��c���I��S����f��4J��;!��U��O��jj��R�}tuޥ�A���g*��4�~��qol��]3�����%�3����k��^����{'<|ݗo�XM���M���P@�.�h�s/�7�Jb� ;"�2l��X$���f*�M�c��㜶��bb�"�rb��)�!�Uv�*�¤z�c�����v��nmؘjL��ȏc���=�(�V%-	���^F�n�D�;3��6�=Vu��"Έ�|�*��t�*���cn����,�{7����9�*T��j������\荂焍�ԓ��c/!�O5Ę}ڎF���ǖ8>6y����	� �{��`����ܷ��s��nT�&���m�_�Ѡ�E}(�E�Ie��7�|;=^�I����H�'�k<ò��g/@�_:��).,"(��6sm��I�m1��Ue�ڳ*�&���yL�)��Z��C��u��CPd���r�M�E��.�@�y�p�}z��j�.�-���Qse'J�@t��?Z9M"�=y���>��W�
�4)�9^�d��Z?3��]�]�D� Z���(�l~r��Ƃ:��W��BX���#�o����L�b�����c2��ڐ�ԣ��K�ʤ��3̻g�dQ��pZ<P�ζS�fI䚏�e ���="�**�ı (�rd�D��d�vHH�{u&����[
��.�� D��=�<���j$}��TU����#)*o��ɗ�B�yQ����z�K,k�Y�cwb���i��.*xȯ���Q�ZOU3�;p�v��9�0_�m����؜����c#��)_ţ�U�{l�c�L�	�1����DHQ���Z��yAp�[���۴�a 1Lv�t��"����ZwM�hSF�	�%VФZ�5#G��j��h�l�n����_J����h��Ӵ?��6�i��V��yZ�����"-m��٧�uF�(o�̉Z^��A�B���L*�r��?����	����43�S�MF4�֗]W�i�վI�Ĥ�����!�-�|���]���8��8���e�FJ犼�ha�O:�B�\�\�$2�u����{5R��K��S��f�9V`��q*"Y��pΪH�'�ņ�)�����F�7�1cr(a� ��5H�*��';�#g�W0�P��B��yj��0��|��3��QB�dH��7R�j�����ӄqW=�
��W�L�gj}J��s�FofցF�Z�QYy[HJ��& �t.D�O+��r����UcMziY�;	.Fr��{OΞ���u����ZG����� t�Z;z2b&�,����g�������=��(�;՚�@b�fL9\/pj�X�c�ڴ�k	���p�;���LT͊����fY�w8Ń�`;�/��om5l~��L�p�D�o�Q�ʓ�<-�Rd��[�*���O<���q������)����9.7,����%�mC�bO�F(�%���2���C_��7l����^���H���hm^�$Y�p����ɦz{*�K�� 9�f�v����9w��XҬ�Ⱥ�T�Dw���2i�t��ʙ���ϐ���f=1�w�WfG(��2���-F��s�f�_����U�!
��X7�!������ٹ�G��k�K�F�N8�̓M^0-�F�t�e˿���`g2f�Z��*��c��vLv۾G�%~���*yk�E�^=��&(e�o�<y�"�\K=>vэ�O� �
hm��1X�[�b�c�[��r��E�_�g��oH)�Y��ty�e�CEv7pu�U�5�{Ct N�_��sP{{xs����w���A$J��An�����G���w ��4ϐ��zsf���Į� �r}h]���7#HK+��l�b�f>ϙ�n~�ıdE�L���`k�>��ѹ�%l��u''���~�<a P���[&{�6��͗;�'�+�AG�k*U��_��=�}���3���{��嘹�#2]��4��$#� �̔�EG��Hs9bF^��a�`���$���˕�\�|D����57�v?�}�->=��J����E�Y �P2p��z�$WmGJF7�O����~�?� �Nk�x�%Eی�&<��E���<+�x��۪��,�S)E��t	ֽ��/�>IlY"�V�ܑ�r�)����o. �?��qۛ3Y�e;M0ŝ��F!y0�YC�U�#_�������i�JM�;��J2u S���OX���=�h���V��e�i��S���K?�;Z�t��,0�/��_g�����|�Xy��t��Q=��)v�t�PE���bO��ٸ6e��%v��iQ��yߒ�����S}*�/Ę��fH
�=�RΘ;�''ҍ�������(� 9��A[�:cŌ^N5
L������ʘ�\5��\�x��.�d(�tm��8K
�W�jv{�n���g�w�c"�����`ؙB�l
���E}���Z.-�(���%�_u�fc��&�j�	�hX�F����m�s>���z�]�����ƺ��TN@�mWwX�s�d(������`��H��V�HO_#���F��I���9��((T��Q,Git�f����Ǽ�C2�(7�+͢�'M����і?!�!m�to�DD���߿��$�ݶ�t~�t���3E�K�3���<#ߒ�+&Y��[��^ё�0�˪x���!v�[K4��*�_R�?�K?@�ϊz�i��7�L�S�S,���vD�����d��c��0�v=����C���&�-op����@,�5����3�ļ��cān��Hc����B��L�4�`����g���S����6�hFvx����c��#�}���c��뱗�0��y6H	��_V3˲�!'��T��џi���a��x�J��.���VLv:��q���{�2��2��}Ipa��u*9(W�w���L�ހh���N�Z��O�q��s���=L�3e�^�S�2�)���3s����:�
��r�i7�:�xn����0Y��K���Q��&��3�5�E�f�s�	@�&����w���6&�/����fc ^����m�H����o_|R��)�E��Т�S-s)����K��^!A��f���V��GH�%|���ʚg�ķ@j�K�>B�RG�c�ވ�sşrϖӠ#�Ô�|�<�����T���;��9u1�`���ɬ�O��cF1o��}�#Kػ}���G�H$\��XM���}��9�J!	�z�2y�����HQтV���~-Y#C��cӤqV4��	۔`�R>L`��ǧ_�X>W~g	L����"�����,���*¯�3���j+���|O%�4�C1U?�B8M�K��Ů�m9V��_�6{-��S�Z�>������VF%8c���U�@KCd����KWK�!��^�D@P��w�C5���v�����&��;m��8�R��Ƴ�QN.7=y-+�F6�>����O۟C���"f��$�0�@��S�8��(��,+_��ͯ����c:�+S�Μ0��p�Gq�9|���e�~��L+؄���Q�0���Խ���asd��R#� �'�	����!v���M4����7�Ǯ�Ӻ���G��O`o{�V"�p=��L�(z�O��ةbf�I������Н�����p�FU-Z��SxaX�i�Ȗ��H�ۺG���RC��4���c��g��O�W�m��_���ZsQdFgk�U)�x���+��BPr�Vɤac�� �O�>��Q}H���2r' ʷ~:���;�`h�ݭfZ��u
\K�F�g<��ˊ�F�ύ�zdR]�F�G�{��fD��â�rP>�(��L�#G�/]�5�҄m��t�~s��ۑ��~�nm9�=Xt�S}�Zv�E�����A�Y}��� UOX�j=z�2�����@ە�g��]��Q���n���ޤ�3.sN)R����*�����P�QJ�m�_j3Ǻh)Sz�<�S�NɽJ/,����p�uQ�	V��`Pc_R����Q�G��^C���������VP8���+dC6~f���"�~b���RJ_`hڝ�f�(PH��q�Z�P�Q�-��Ƨ�ZF���G���1&�4Ԙ���;]y�7��{@\�jr&s��ߑD �`�%�e�D9[u3p��(�x���d{��厈���i'���ғ�Vоs�������̰��'y�Td�KW�^����w,��E�{��m���ylj�m�4�?ǫ���Q�8J*r�n�v���d���:�$]JO�<��;O�v�vd��C-��,d�B�ś�9��0R�SS)>HD�>���,.^-<��$�ЎI�%�ٍ��2���y���9A,���Bg#�UAk��d���]@�Aǘ��ľ޺��ڋ��ߥ��?+-�#׿��l��S�$eOV���ޅ����A)���b	|�Z,�pw�i{�ϢeU%0j9@�:Bs-`�N�$M���V�D �s��#]�w֒D����~I���P	��e��C��v��J��7�Sj�y�*��՝[�ܴ����k�������Kf˦ ��Ae.X�DA��ݸ��O5�����
��u1	�rIf;�xB����ڞ�41~���<�	.Q5y4�f�=~�kmYH���ȑ�a,?�Ajd������/[�Ũ�f�|jI��V��멠��њ����u��\zܖE[�hyv�"�Ӓ����w� �.������|��D$�t�y�l�t�@A�f ��!�¥A����������i0�f�*�5K��,%H��0�<4X���BL���N"��������B:�ŏH3㌿�Ȥ�S�yi�W%��T$YXhH�9L�LΘ�<S�������um��h��"R� ���yTW�:���R+�$M�u�����)Z�n�y��*�d��h���q��O�ܐ��$�~��>���x@�Ԃ������n�� v^.4e�%��O�`��9�#\]��d�qk��5QT��=�����`�)(�~S��y�=\g:f��9,�8�ׂ�W�,���ht��}���{����e	�����?S+GM[�N�5���Q%y���.���,����
O��C?�u�}k�N�7�bi_�4_��H�t���K��mW�m6�E�Nj��B"��S�Qr0Kȧ����t�[gY���㭣�#�K�hK�~-xL�����A���Ĩ��Aa���社V���m�?�c�i�D�N����.Х��2+�r(�*H��2kW�!ZkP�����2�Hg�-�Ǹ�
-�IP�*�A��+�̸��&�HXfBkv���(����l�1z�5i}���2��@�a�F V�鹜]'��U��>�E���8�z�2UEA&X�%]7��G���a~�� �SU�)�Byє�ye]z��fЫ�6/����)�r���U�Ꮋ-JZE�B�5k���0,���g�H����q����׭�pe�9���D�8J(�Ɛ�����:���)l�.�VJ`G@�3���(5Y�sR��"���M��Ö�u
�:ׁ��;�8<X�4�sr`*S�bϝ�ё�[ !���l�� ܍��L4	;��3pHEv4�?�,�RS3$I���9�س�E	v呢���{�L�QߍQ&m �6Y�e�%��.8s�٫tI�ٓ��x�2TDp<�c*�x�hQ��Q���4�����q0�K!��v���`(��M�^c"A-�x���땊=�1x��`C�m~�9��=�����̜k��a[���~R\\N���+	FF�C�)�D�>��n%o��+anm=R�6m^*�`K���Ǖ�H.�z�ڇ��G`�Z��v\�;���Ɏ��"Yǚ�B��6����ZЃ��Z���������u����J P�j�&[����j��wcWC���П�VI`�sTr�Ӭw�eűk��/iEN�b�Q'K�V	&pV������(�p�)�D@�4G��uy�UF��)-�����T��,i��󞣔����}�2&i�-�qi�b�-�;�E.��ߚ�c�d��� wÿ��������T���N��h���1�����O�w$�V���ܟx\����}J�I0��N�h�'���Yixʣ�SO0yRl�RM�i�1�)��G��~DHDݟ�vnip3�Aj͵���k�z�j�Ѫ�7�>�2Q>0�e�Ͷd�w������0q�j�~�"�ȶ����t?���A��r�Iz�3ve��ǌ!�経o%��5��9S�Q����K+e���Ccb���69�n��d@��-�ˀzEǑִ�
Q��]�hzJ���6�z�^�}q�%3Q6VN�鬌�\ ��zȦ�F˕DX���7�?ii�r��x�3j۠$V�
���eS!�l��2Y�X!�Zo
:���0Z��j�<�p%��d���A��&��i��/�j���}�Ђ��o0��`����6���[�o�!>^���$ZP�͛h�b���!�j����j���A6�m�2~u�x��Cuz�3e$�����u�P����Z�ⓢ�<�pV#Z�2"e����D�&n�Vtt��E_9J.��*��Wڂ�<�����;��]奷b�QUG��.���Q�,ذĞt��ҷ#�x3�i��)�G��|n�J,h��G��)yVZ�7?o���Z�_�����õ�dҏ�,���Qn0�:mj���F����s��7`���(�9`o_�.7!�{!�p���Ra�N�-> �f;�8������QT*�o"��Հ�ni�1;`��$���~�a�C`�	�_����w���'�Z_�u-�d��0f�j�5��Q�{Җ�����V&�#�5��K�8�%�դ��w����Ac��[I��Z���X"Qdf4�p���;qL�}��/�'��tB`	R���&���$j�Pn,cXX���"�>ѐ0u�=���)�ד� f�Q�_o�
\7�}���^b����!�;��U����{�Т���}�{b�%��},ݮ�X�b�l�v��o�qxs�[x%���u:��V%9��cd�,X�Q�r`��� �&<���#��:�@��2���F�R�BK=_�R�nm�Õ�K=���2M���9�A��=S������{�^c���8������n�rqe#�K����U��y��\�R���J�;��um>e���s�����f�/ð�}�����(NpY	`�Z�;u9�b$��Iڙ�K6f����e3�u��q������ޞ�@	xɱzq�
d�Ht�qÐE�H�/��yJ@%~]���y)BK���#�M��)�;��^����������`1B(����{���L"��B�8{ E���� h0J��o�8f?0s��� �ڡ����yD��"��K�A;j)xcKo��pj#�g��֭~��5�C%ߐBM�����:�	�F�E��P��Q~Ӭz4O%�I]{�0�H}Z�O�m�eaq���v� �x�[�}A��dM����/�/m�7m�2yjy�����iSxp�PLu�[�7�@F�j��K�+�����7�3S����̽�_���n��N�{�#A=�`#E�Z�$pr~��,��J}"�D:I#���*��x:fT��C);�zk+����~�d�u�>,x����j���4�!D����4�����,�?�'��>I�
)��lj+����I}�OH�D 핏(����Ȏ�A��O΍�n�10tץ8?�FGDg��dV�YU��(��?{�Z6Ἱ��?�����3Pd��q��T.���W����ė���(U�����!������w�E�8L�q��櫗w}�`jh;([���0���FM�٩{~�{�^+�4UE��V�v��=�}:xu��[��?����cl���T0�ѓlڑ	���R��	e�cY�zV�>}FH�$���%��9l�"�?�CP�B���>�1D~���Jp�M�FK֟Xq�w0�m?���U9�ai1+��9�VH�*�ǌ|�R�w�f}Vn�7�eI~���^�%T,"ZfJ#���a~��|O�����m0��\:E �בS�d�������=Z�qΖ����l�;�����o#�Ҙ�S{�PY���.f���b�"9����g���P��ˈf�́m�$R�8���j�yw'����"���-[���	q�@l�T��]��Њh%����`8��u�w�JX!3�O�l�,����q�P�W��N�����}�¾c@��K�����i�y�<{�*�W��~��Q��3ߜ���M��h
*�pT5jc8��:�N.w��eK26A�l$~j���vf����P��d}L"Ly���fB��著�P{��㛴��	uY��udۄ�m܍��@�I$*~��JL#L�'Iˡ:!+��bz���'���L]b*6�E`��Z:MD(p�����8���hp�#���S�=�p8����5�����m�@}05��AOHnJI~��T��5pg�x�U�\X?�P�&Ix"d��+l�v�|�\/጖����#���X��� m��M�-B��â7���Q���z{b�b2\R:�bv5C]-	;�K�Z
�LӠ%p���TUݗ� ��?��a�$bQ]�����K�Z_��`�� ��ҏa�c�����8oa������8Z���}Y1�%8,���bß�D.9�y\^,m�C-�A�=�"�2�����?�EY�a�H��G���Ӏ�$���۩��4�C�J.�C���������Jn�!WnͶ�6�=Y���ʪ�N�m��~����Z�s+��#�uUuev�RxKF��Q�	t�A��.���t���;����\J����u�������q���Cb4���Yl�Nij���2��Y�)��x����te�'�?k����/Wj:9�Z��b����Y�{�� J*��KAb����MM�M�B�=�f� ��⚹抩*QcS΁�b���F��rG����
3���I�gq���3ۋ�ng�=���jOj�v>��U����
�4�{H�l�q�ŗ+9�迈�=g+���j`:�D
7n��k�#:��j�Ox]j���s�V�����Z _6ѫW��+�#�|�WFs�����Qq��h��)��,�eig��YD�W��ey�v��Ȩ�6vQ�(FGj�qH�:e�D��E��귛����d���[%������I��a���TY{þ�Ʋ��p��I?�~�����~ =�����&�;W� ���{�I���nQ0�,L���cg���2`���PH�4,q�9�AW��|�@�99g��U�B�.4�7��1�3�@�ۓS��)��={����A�2�� �'p#U̻hYH\V5+������	���BE+���e
H\��#p�������������r�2��t�d��R�L�[s�;�ee��ߛ���'v��F~�A+sx����Jd�A����C]�2?�t�񮴠�Fpxp���,��B�F�(W�'.+��d�g�!�`8�� ��k�Z����2�H~?�65%!��%K�`�[����ע|A,�<:�R_.ߜk9	]��F�1���r�N}��j�oF��LlS��g���)�w�����v�	4��p�f�	�������$]H~l6�2+��p���y�?��ŭ����t�I�����S��P����.ˍ��Ex��X����yj'��0l�À�����,��~�5�ˡ�aЖK��9�Nq��)ɶ�(:����j۩�M�Uw��B}�F�U���	�V[D)�HL�n}�*f���NJ	dD����Tc<�(�>I����|P��K��t!tSQ�> �u��jÞ��7P�ã�8�}b��k*���gY����L�Č�.�z��O�n�Y��aLa?��G_#��V�9=��W��N$�5�)M����Nひ(� y�D?�Zµ1��<؛ r�m�-��U6��%�lb�^sh�u|P��ڠ��g�R*R��H��|��gװ䛩��{���̈4gNș: y�j$����'@Z�G��͂�KF�ޞ�*A	9�?��B�^����ծ�k(b�cRP-��q2���1����rF��{Lt��0��5y|P�xyu�u�L萞�P(#� fB̊�T�N�Q@����m�*��މ��=�mRX��s��F&�+�:A�Dg�_���8�+=�j�7B�9�C�.0{f�{�����N�5��ԋ%�*T,��c�N&�)"��w������v�1:@�%i����[p���J^TgD�-���Z��jx��sf�t�ܔx�w�A����-�?T�%�(yԚ0S.��c""�mv��V&��M)�Y+�q�Af����e|�����/�%o~·T���q� �����D�I��.�ʔ��0���X��)�7�2#��3L~�jcE�T�z>/�=��e�W/�=
�V��Ҵ��KC�T1�=��1IeD�d����z>a�f������Ǒ��o1��A?U�z�OŜ[�yroS���ZL��8����R{p�/�i��e��L8�}hQ=��*Y�wh.�*Yֽ�|ҟV��ci��3��k�K�.d���9U������i݉�0����&�`(��R�ޑ!�c��z�xv��K{S�\��a�a�,��� ��o:X������#�e7���O�K?םnr��n��59�v��7V�3О{.ࠇ0��j3{GWe�X7��S��9��*�RJ��v?���	��KPI��-�@�nE6�.��Ur�I#z3��b���c{��3&��4]C|��W���E�۸�'�#a�h-/��&������@���+t���h)�;͓���"�_�	w���2\e ������l���z�K��OEI�o&��qJR�ac���'��j*�>�W3������1���遉�9�V5A�`A7|��k���L/^�J�e���}
 j��Ђ0FyM�X@"m�E��A�:Q�)�CLRa�#����̦
bO�SD�h �0Cn9`�+�8�����wz���T���i���f)�a.�'("�LI���`��\-V(��W���c���qF��'@SQ�iB�Vn��2���Z�6���+�Z�;
~ ���xf�>.�p�Pr5Yf/:,�����D�����Dx!�� �\�-��ِn%C�*_SвQLv��4a_����
=��� .,������!@���b�݇�7{�ML�s�:Q���]����x���?M�&�?�~	W��*LwF�$¿���������]�y���ߩ�UZ\U //��<�������
{��p�t���le��W`/���#e&ل�<p���MF�����>ݜ�O��`���3�,��Fhe
ћ:����M�[�p�0�m�ai�M�{�����2�*���G�꫍����1�x|���Eawt���RFxm�r<��C�ڭ��"���Ib�K5�G���ۡ��I�#����F���$_OW������v����(�K`�4H>�Xǋ)s�%��M0#�a�kG_��AޤRo��$-YD�!?';���c���R�¿C�qFq#1�^�����/f�uG�l�2�,F:C%~(/
 '� 6���V�y��
�x�<r�۷��K�f���m8p��-��ߎJ���ՇX�v�����b�թ�܁� BAQ"�`���@N�ɱ��XU1��Rv���51�9�2Ʊ��N�ws�Z���}��{�7 ��/��u��y�	V&�1��3������YEN��Ԕ�U0��h(e�k��%n9>?�q�
6+�u���\��;p���]�n���T��i�+[K�{�GJwW�~
�Q�J���[,�&�E�P�j�;��#�Lj�G8���'��CQp�z���L���ϧ#=����tb7��Pݏ�*ՠ��;u���G�6�gH	wB�F������V�޿�980OZ�\���+����'�`V�w�FV���ɦM`�iRn3����Xi5���������V�@A��\Mn�L}��D��0� ��F�4���%5�2V5GO�,��N�_�y@ Ң�P�F�^j��H�)�����+`x�kv� ֳ���}���X�ȱ�W��a��ATeK�*J`��o��fo��e���F�����s�Y
��5�L���5�������1"w;{7 �oU��?��<wN�a!(늉o^���W���;^�F.B6����ց�W?�p#�7	��x����}]Q.zH̓M~�<�h]� �䡥 )Rx'D!#��g�I��������{�� :�1_WN������>j��e�6)E!�L�1/"��$����_��.i�5.�^���P�+�z���5�3� I#�o�~����"��K�Z��l �mG���)t�i��Ho�p�����L�k�NJwD��ԅ����Þ�̔o��
|�jn���ޓ���^���ހ���e���������ߞ��}��d�
�_]oH(<�^ Ǭ:��E�Qn=L�K\)0�����3�z/��a���$k����L�|��F/�J��.�[�C(�%�tL���BD�aT���a//�*�Pβ.�>F��b!�u_�5|#�y�/���jjv������dS1�X��ѩvøN��f R�t|��A]�i�2E�0�!�5O��ױ�@]��HVK*yt���W*��O�3_��@9�v$���y� }8��`Ӗ��2`t�z�W�y��/�x�YQ�t���dUX�M��l7���P,�[� <�#��n��.[���������{q��^�'�Y9男)���G�d
ʠ��O��@�D��y��[��ꎕ���/��UہB)�E�B�,�u��&D5��;, ���[���
�^����P���6�8��)����Y᪄����;��ǧo�TE3��a�[��[^�Ir�RABxX?8~lP&7)I����<�?�U�Zb~6�)PYe�8@V���3��[�r�W<k9pTo�Ϛ�[�sމu/s5,����<���ܾV3��dM?���-1�s'���=���).�Ӏ��c�0
���M$�0���;l�<B?H�D���O7)�<$>�G�y:�{����S.�՜n,����:�L��Y̷'M�k�p�])�:���R<�oCr�VG��=�l}�ܸ䃂o�tʋ<8 &�Tء�6ЋvUP^D�]����4
�.��
5��p�Ψ��d,��n�-^�h�hN�&I��ל(2Ƒ���(�ւ�j����͏?<���M��U�B����.�\���\h
8�Q�EH�t��XͲg%������œz�Q3�+�%��VX�ŏ6�qX��~�Z0|���a���'�����{�$GK�n��fE��m�[�@f�q�>{3�A
 ��Q�i������P,%C�����(bn���Q�y^A�LX�j�r��:g� ���fZ|�r�I����Z���������#��\�cOB��&b،Ep��%h��=������U7{�kt6}!�����\��jR$����s�t�-�{�-X���=2߁��Ԉ(Ks��1�|�E���ũ9ř�e��-��+N�~A���ae�����	�_�?�Y���5p�M�E���9�M��[D�-��+�S��Y��l�	�{�-������Y�,}��(`�Z'-������Fͭ�a�7��uЭɎe�S�L'�}b�%q찡���9V%^���W.-��-J|����Fp�n*S����؇x0l������	�K�X��&�.hԚ��w�[�U�<�&��?������=��_���<첅��I	@��b���$�t5���YZ>Yoy� u���(%�t
htT�#�TTD�ҴD�[���z>��vXs�D/\������8&�G9,0fs���RIaQ�^%Q�F�~]�r�16 &�IUZ�e}3�s�&�)K� 52΂{I7�_���5�(���C�[X��O�\~&�o� s�ܺy�Q�`�Iep���S���k�����cJ�j�S"֔w2�笧�z�#K�u�g�L|�%�8�#EV����]��C�e��VZo�2���!��Ae��H!!cw��$�oB�3�b|�͖��MT�r����~>�A���lc�a��Kϛl+p݀HҀ+���0>�n�9n���;��i�����c#Ƽ�#0��;i2$rnT�nZ��_r��z��{��R}�yB���^�<��F�M�:���R��}1;�'�թ�,Q@���ٹ�M�֖j��}ך�b�qŷ|5�FM;��l��ף��6���IR7����`���j��S�����̹���S�u�������/�Σ�z������	�h;�U�T(_��rUqfR
a�5y $?z��_I���:	Ǵ�Ъr�)z���) �lK�ǉѶ:Ǐ��dU�uRp�`��	J8r5S)�E[�oBĿ����溄bMXy��u*m��X�W�D&t��]�I�׏�JX��.7E.��a����b���k}�>�v>�������b�L �*@�dCO6�3�w���v����B�x��텪O�h5�9��9,q#R��.%��m^;�a~��Жo}@{`W��5qb�ܨ�3�V˨�������'���Nf��f�~Hβ���̙{��h�N�ɂ����c�Yn�@#��ơ�v7=�w��#i���ʿ\@�.M�y��Qt�S�{(}ls�[�-@��#t��_�j}�0ք�=� ��O�2x�"����|�� ����F�x�Y���/�V�	nO��`y�GQH}y�ꌴ���9���-��q}���
��?TK�dC�B��_�/e:�j������K�
ýW�+��MO��K�D����:"�'�N���kO�U��0כ�RUE�/��ҕ��+"l=+�����ԒD��)�r��(?ك]���" ݝ����+��T6�6�J��гעY����@�/�����	^�+W����A�o"~o˥�l�Ӆ���G`�F0o
!Ӈ��;m�]�pU�wښ�|���d@q�e�,�y�X��r�m��=MeS	��Q��V��n���Q�dh��)�rN�F7���������5����޸�V !2�������!�������1=0�zF� 1���|���ȉ�k�6/�e��+�󀘡���sb��jM�ygz�Yh�贐�}(��+ω�&u�G�j�qR ��ゆ�s�+ '̑�6������ں9&�|�j���f?S nX:���y~=/��TG�-�5D�Q�t�+��n&�r���ËH��{�kA.�[�dv�d6�Ib�H��L��"x�'9s�I��7�Τ,u����q�bEb��!c����<��s�W�_U�!�ѵ6�p*ڕ�����~{_��ȈL�u�o���E{e!+ق_�clb��Ԝ����n���I�RI\�vX��	غ������ދ�ڣ_���K�K�z�0
=@rW3�o�����9ZJɫ�S�љB�T�*�ŀ����i����s���şr��)<�"ǧt��00袅����1�J\�8
�� ����q��hyB�*fi=ųh.ߎ�;Ue�NP�ON���yģ�`E@\�DM��V��%����)!��ၒ��c���zR�_�U� 6ɼ�����С(cr�tԍ�����޸�!�=��o�[?�e�i�b��l�"-� bO�ϳ �@P1+��>j^K#�������Q;���r+�	)?��#�$�C���8Xv���l��d�٬�H��<t-ի�4 bݟ���w`�<B��c�|�	m��K�d��_I�\�\H��r@���c~�ȉ��� 2Ȭ�Ŵ�b�����ch�5<�E����pZZr��9�/�Z��f���i�U�U��T!���:gv�C��/�����M�i��N��R\�g�/�u�W�':? �Q �ک�R̈�KL̛%V�VʜxN�j92X7�U؎ҸBP�ܙ(s���O ��N�G.��$e`O�@���I�Ȍ 5�&��>ԮJ xʈ.�����'P�O���-jY�ߔ� ���/v4̀ۇ���'Əڸ��l�<u��,�`DLqQ"vms^��Z���\q�v�%![t�Ĵc�ò���J���]���C��w��$�;pFcqgD8 𖩗� n�,Ӂ�{�L)bRc�����ܨ�ۨ���RB��1�2�f;D���獜�4�r1�2��<e@�{T�>%m�ք����S�<P�D��>�Y�!W�W'pp��5�`B����=pI��ݭ?��4�A��������=��R~���� ��k/Cfh��G�+��t��ʾg>��h�wx,n�1���Oe�A!��%<�)=A;ͤ6�}x��b����1?2?*q��l���ԟ��������Q3��za9xQ ��N�"Ԣr�����ѱ����������ɑ�k�r�I@^���?��J�G�ȴ�?,`��o�B����U�Rv�����e�}�����'��+{|K��z�k?��S�M�V�� t�񇤆L�-�;ҕ�A��L%R�u�y�3A�@L�η� �~ �.ýcV�;^��`��7ҡg&!f,��9�:q[/K���S����hl9_����~g8��(��!��V[��&��>��۞���l���Ĉ�(C�"ve��=r$��L�,(~o�4���˼��]���Ä�#�E	B���u��S�DHM�!��(V8ʇ�n��ǟ�A�ă�!e�
�b�9@76N�#g�	��,�'�2!�CG�/�i������;8�P��c
D�0�S�{$���=��XX���n3���BɆM[k�Ɖr"��ÊZ�?S����@�(���A�m��Sz$w_ʟ̐�<���q��y�蠠�a袍W���hu������F��g���kG/;���h��ֺ�5�#n6��V�N�Ē�S�g	�0;�n�'�Ȏ�@i��e1w��{�/H��pגS�F�R�.���"�6��
[%��Z]d���BO��k������RT�F*i8���vRC����*}8���Z�'����cb�V���b�x0d�i2�+�py-�籍�#>��g��?p�p�����FjA�6D�s�dΣ$Xj�ݽvCj��}��ړ��ܿ���z���l
��zf74�Dch}(�UQϰ�U��\n�+��5�G�>D{-;<{����d�}.��
)}�����1��41bx 0�lr���-�u~#��N����l�-{#NGg���������PQ���y��)ѭ���~Ǳ�q^�ǢY{KC��6U2݅��W����7����{�Wi<�@Ţ���_�5���"��!�ÇU"wg�E*ts�s����"��w����L<~����6U&	��hD��Q�j	3C\����-W��̮dV��Ly�MμX�Ǎ:Y��w�Q�W^L��}�7��"`fuG���fGv�Q��P�}X�:��$��Ւ�?�^P��?�b��S��Q�B�A�9ᔜ�1��l��⣛�D�nO�/�����k|����D3��mlp~s��x����p����H�m n�e �0�dw����Դm���6Ky�G�ʚ�1�+ �+��5q���_ �y�~@v���&�K>�-1�����vm�b���R>3~c�a�mW�R��gM�h�t:�'�<~S�����e��qW'�zO%���< �N�e�Մ�]H�|�B1�c�Gr��ǽ~�ov���n>�[���KD,'C�Q�������jM�����I���f@��G�%�|���$�����h,^�&XH��G��B�e�hԲÖM_n�|)[�ʯ��!�.�YmK�Rq�3�s�ϧ��cj��#����s�c�<f���}�f;�@j�wfƖpG� E�M�l��;N�]���J�2G�ǹ��#x��5�=�5���c�oNT{y�^̮:�5�-�����o�ܮN	���	�w�Q�Cl��Ö́YH�&G�v���-:]����AQuX٩A6���-��!�_3��M+<������O�����:����J���je�������_���P�C^��A�t޲(��b��nH�7w�@E>�᠂��>-�h��d?|A����gQ�K�fqs��ץ^=Ô�a�k�L�'0�9�Y���u@��u����/��Ì{O��ӚJ9O~��Q�=�>�!�\Os��m�$�����8/�Ml�tx0vo���;��@�2��$��a�jb���,�}���0k*����L�8�(�����W�k>@�K]&����i��\RQ�+ sZx�iI�d+�V!�d�i��8�]1B2p�{�M#����X9g���Εm��a�Q�l��~e�{��<'i�`�tG+��Gہ;�A�N����դ����w�Aw�<�q�G��9ī?EPC�5�v���'��[ʇ�]_P��W����[���V�??k}���Uē�����<ˣQ�"!2Q!G��f�.��KQ�	�r{�M�df�a
�Ǿ��?�\�i�2e�WI��L�⑀QZ�B�;���o=��+vg��f�)I��V���o���/;�|�	\��t��G��;�Ň������x��)��0ޑc[&bnq�o	� T/<�ߐ�i��2+���&J�iw���[��������'JNđ��Y�H��]�4�3>����خ	>9a4��ɐ�A6čq���&�`l�:��c����3������A�t#I����}Hq7L�p[�j ��������|��6M+�r�w�G��9�}Pn^Ж��w��k���F� ���ҽ!Q�����પ)���HN���4�������n�p�F�b/�0�<$?��=D�y���ej�h�7�$�<9R��$�LWp/� GO�M�+>}S]ɩd'�O>��r�l^�s�@ٝN�}b�i����4�7�O����z����6���
����T�ʑ�u��iD
:��J�W��~J��h��Ԣ2����'閤��� �l����|��,Z��i̇�Y�6ә�Ah�Q����4;HL����X.��ת)����'����墧�]J�F����"����@1��?�/���X�Ozk��E���*&�Dz1�3޼��v�U}:B����i��������~�(q�WF;nm�ג����Bs�u��?&-��[a���	JIF�+k�,fc�d:�ţZHi`�M�<���؋[�p�9�E ,u�ݲ �5����Q۸��[c�z�@��j�7�ށPVؓH^�{����9�?x��'��8X�D�/�n����Vq�~V�mb_i�sW\	 �~����;��kA` �&T��]�8h���e�\.��DNVx�7�i�hO�Q�[`���c�d-��]�-v<u��Z�v�޼�#�~~
�Y0�	����.�kx���~R���l�Ьh�{��+l���:��'Cd��ԍ��G[�<`7
�� � `%�Gz<�/�K��]��qL���0�֧�CA"U��*�I�c�8�r� �',�[������s1�������xo��~�@��!����ȓ���n7���X{YG���w�[!���W�R�	�@N��=1�!�d���+��`�ɩ��4��!y���h_���)�9���bב-F.��	�A��T 0U�)o/g3�f�\�$��&/$5+�O�+Ǒ�b�n�IR�G|jf<qwp0����'�����H���QN�ם8pz
��%����)��ID�D�<#�	�Y� �5�Y��IH��M׃k؇�2�y"���K?�X����������K�6�LS쾱Ӄ�MԘ��rw�B:�kb�4�)���H 5e�=�Rd���E��z��h�͏)�@����$�1�<��r>�N��r M ������� 6q��^��Ȋ��HTs��	$4Z,�0��e	����Z��3�7]����1�>�~�m��h/��� � RX-D�b3�Ƞ�������N� �H`������Z�Gڹ�Q$H� 94$%f }O5����P�FQ�R/d��1�cGߣ�~8���z��w�#�+	�/*�,0*"B�{��������P�qz��^q��}I}R.l�I��8Hn��`����%��㒕I��lڏ���Sa�����Z.+yK>��#"~P��x��"��ǂD�"�?�c5��J:^�1L��*9��K��4	1E rÂ���.���-XF)ǽ���I����A�k���Zw�<
6k��3����9��n?�k��~*��XBp�������	b!2���F�:�-�C��P�(��.>n^<���ƴ����2�P�׺&�Ђ'h#�tMb�BJ�/ԃ�H� H욦���_��3�<:�cT=��-V��,X�
�6�Zv��`�W��p���	��I�����A�W���X-� ]& �c�lC�k�7��٘ӫ����/�/�iB�ګD��y�@��ǿ����N�|���ֲ�"e�G��8�YS�	A��S�H�j��dN@c�>�=����:�)��qB�o��	��\�۴SZFJ���aJ��{��������ʗ\�X
�%U? ^���r�	��}^�c��gR���]��X"�H��
�8׎E�8#������=�r+-��,mـX������]��#�����G8���n���3��EB�k�s�ΦہI��޸�K�* IA��:�ȤI��_b'0|�F�<�u �R�C�a����?�5�2󷰛#�TOBaȍ?���V�3�H9��R�R�t�Jz���*��=a�#OE��d^���q�Ο	b���� �Z��5,�Zl=�M�����Vxŏ.��`�9��������
��0�qQ�.�|	ő9ӧrD�J$��:�� ����L��ܖ�A�jf�C�@Ֆ�U]%����!�2���ŵ�7�� ȼ�CS�_)V���I������LΤ��[���dy�hb@e
�j��f��u  �Sȟ�h�W�|��w�ҥ�O[���<�w�)����&���)Ρ�5~���L`;��e��U�;l�t?�!Y4��a�6��P�����J����^r{ymÅ�F���Pnr����;�Hj��K���D���T�E��y��ǯ��_z�Ixѭpd���  �:���u��̦:+Î٥��M����k���S!g�Yf�N8�L��ՈI5c���� ��#9��i�����(�u#��
�H轙�=�M�K�7�l&T!k����ɯ�w$�Ã(����C׶���T��e��ch��z뎴^@���k@k�*O��e���>z5��@]����b�d*^��ȴ	�e����\��ɋ�o�^�ќ��=�^�P>xNd��I��D�`51���7�w�I�tƮ�V�r�W
���*�ح!��/�!=F�+M�Z�^�yGH2���+�/ј�{8$d&��d��ٟ�olsi6�?v�)\f,L�����Qao/�eˎYh�~��ŹjW?�-OE)��br�uC�9�j��RE�y�ͣ��eM���ݴ�qC����	��֣W��N�0��Mds,�-�J�J׆,�c:��l٩o\l�&��`{
]uN+_e����f05R�t����� :��7-�rc������J^��#,���(�X���a��<i�,K����6E{܎�y�]Q��q���]c�I�"�ܭ�7�G>ӻ	@~���q���x]K�Wd��h+�?��d�u�[Mul
�K���+ ���v��`[	�48Y� �gZS��ɭ��4�E����_-�ְҜ�˽0�@lUr���^"�5�Y�Aj=;;�9�C���?x�џ�%��z�ySY<��B��1�y�(C��1WԚN��C�� �
z��|��%ȷCʏ N�����(��)m%�<���_��Sխ�p��?���!�:��'Ž�5��4yl0��[N̴���{S��Z��4e X�� ���GZ ��;~n�(�7ʊ�*��ʾ�����:� �j3�j���-ET3������	MǁnSJ��{����F�����'���f�v�<F�;0��Xm��u}��3�r�-�;z6)�5��c�k�8���`DG�]����o��&9d�,�a���.�*�?%�r���k&-8�%�7����gr��5d>��%�[t)�C�i��K�b(���t���.���)�,�WY�{B$��H.�ȡ�^�j#��I��P��%9�ʤ(ҀZ�&���XWe˔ �#�%�K}���/�)��&4��M���9�OׯL)�H�`s��A�����x��	�t����Nد�1~�+���l��[~C*-��{%�>K��}��]V��Ȗ;���^S[��r�ǔ)��f�2n���}���l�(���l�e1)���H�^�'F���r�N�S>��wL�����Cs�a!	8u�'J��Di��Ϧ8���7�EJ�����v�������*�AF�>�lk��B�Ҡ��u���N7�o���m��[Ei�����d�ZQ����:�k����#9�o���(y��:����ap�ɯ���Ӝ�Ie��k�z���$���de�y��M�E��}������߻5��X%��~NE��Av���t���b{.�Vm�Dd����+f`tŨ#ez0�\�����U�xQ
b��.��yp'�����wh�߬��!��� � @��֭���D&w���?�'��V���Ͷ��Gk7���_m�5�V7� ��[�!��ǡ���|�C��Y�^�'�-��Ǚ8u5ri޹�vE����zhQxf~�q2���6�]So������䷓pɏ�ԄOZc5$��5�0h�
�Tx1� �L��!}	:$��c�tI��ǩY�<�]�����Ɛ���9��%49�A!�����E�J'�g=��0[�K���㜿�
�D�,��b�{!�r{�lk��(��_�P�E;���*Zu�2�ا*�t�Ԙ^Ƽ�A��d�ZL�[��h5��_��v��1�3���S��B���B$���x����(`S�a�� �.���|�,�
�<�C�j% �U�3!���afj̐T;�x�]I���)�~L�����G�K��Z]M �$�q��?�e=��� [�&�1?t�8�Dv�ɠ�(k�;�"��)v*Q�Dnc�QfA}�M^F�I�=�EC���Bc�������"[!5R!��7�#��n���=(W���mC�M�>D4��[*��} �ȩ� � F��W�5!�i�/��hl���
����[d�ϼQ�岕m����v�pB�Y�拽���@�{`M꘶�B�< 2�Q?��� ]��?C�w)����2:��H��I?�#J��$DT	/�����T����Ee���jT7<�\�� r5�^������.Mu{;�t��Ub7��`a]ՃY_pZ�����ɜl�Z_[jӥ��W�����֕����1�}q��>ө�fF4��j��32�t��y��D0Y9��N�N�!M:���`=���&и˩fe����f��cS,���Aۙ9Y�.T ��$�ָS#��h�;��KaA���P���򛘡�5ꀿ��L(��F�@�d���a�"�ўd{$]8䧑w)�+�2>��姨���[9<)�����Y���Ł�\���no�hb��5����㬾H�4m���3����w�����+�@7�u(6&�� �G�Z��y�<�/>� ���m٬����BK@�r*�ݟ�8��Vz�8ɾڴ ȯ��P*���i��)��J�s���� ��$G�A�ܕ��E9�d��{W��U{���Z�Il�j�h�����8b��
�|T�(�:�63���f��2�zܭi��.d?�#���J�H�̍Y�J��M�����e�d��4̵�M&�⪢�\ů���mđl�o(�:����b�>���Hj'rJ
t1��ݲ�����N�C'B�;��Gp��ګ���"#�����7�iݲ�A�؍��/S��Z��]�U��Ȝ�=��n�>���q{#��hM@�`T�Fz(>/O_�p}<���_)�����]��q�o&O�b�0P0Ȇ�^
��:n��+>s��D�?�x�־_`i:h���=�[�6��9�P~��Emv�ЛJ�&�r
��-*fD*��T� ��L�g��[���a>z�CMOK8ځ{A����k�Ė8֏�+��AnR��s�aSM�*P�9۵ޯ��E�h҄'Z�o�?J^��=�eP,�W�#��Fl�&�X�dj�؛�w�bO�"��{���_ ���b,@`�:�ĄCt{$��َ���{9�*�	�0|]h��\����#7�$�l������������{�~,����PW��[7d�����%�Pm%�.��=��v.7�fv�+is�e୻Z�
l�qS�����@m>%���K�>97K�3��y��:��Ɇ�rE�Ҵ�	:[�/��ؼ��~����P�VO�za�(iOن��̕��X_�X��G�v���3sKd��F�_�L�"4��zXѐ�Ǯ�oj�y���1�u ����t�����5�b�E��txY� h��.Dv�~}e��1�2�]��,C ��������Ws $��� ����V��WG���|�W�%��~�l�Ͽ�ÿ���  YbxkM����1�İ��~�N�i��|�si��|��?gm@P��70��V��!��� UQ��4���2�HD���g�bVrްI70��N&�b�n1�\�bv)�����#'U01���!a�.��f�x�fI����#�| 7� �?���j=��_ۆ��0�����=
�y,f���mɦ�r�P
�9�e<w���urJ�T[���v�� }���D_HîjK\�1�5͝���㤮᰿\��Q�����t���{"\&7"��A2�?N�1�j��ptOBF_���ңR-����DQ�G%/W��=�G���z����$1�N`��zX��k~��e>~�XK�y1f�6���-ڜ<b�� ^ZU�	�`|�iOXq>ic@��P�T���P�(2.L7ՠEAh�ar������I�[�*x����b=yrQ*D�A���>?wy���ij(���l���yOӜ�SseO�+r� lح���Rd�S�~���-V{Y�O��U��b��1�Y�k�6H�i��_�܎��٦���>�ʺ~!Lw0F�G�W��+����0��ҏ��N��ޑ�\�X�;[grY��v��P�"Έ�l��"�J��fe��"=3��8����(u�b���S�Aj���gL�}��o��޿��.�2��΂�5q5��g�t���x��r���ZA��Q�H<Z�Eq	�C-}��R�Όh��g���;O�Ͼ�����h����Eo�w�r�'M�j�u9y�˧ �n�c�n��3,Z4?r���3vXkfcϙh9pW�ΛgJ����Y��7ɪ��Vi��n�ji@s{
�6�*?�M�M���e��t�:ɶ8b�j�lA1>!B�J��1&��^.o-�����WPZ�D^��DP�6O�qA�F�2Vk�>��+������� JX攳��w��KH궜̶BA��w�)�n����Bj��~!�]R�� I2raE?�ى��)������?s�	��ٷH��|m[�t
�}��ʈ�q���?��if��u��Ĭش��iD���L�&��N�9���o����H���u�z���w���V� 	�Ӏ�dR�$b�7��$;~6Nj���C��U��g��t酴�?�:!T"l�0S�̿�Օeo
C!t�R�b߶�f���pg��w���������B9��d��〡�F�ŷN� ��)v�L/y����'��b>t{��NX���u��Kѕ�����Ξ��ᴡ���=T���^8�`]��9���|_���~���((�t:j��pÞ�aE��?3�O/ԡ��ŀ�^�'�"&��`x�c����w��o�6_�3"��F&�'8O�;ҋ�Vp�8/�ᘢAX*���_�g̽_j���_�^0������aߘ&���x�i������A&6��T���YnĽ�C�&��A��e��x
�*X�d��nq|(�ӟB��x�eZ[HtV3�u�\6r�7�C{������t�Y�clu�U����4Ң���'�憅����TYb�b=�w�m�~�	'����Օ�^U��OȒ�'����.��-s^���Ȑ8�ߏ~Ո��S�����Qw+�.�Q͐�R.��(�h#�(CY�ϳ>A�AA<�
�e9��C͓�����E̪B���S
��e�H�b�A�O�M��d����Y�Vp$H������h61��Dk)���Dn�r�̐:ξ|�`!����(c1�.��P��@�Y���ކ��Y!��d;��K_���ֳ)�B��2P�_���ʼx
�-~��	>w�k�r���e�h*��+������3�4:q�A�nDL�`Sv����
\�;<�I��vKe�6E���X������|*�~1Deԅ�(c�k���I�!�%Hz�C��ĎN�������i�W�e�U����?���B�`K�<z���9�����j���E�������+x3����S���>�����b\�)�@���4��N^����5�����9����S��w��xY�\�
r�
�2�`�$r<�Lm�2yf�[=�N���2��9=��M�U
UV`I���xnH�?{�v>�1�Ygzg�S�K���X\t�,�k� ��՗�@<Z��:�ML���]�C���>�[1Fߊ�0O�nՄ�*���k��μy�w�wA=�s�x�v�i2�%�ݹ a�QEǖq�L�!�L�����k�w��Yi�Gc�8�k0��!���{����Ȍ���$���㓿� [k{6=���K���JU詓~V�C��&��ŋ��>�D*�Bc�w��К������fXh��?�9��>E���:�7=Q՞�8P��<�PW�#Eg�t��&���:��A�iq��skPp�:�
6��Q��	xei���S7��EV?���rݻ�L�'h�A���w�ǯVx������s�������D�LX`6�E�����ڪCY�'�b����\Yz:�*7GF���P��>f���}u��i��P}���|N��ȟ�h�϶fj�d���j�O��Va���w�֖X�Gf�z�癆ñ��#侒�?H[��)	�P���a����Dd�|�W���H+��@�Ɉ#;A�4�@8���b�	��OW)������*�A	4��jh;��q��8.��GGSi2��A���]1�f�yɯS���'��Z�
�x�cJ�5��0���Bh&�w`�hm��z���7��Řߩo�a�|�*5�fj:�2&w�h[�s���$8�m�92;"Ɣ>D��Xn��]�!���G�蘚���&��+P�Hc>��=}�(�i�SMq������K�w�����t0�H|�T�3R�bL@)�����*���RRq�@�ٖ�T�N�ARNf�����xcL��l�������@��(F�b B˙l�JD0�4o-,��C�R�!n�
�uv�%9�0�bx|J�������P�X�\��ʤ��>)`���:D��P��p,��LF��{5<�x?ʥ�m�t�:��-�a�����լ �3��T��H5C6-G�6�UK�����t-���_(�
h{g�R�y������eG�_4AK�������F������BTO�I�M&��n�ec{�6���]݃SS��\�(����q��N�&��V�F<�s�62ߑ���!�\̶|��O���/A\0G�+�b�u;z��Uqѕ�\����ˀ{�
~5帉��]hE��P =�d�88�>{��3�F�0�Ϸ,t�+��V�< ����l`�	�3ˎ=:��Nq��d�:Z�g��0���3���Rh��~Q�)P�u�J���ə�+"�����3�O.dd^�����
�j��%�1(�V-�jI�,�aDl�F���� lK犋'��'Ǜ�*�|��Q�ӡM��PGT����8�9߯�����No@\�4�.'T*�1�D��61O�5��@�C������MJN����n&� f�m��Hf��ᡱ��A'��r~'�j���X|z4�t�x)�y�F�|�U���~Ġ���Z�E@ �#��w�e���m�st�dD��6V�|�Ô�-�����A�����H��߁Ԕ������cϬ�A�����>�
������gmoUf���r!��
�A��NR
"l&�+=��>����]�J^���2��g�v\9�grX*��ή~A�<����i��RLp����M��,h��������{%��v���!�j$�}��9�JR�p[Ht/
�arR�KT�-3AB< �E�^=��jN(f)$#��쨠"��c��^�aW�#c�aC'�e ���Z߫�Ӎ&u�]�'�&�h���9����W��lM��V�ȱʗ�0�[�M�Ca���P�������;
�6zt�1�q�s�稿��� �r����"	y}�V�B��y�/�I8P����,U�J��?����\�O\uB���)]t�>o�i"�IUu�D1a��"	0[╅�3�-��=���d�p��N�;�=�a�C�7�D�740 ��8��J3\'��ֲz�Z���iL�n�
4i��{���ف
;M֜`�9�R���~�q�ͩB��X�	T@��9� �wlëG����k�4�՗ʡ��][t�B��	���5�P_�;����ϲc��%z�￧mZ�J�?�#E�oc57q=����7)���j� ��Lp煠�����5	V�a,��+QmU	�������ĳN�+���L��.#D�!Q���R�[��6m�t�@ϣN�ݡ��l� ���
C�9.��0�~�MN�x3��Ƞ�Z�0���BR�m�jg�ٗ�8���:�r�eJ��l��ZG]����Gx��+5i��	D;X�E6A����k`wS{���ϟ6������;C�ݯ����H�DOk-��,cR�σ!��������oUp(����?�^�ժ�����/�5qEЌ{�g����(�R�����v��=Z�`Î"(����#A{��**�ҟ4M*��[1Ol϶��f��x�@X>Vv��K�>'�\Q	�S��P T0bj�ܠ>V��Ş�$�e2��6;'�vkx�L.`�ry�Zv�����Ix5ke�7�Ep�~g���� �ᯄ�Xi���W��`J�BI�"�����2 DN�y*��G�z�̑r�N��&%{%B�ǈ����n��V��ae���<���0��$����fQ$I�[Y����x��m��|{k��?�a�s��G�|�Nh��餂Jp�������3���R}>JA�',`{^��B#��h՝��^��B�O�I ���� \���A���:)|m:ӯ��~�"��.�?��/�j�x���Rmu�O�0r�J0��q�܉a����}�[�-�{���-:�0�W�w���r�Z}y�9�gf�Ho>��w_�x�#�RF��a���s��J�ŷC�o��u#�SOe��l���Dh��ܦQ��$�� ���4垦�7ol�����wK�FH���( F�f{��S��k'|fpF�G2�H���?bB
v�I��~U�1(m�W���:���X�[v�m�G��禐��9?�K.��Cפ�_��$�Ƴ�Jb������4Q��v�$��x���RVs4=��{�Ks̟eA��`�������맣�;���J�&h|X�\8�ߵ0���3*%�g�}i:�ݺcr7J��&d;�7�D��V1��Lj/G�2}�{1q+�j� %�;\�5�~e`�$^�op@[��{�OP�*����
��H��M�;�@��S���aH�����:W��<���b&�̑�J�^k���
QM� NB�bw(���RL�2�$f�ь��Cz��3a��E�^��a.�|Q�z��z�O/n'�Kl;(�d����'�.�?2�ׂ�L'��@;��a��p��I����Zd�Q-�=J~3�F�q>D���5��Xx�Z����q�9�B�rc�l�m�����a*�s�8Y	�������n�-!ڢ�b�bb/���^���=��d`�8f���/�	�4j���>�٠����CbZ�`2y6i��q�������쨃А;�Hs¹�!���Z<3cH0�3�1�Aν$<>S��ҋ�v��+�I��H���ꜱB� %C6��c�[x��Ӗ�*W'���K�a8h0�D�sY�*%����y����%�L~oU�ˏ]:�ic(tɩ�o�Lx#?���XQ���>՗O2x��*�3U�AW���8wB�W5��7۾73�5�6�k.f`�Q�i�dR�����%��T�6��
f�j�0����%E.��)h9�1Z��taEt�Q8_?�ڸ+�|N��`������MD���m[�%�F<#���$_o����3`4p>�vs��{!Bׁ1�&��9WK�hbf��N㫐;�rh��S�y��Eߋz	��ݭ�p�����b��a�8�ǋ�1~�R.�+P�T�P
^R&�[n8₼H�����|d�l��I��tB�D��[<U�����=�T��n�^o�8o�eR���S�{�I�y��lp�=K�e� Ls�����SW��!��[���)7.=�8����&�?~:Q4���(�:3���O��"UE|.��7��2D��Jg�L�%um��et7M��~f�=�A��7<�i ��q�s�Pbj�8������}V�M�C��P{��l�J͟�e�d5�TL�%!O��6�k���[~�E�X�-pU���������i�'I��tMԥuUp�˒t����F�@T�L�n�)��H�����Q���j���Ձ����\^D�z�j*E]��r 6T��͑{�{0��v�� �Q�Lo������:�f��>�9�8{�$�PǠ�<:��z<Һ�yA|KTݪ���r�ˌ�ـ(���8���C+�zc�E�
�#>$>�ȴ�N>�$V66�l����n�&*E�!���
�e%�Y���2��z��G,�:Y${��묇;��o} ^<�_�*��xG%����ҕ�j�d8 ��(9�)�M[���j�\YBA�b>�����Z�P��Ś����Z�C/�VV+ו;a�(W����ξq��錆t�m�6��OR����y�TD��?VO8�2��
��2xnV��1E���#e�H+���`�b���k�v=�����7�W=��Œ����̼�_c-�`��!��� ����E���0���hl*�r\h�K�.��h���a�Af����4PV�w�7Z������%p�����"�'9���ӻ�q�+27R`R�e��G1]q݌m@R�����g�ń+|�������*�x8��2�]'3��X���T��w�'��"g�DU���~�]p2�3�ekә0 ����r{F25�4����x�(�����5����V"������'���2s�|�b�1�} �ˢ$S���d�H�>�e�� �R�	u&���Ui`�>���v���rG��	2�?[���F��3��$�X/��#X@�; v�� ��D�C��B�h��	���y?�M	�~&��*\������r2� nW te�Wz��7(y8�����G7�<�oĮ;�L��:�_�o����=��nN6N���Lg�g��qÐc�Ǎv/�ߵ��K��5P"���p�����C�P͛���	�y�0~4Gr-�D��b�<����9=tB+B0�=A����)K��'�A�N�Frw����hc2������Ng՘:=��Qn�:�m�Ҫh��qU4X����ʞY�<��7��b	�I^W��� ~($�s}
)*6�u5|%�`^=� ���Q���iQ�۬�e��k3dR��̀�e�P	E@e��ac�N��P�d����$���P�G\�>o���P�x��=���Pg�$�`�W���Tc���Ud���A9�B~ʽ�~Đ��w;{�,��(,�>T:�hJS�޾��h6D��e��?�uC�iS�w�W�����Z�}v���4��%�VQ:�ӿ�/_�h����'���^�t��z�%M�@��v�ʢ�;Mg���~��9cC�M�j'�Q[���RҺ����d�t��`�gC���rkH���z��Rɮy�N�1�����MU����^���<�8��̖fYZ#[���|m ҄��Ԯ�`E����As��W6z���I��.1w
e��&��n����},99eK]��Iw���:E d$]�yuke�:8���0ka�߇toR���A��ن��U:BT���=�V��z�j��/W�J��������mE��n���SUp�j��Q޿�[^���4H֒��4u�vWy�4Qu)���Ɋ�?�|�_uM�T/6�{�x$���ѡu���t��8
�#dhL�[;�uv,a�rB���)dW�;L��悹�I���E�+K���|��j1�k��	�s���E�����zE8�&�i���'EIM��D!x*"x?�2�p�'�5>��~��Gz|7ؾ�gӁSPmC�SAX�ns��aP���w�<� �#Wo�"���VF���C���fl�E��s�?D^�$ZzbBC �e�ȦE�n�}��f������c< A*�x_���	߳ a߇0K_"�%���
D�0j� O�9��P��������a9�ZA�h���e�j5��|�$Ml�4����'�Q(�憎dw&��w���K���4_� ��49�g�j��bܴ�a���N�&��)+Нr�Y�~�8�k���i�H�v�ʔ9R���ø��ٺ��q���&��k���3�	�7�T}M���3R��9��2R8���~˞N��RS�Jy�*O��p
-�����[�J(W06�B��-����fo�Y����~�� �����qG���h<�sx湜�!�
%l��(���X�f�'�[	� ���В��)D�k�R��]���6-|�~cXx�@g&ݏ �	��)��[Ǩ��q�$��2�q��	�$~Y����WuK�os���H���\��f2�T~�ٺ�޵��9&�;h�ˑ�5φ.Hl{��/X%u����c�H�rx>y���cL���a9�W��`g(���s�o>]W��Qb���1h�uc
�׶	)�Pv��o9�P��Ѫ��|u���9�0��'�z��ΈA���8��!�d`�66�]0��T��H�<+e����m����Dg�`�Y-�ؤ�nHB�}���;�l�X�E47�MA�-���*YoF��dζ7k΀M81e�x��H�#/'oG�p��TtD=�V��V%L�����AP�5|N�Wn_. �*��������cF��r�p�o �������=ڵ�"wV3�y.oA�����	Z`Ԟ�6�Y�v���k���^�֫O�Q˄�)��{�j�^N�@�/��>��i�y[��rC��f�p�xݱ����H�0^�j½�� /*?L�;#�,��8ʈr�Ƙ���b���"h#��z|ڢ�3��;���5��P?�c>�bd�E�&&{�a��W�ia˄��!�q����<�򂢉��Z�B����ԑ��3W	����?�y\�FӂE��
�ػ5w�؎��DV��*��
���Ụk�OO�3���f�zik[�j�m6�I��x��f{U��Q��(ލH�3f��֤��t�ŢT�'�-H�;�j���~�`��i��~�h����[�rTȿ���9�itCLnբ+��X����[��_���eSq�'�u�(���j[�-
+��e,+>d�q!_?ķ��:�EC4<q#_��{.��ρ�Zq��;� �kxa�;���D�,\.̚뾋T�ó6��JG}�;�|��CP��b�;S��+ɟD9�ya��H��������`�N:7lQ)3v_N��r@a<���̛fyv[�E�3�<���b��b�6+�}!w^��U��ūA��2�7x/��Ie*T�a�vv$�V�%�� x~�Vrnh���~�J�=�fR�(èď�E�$v��s�.��v���Y����AJ�[15G=q�o��;��V$h������N�LG�d}��s
�ᦘ�ūY2�����D���2�+�'m����C@F�.��L�<2��p��~�ވ�}�PzN�I�VÇ�xN�B�.�T�v0:SG��������/d��%K�:�O�g4D�kK9
}��!�z�d���5u�����@�u�0ԚC_>0�+�@ȓ-����w��42y�
���F�u�CHX��%@˪�-#�h�Q��΅l�L�V?Oz#�1�4�� �Sב�B����a��鬾���]�{,�c#҆67���Åzn��!�`��.�;"j9�AP�-/S'`���l�>U9[�gpJ�1Q�5�_@�����6�%�޷�]��u��i8'鰝���b^�9ƩЛ�� �'����RU�Z��M�R=���t��;{\�`��f�|8%�6cQ��i>�����&�b	�b)W]�e���{f_��ѯ�HqK�ܑ���M��Rrϣ�s�:?�_辰{醑��B�a�~U �p� �ǋO%r��<���i��"b�Ylr�l��v�jV��('	�> ���N�xL�����LS������ �����H�j�l�>A����JF�(�b���ЊSOJ;���K����.���Z�ikm��-���k� �dʌ'_JM�y]��|H�C��Q��j��vBSV��)b����x�ftڳ͠�jz	�64B�	����7���K#Z\c;�m�]�{�m��0��������@��E��Vi��hh�=o����*�yI��	�Jt�~c�a��R{o��_�P�����i�[�*��O���u�����>����F�*o"���q���9AҒ�T���_rL_m��U`�i�#��#��s���*�)�5�ҟ�@$I���n��ţ�`�U'hb�J��_x������Wf�Pvl}Ͻ�\�䎦l�S?#��A����1��)`PUogXk����V��$ˍ A ɵ� T5+�R�y� ��ݚ�r9G���&�Ή�mj�u��ٛ�����ri�1Z�]V�2��e � Na}�3ܣQ���t�x��fъ:�;2��v��ۓ��aV��~h�Z>�W�u��t�͆�چ�ĭ3oO����T������r�[��� ~S8����ֈ-]�~M�2P�i�Ӥ�~JP��
;j��ˆA�����-H����T��'���@#oa�q���� K˜3Z:e8�J6��5$(��׶l�?4rh�������7oa�@�l{zXo�a�R��Q	�d2ͯ!Tְ�Bp%u8��?9�-���}��M��e�9Opj��A����D�Fu;R���S�����K�;)},�vE&0��B�m��a����L)ls�t'��C��9 �g5�u�z`���,���h$!����z���R(��˫ԣ��~�<p��!�:��@��앀AC��&֚�(;?�#�2β>KZ�`g��n��_�HqP5h�s���V�b���)�2&bb�}%ӡ;�ﺒ��Ma^z�ۑ(��D�G��n�X�����
�}-~�q\��F��,��E��(����>鸊z�{ε�����^�Yᘌ7��/�����T`ϊEqy�2����Q[��o�AV�>ʥB�"�_n�ɲ%r2��/T��0�b�4�7\y�����f<�1���Z����z��/6k��y�k�|m��B���n�����7��5�%��7��^���;e$�zv�\�ۗa�[ƴ�#��8�4T��n�PT��)�	�K3��W)>�����[E������� c��/��f��	�����-r�[���;���zIV�>Y�_ȹ~h����� cp�+�'-sn� yx�� �+�)a,,��W/�N�[���`ޗ��_��ւ�����`��V�oa6�">��bY��6{��s�R}����/^�7y|�<�o�8S�3��Z5�81�g�u~�a��C�~�\��
���"��LrGnf�D�:�����P!YS��Oq�	�Z��q^j�wj�ET�7���(?_����w�������C�Nn
+I���hOX#��f����a���U�-�>^v8Ȧ���Y�!%E/�0�����
q����c��Mɝ<����X��)LF���Ak�M�t���E+`I%9討i���!�M��3T�:)��=Z�O���?���BS{q��t�quWqo+�h�����hC��cJ��2���U��1�t�n)�{]���߮�:iO�r�4	v��j_$�4�A�)(~V�D��˴�I�f�U����*�Y�'�Yе��7��) �p��P��������V���3�-:����
���k��t��B�B��<�K��t1nA�ԜA_��s�:/������z5�-��<��U�d�̸����B�L�K|:�<i����^ ��Z�_�\���u�IſAMT���Y��T�~y==%���ݦ-`��w�L��}����\���V"~��V��%�XdMŌW*]L�K59�#���kD�a�ٜ���g����8�ӭ�*ʂރ�I�=K5¬�nX��rQ�1�fܝt����2��8�������eyv�m��}g�{�O1�^."1J�4� ߡ5ȞD�����W$�v��������N���1�8B_�Ax�����o�2�D@+|r�y%�8�L)ꍛ�]͓�ϙ�!_����.��4 8���ҝe��@��� 'p7����#v��p��=���gu_�>'�ZT7^yO��Xh��,�z=0��:��0Z��@X��ˎA�|��*��;a	����yۉS�B�Ͷ��M����#R���?�2@I��B�X�2�HC_���
���z�t�.�l�� �|hI�I�c$��&��r[ÝU�%7�Ҝ�Lܠ���{$կ
(��%����qY��8s���7�@�����j�K밋�H��f@�ަ�(L������>���,6���pcE(A^Dd�^��(!O��]�Jj��1���RVL��9�D��+���P/D��Ǹj&�T ��O
���!��ܜ����8֥#�\%5ث�)��r���('Ӡ�%���?�o͔a;1��B�k�#�@f5I�@(�����/ z0	��I�d���;�aĚO�~�wg�vL�Z��3��{�do��ιK��$�ñ���>ՑȾn�z��St�[�����G�CjT1�,K*ն{��L�AY� Q����q^jS����q��ʡ�X��(�}M��Сv��vʹ�,��5Shq"�T��'q�_�$��XW���a{��� ��^�֧<�̻��*:��.�lĺvª�7ŭC����.�����(r�N����܋�"DA�%J�R�2FM�Ģ�}H�LY�s����!�C:]	H��[��%�.�,]V,j ��r �q#!������i6)��6'F�{ 'u(.� �#_gH��|} `��;tA���Q���[W�ugm�������G2#���ūrP`�;��^�"�h�I�p�
;P���w͸�6���R*
A�%�!��'m�L/K{ʍw	9���I�K��J���C���0�(�9���� 	�7t��bt�ٙn���[��Jx�vaMa"Z� ��r8tV�ӷð�4��6��LPx���+f]�S�9g�n����-�~t������#si�M0ERf�k�N�$�GL [{+��|�_�-�})$L�����y���&>��a�����inZt���r���)���CY60�j��^X��0<+����֥'2U�@ZU�RZ�_'�K�D�_g�?�efF�����T�FTCU�8�F��C��'������}�H��,1�$r;8r��_k�7P|o1���뾝��*ςx�S��=s�S���0��)I����X��?u�U����&������B����+�n_D�7T���_ߦ�:;7"�ښD�ofn�"{uxԙ�Z�yʉ�8�E�Y.��g��(�3ޖ��[�V��m�xÂ���\����E�W=k�tӁ��7GE )B�|H%3�! �d)����N���y��cr(3�|����V�[��	8�n��v��g�/yb'U�؊ �&�sO�e�d⨇�|)D�Z�����a���Th��U����N:��xD\��{�;�%�$�/oGĿ�y"�4>���׶���	�<�«��<��x��\��w��//��^N�jVU��[��t�Ǔ�\��DL;�G������2���,���e3��yG�Gũ��!���k;ߝǖ�v/�k���+	�#����L�����S�5v6�#���`�� ��q�&���^�X�GDG��;��1F>�`����z~�Ϳgj{(Q̅�E,� ��c�NK[Cm�UJo����vF�W�'���xg�$��N$�K�jΐZ��U�N����M�T�kۊ��*��Y'bI�Cc�+$_O��Z���TҶʴ�DM�L�α_á;g�2��(*���W���MY�EaFPE�[�)�D�k�V�;���= �T7�,�����Ic��LҪ���
�3�J�z̶�{}��Ov�"�Qof5���g�c%{5�d�>@�Sn�{��;n[� �%�l���h�_�N��Y�T?+��J�{���,����u.c�H���E�e�6I��˧���d�����L��X�+�q�L���,~|�;~r����ȓ	QƟ�Z�	�����փ�'��8�x�����^x�Kzo�j�i�}.��{��s��3,:��������%�ר�����~�0���Š�<Q3K#�Uif32l�X���R,Jy0�se�<Dt��K�/�O�^ _̘���g��o�+��A�m���Y��e-�1�	�7���!o*k���Pܷ�N~��S��U�)-�!o��4���|x�^Hh}�d�<T�Dwp��]��e<�t�.�����nlm���E�u.�:��[���Gi�Z<���H�{�`�H�f��iI�rG���ug�o���C�ss�W"E�ō�����y�WUj�µ`�?�%"�G�NUl,Axv��`-�"�sGBy^L�-��Q��&�ܶ��´���"���X�*><��Q��u��ep�d��ǲ�Aɔ(�
ʎ��Y�+�na���w�Qe��;�9�W���:K�Ζ-�-lpMٲdHT{��/��EZrM�
�HMo�[�HG���K<���"79�=�[��ci�
��@F��@6qL=4B-B'��q��ˑ�u��:7�P�v�Yh�jGxN%��ٲmP��Gg$F���o2��z���k���UQ�[ck�<a�����f���{`F��Fp	!z�y������B�g��[�
x���2�*�f��O�[q���_П�N�6�_;Lp/f`:�7[�'fe����s�#�,1���gJ��N�N���������O0�C�mms0U;t��Ք�ﶹR/��SI�g���:�e�]SP}�!���*t�ʅ�ox�O$d�"�y��[��J��^�n�R&yk���W���4Q���?Nk�'�I�n�𚟻)Һ����N���b�B�$���/vѥ������<5�b�*��l�tz)s�q'K����U`��Jx��o�c(2��@��gE:N�k��ܙ����(O����!X���������'<��"��Lߝ�r�`�Ng� ��>��8�\5=q�ŝ��;���5�7&`b��H�pZ$��	��9$�x_��<ۘ[�rȃ��ÔO��jE��������Q�ӈV�"Z,#MamCo�Jq%&�퓭Bv:�.�ڪ�a)����	�'ظ�&������FN�3�˨e��[��S�@��Բ��9P0�|	��9h[�'�V����fϢH�W0>�k5�+�z�P��~�%q��S���b�<����3_�/m=���jH�)�t*S�Y��$F`�y�/��-|faq����7I0@��L������Z}�<W�c,v�ȿ?�q��%=���=��njBv.|�q�vϱ&�T�ov�}�VW.�( /��u@D=�n7��-QҬ>K������\�����YE7����%n����熭*n)�#C���Q_}��,~���O��6���ԺBv���<�p�,����AE�W������'$��cF)�NV�wi�e�" ��L��E�������gwV���[�u�*��<�dr�y눱��1�~*t-,��?�xa��G2��t8&L���^�~8�LB���
�
��S0o�ꦘ�=�Tz���ѿ�u��ҩe������Z�=��8��g-���ZG}�g��\,m*��s̀Y[~�I�|��4�"J~��l�����ڛ�'h�����t��hyW�/���[��S檾�3_��x���Ĥ 	nP��p2�V�ӎ������
��1�t�aaσ!������)r�Ɉ}��F"��
���+�V�������$*�Tҥ��˛�*Yt�\��A�^�_d,���`<�����L|ʰ�u+|*�8i1ScꮟX�W�i�����:�H5��o�·�>�y�1�� �[��䳅���|.��} F����"*n�;C&2��ڳl�d� �d�aՠ⩂;�����ث[��FY�J��v䊟:�G������g����I��w�ȢB�!�ZA�!���q��1됛
���C�۲m�'(BL�P�Qek��NƎ��E��[���K>��]�#` <���� �K�o�p%z�U��Dq|-
lH����Q�z�>��>�8��o�c���˴�\F%���q��������:��!u\�2�;3s/Z�caB���M�'��e��6�n�E�%�p4�ҭ�TFh�#�W����>�譃�Y�+�~�V��D,�� �{Ē����Y�!�f
�������i{���Z)m����'|D��ގ�*�)b�ɅE��&;M\���U�l�x毠��������RyЭU��+5,ϋ}��I;7 ���V��}rҘ������Iߝ���	⻾��UG��p�pdL!z㧒��vݱd����9@�,`��!kd��`�%���-�OX���.x���g�S�賾��\�[���^s��hq��RUL�w����֧��� �wvЮ@�c���^m��\8��?A����=˿1�ǥ �����
h~:�1��wē&l��ę
m���f�)M�=7��.�*f������|���,]���1�C�B�3m��B�?����9��A�j��Ә/�zh���@Ts�0�<6���qmt�!�<�k�I��17FK��c��\ƫ}7��O�����7�C��W�N�L��������N�����%����Qq��ީ��o�U,�l���C�z�9��"l�rbky�^j􀮟J�ؗ28��J���<ɫ'�_���3۾�h���y��8�V��%����^��8J�B���T�	O��搑���*��ߔu=���uM_W����h���*���:�g�T	m�YDi�;�v�n�g��غz�eDs@��n��'z��-+`����'�������͈34�ZLa�����R��W��{�r瓩�@�Ԅ��E+��xw�!���ү���M�P�?���7��4!��A����,~_�0������swm�����$��K2#��2	�  	8��|����c�Lf�]_����N�Y|PRI47��Q\w��p�̼�E��hT~�a1n�sJwU�a�>fqE�]�Hk~�[�/�7�ԗ�7�9i�ďs�슛�Q���,&,,�Õ��T��!��[�����"M�u<p^��Ś���<��r'���,YFt#1C[_�*�r �Cױ�a��4��u3�)Yˤ�N�s�Ix�#JqiT�@m�m��x[)^�Ü�9��x�}�d,d�:�q}��OA�����P���Rz�Д�=��+B�*[�S�6�fc,�e���^K�������g��g�
x3����Ӻ�K���UR�œ�>b�S|&���j��9����u�	��,~7�yOA?�]B»А-fʡ�|��v�m��"���ew;�d4���	P��\����.�$�{�� aבu{��d!(șG�z��E��絺��G*�|�<��|)N�.#� u��c�iO;R�O�d<���ǖ�e�黒�|G�W0��	qg�.{Y6)�b�V�X|�#�@!��`P�\Y�!P�@R[���(�/P,6���zF�z�h��HU����Eל�e|������i�_���'�UW.��1����wRWA�rh�aVUꇟ�B��x.�AC�ط}�����	�b����k�t"R��+�(�����Ə5��1 �=��c�K#ľ0!�݊s��N.�/�q'��t7��7*��;^�J��5�r$�~<i~�������ujH���8�؇,���D�ݏa�&��Q{#
�A��_ O�(���<��;,_<��?\.���_� g����Rmm\��p2��������`�
� �M`��Y��oBh[�d/i�	��Y6���u,�%��k�@�W�Ó�I���˼-z��R�&��!� l�S:��GX�ak� ��ݭ;��#R�@5
�&�m��J�`��	6T3��m�6B��u��/47�/i�r��w���mܮ(xO�D���LX��l���2Ú�%`E��+�ݙ!]MU&�,6��Q	A�A�����;4^���҅��͸�kh���`�i7���R*��=�TסH�k��M�����~���E�P��`�~MK��xqI������t�"�7�䝕�XH�p�;<����f��3v�Lw����c��j�NV3����&6aE-�յ�Y����~��<fU���D���c�K�����Tw�+��,5eL&�����<a#��?�aZ���� �&�p��ebD`�������U��� ��H�&Dü�Rnɵ�m�"J+�Y�,%�e�nk!٭f��1.������B���{�(�r11�Q��)�󸮂�hu���oˠ�G�j����jk�˴mc)-ޡb��Ξ�6��/n�u�#�����'��:,~%�e����G"�˼[Z�֙�%ʃ��P|9�U�}��;��Q72^!����$f�K/\D���r�մ�,���$��k7!����m�D���;���d pCIB�ewCz*v��{�t~�LXx(�J��}���	�6u���T/{,,>eIj��<�rPr'8��Zb�(�6���Z#�`����p2;��v����
��>k� &��Up�v�OU�O%pFS�Z���M���t0�qضk޿�_�o-�I3$.^��!��M^�V�7�y�x�/���-3�qr>f��x�6�(X{��/�a֬O�O�z�iQP��Z��Zk�zDRΟV}�^��O�N(`?M =W���t�]ߟ91�S�;g�R��y�c�bHx������c@�Ig�_F.�Ђ��T�J�/_x�xB�^�lG����.���L(ͤ����&�I�E���P�s`Z�p�z�N'i�ޕ�=�
i0S�Ppb�RC ��:  /����cD�wh{$��*��e��ҀO?�]z�-����D�)�����A4
�2�ڛXm�7�S��[���	�\�M��y�����x��_atH��z����af�f�����Ƚ�������>�{����� ƨ�lq�<s+����*�v:��%CR���%�B���">���/U����dwg	w�o�0� 	9�G*s^m�.V��~���|��Ɖn	���������>�
�gm��
�a`���2�m#Х�s�̬Z���/RA �]G��W��gـ�ޡ]���V�̄u-�1�����%V�W8F1H���c�)^�a<�v��H'�j��l!�Im���Y�����_��~�% �>��I�{|��p��+�-h��AS��󽚿��0@V^6VA���rWq���=�&�����Y:)�����!�d�{T�����?HT�7��"���ķ3����4���(�9nl��<�qf�	6��M1��p�&h��*NV�Aq4!�J�ݚ�`�ޯ��MS�����5�4�NU=7>�뱈�c�!��o,*��>)+z���Kx\m��|}�FG3�$ώ��S:8����c�'�ᦋ�6WƟ=Kw	��Z�����%������9����"[��h���! �'�h3��=C�;�o?�H�p1Ntj1jy��V�7�u�3~,{�1�A�����Xz�|B^-�(�T��)&C�/�*�V��'dW��g��{4���uzz��������3�d*A�?�?�]�`?K���u�$�EPi���-Td������%'1��t?BF�x-����ydPo$��l��,Dd���@��8�l�ˁ�}wBw��K��������3=ԛ�%�FH�9�5ѥ���\	`{���X;ZAnh�C�w�Kۅ����(�k����)�m'y�*	��	�B��GM5ȷT�+@���G�i�rB0�F��%�ğjM�F�8t�_ֿ��?`j�}^kf���f�{zo���?3����2?�-�����̡8b"+*��Cs>�@7fz	�XHCȧ��x2��@@$a��=�
�{���7��`�0�cD�J�Ę[B��״�����W�>���BR�vI�Yk}ϩ�j˗��N<�yR���L���Sr^w�غ����E���A��`���|:��(�Ȫ��#ȴeeܾi�H��0}86����g}�}��t����:$w��h[�P��6A���$ա"RyH�y��M�(�c���4��JqP;��홸����v[<L�����IQ�+�@�p�<*4���Z�^Jb$�u�~�ב�i���� R2�����8ˬy���s7�����B��t�,�&�|	��C{!�|�L�~�jq	��)y��l^�=zGo� �����˿Ʊ��(U��� K?&Q˸
�A��|?D�M���Hc�������+�^�3���"j�@ľ�B�{�N��e�(�1c�)�� �6��/ɜ-'���� �2��^8R,S��V4�2rB�(�1&���d�J��+�W�9HX���{��x�6����FO���LR�N�t� }�g��tqE�pAO�|E�cr>m������9�DR��ȧ���/���K��� ΎC���[3A9�K=\���7ԿL&���Vz�'C4����z5��)�m{�s�_�m[q<C��"�4��Z��ZBQ8����TJ��;쏖G�OQ1���C�Q|�e�2w&Wm�=��[4���dO�p��RA\�\�0�.��i�- ~ZkeT�?Ӏ!�Mbـ�I�����K��d��_�}%�<(P~@i�|��5��y9�K�K,_���/�G��1��`����db�L��:�.��8Ê_�PHG��H8��^|�٢�ORjMDbݦˎ��oύ�qxU.�����rї=2c�b������͠��FG8��qּ' k���~!UXe@8_H¶T�|x9�4���N�{,���f�T=�'%�����PA�:���>�0iiU>�W��	2���z�b�I�AFrI?�'��b���O�&���b��g.�OX2�1jM��JZEr4ٻS�N�����V�>��-�6�9��������"�2a�ƙ�0��9f��=�ܓ�n��������L0������X���(�kGO�\48f�1=:���O\F�6P@��}��[�ڙ��ڦ�Z�n
/��I=υ�ȋO0�u]
������)M�G�z��6:�K=�Mf�Uc!J�"��&U�����q���+�	������u���J/r�!�a�DHO�iD	 ��fڧ���#T��ٹ��wC}\�{x��D�M�|�rP;K����j�A=�:�r�f�"��|[k��g��<zN�V=B<��\�j6��f��t��a˹��T~n������#3������Q�OZ,�|��$C��)5�����|	a��=%�n`Fn	�}C��YI�XÓ-�]���0�}���l���ą��K7ոd"�5��"h&]�p�f�8�
�:6��.=�I7�.����$��B� 1���$V�����A�@nom�Y�Z��g�y� rDޏ:�\��&xIw� �"%��(��v���s"y���`1ȠΫ��]� ���[���pE_�2��<U�lEɮ%=�Y7���/���$�@�y��p"�.b	�yҠ�@��f��x[3om;���DR3l<A�ʥ���5S�o��-�旧�zB鎋�GFa��s6m�J?�\܊%e��kw��l	����j�Kt��D�8|d�͇6���ԙ:�_Ɇ%��ƥ$DB�(}��t7Fu�=�ګWt|~t�l�? �<��E4K�_{��׹3�ux�l�Τ%�:���E׼e�s�ģ�&%Q���=���γ�r8��L��9
��sӘ�R�#,�-�"Ԥ2���
{����#�vF)G�8B�����̀o�y�H��?2�@W^w<+�)���l%-KΔ�]O�!�v1��N?����a��qZ���z���VBPNq���y�A&�k22i��8��KB�lO��FNh�
rS�H�8~���H�v YP����%���;�W�pK͘H�(�P�I���ݝ]!��Z�1.��C(;�R${��r��o�k��=�����K3�n��J9�oA���&�Ut����u+�3����������s]����"��W�,?I.8չ&����n�U�Mň�c��qb#b�,�����[W"fM7�
J���u�s�Uَ�[���7��ӑ����<��V�<���<\�a�1�����8O��zT�	��"s�ξ��ia�b��O�x^A���هAn�)'��ȓ� @���0)������5I��J����n�a��E��������S�G��;=��4����D߲)p���F����p;$@����@��
P%p���M���I١�Gx�s�Gneg�ωu�hڽ����l6Jĵ�@ �&uܛ�܅cō5���oR#�6tFR��"��<�oٵŬ�3�(hS�h��I^�);o^O��̌R5wŹ0x�\}"=/Ҙ���Ec ��z�$�_�8y,��K#�et�[�)�毙�VW�X��>�R�(��lN�Kyʂ���m�{p����$����&�g��O��\�+�ME���Cg��C!�I��_�S^F�G.�D
��H����yGbjOz��/I'A�RҨd����M��|�Y�ks��BՈ
��g�;&&�Cؒ�d����[/\��ɐNXڮ��W����<I��2����m ��K�}D��։f6X��;�J�tg��#�,_������$�&��g4�s��w��&���v�������PrJ(+��t\�m����lZɌ��sm� �����2���Z>'!1�(�9�6 �IK5Fn%���̅�����PO�5�@��H�;!�ۇ`��:��e��i2���㬘O�5��eۅV�Fً�k��3:��gC9uV$�&5S]4*�:;�����.*o��rZalOS-�_�xρ.P� 	��Q25�UDS�pG�Qc'�H]��at���ͪ�����U��o:Vw�|:^�����t����9� ����窇�uU֛�ף��ӧ��@=
`�"��� �?����Ѷ̌��|Ϥ�屪V.��	�P}23�nLu [HM��j�7���8j���ǳݩ�����P> ���9$f�U�g6���O��o_���e�+�e�w�;Z�ߘC[�h��u���b���#q�x�bmCD���i���V"��|%ȃ����)�s��� "�e��m/���K��w ko��l�`�8$xޫ!L���5���$��F ;���~-�#"�HmkP�������%-�Rl�s�KYH�c7��s���+�=1��p��N�t>Z<'_�x�t�C�0�",�^���y0%�[���u:uG����ⴥv��B
c@V�zĜs���TÑ����w�h�����
z�VFL(�SK��-�� v4ЏK�6g\�Θ���b�tB�o��ٍ�,�ӂl�{�| �h�W����<�R\T�r���N�'��E����;o�����]���QK6�넪-��!�۪'��h& YSbC3�ݿ:��F�C����\1������71��u�ȇ�=��h�M2���h��@�k+J����*�iא�m,�@��F�s@,�N!.�[a3��M��|A��.���A�&�z���w.R�����V�����:p�*c���t�iD����_A�bC�~&�?������T���`�:/��s�S�����m�wb��e��B�[<�Ne��0+��[�V|�(ʜ���!1����L}�pb�#�H'[�!�Lj_�<TS��鲝�Km^��[�c��E��B�-��Mi�'��]����07&�E�e������5oe��Ul��%��)U.b%�+q,1ı�u �f]�^Za�1�\zƜ�f/��c�� fn�4���ǔ�q�B�9.Q�;��m�,,�R�&�ikb��T|94�`t��1<7 ��Q�������u!�.j�|�D`	֋��_!
�ޘ���@|��x��!�̺ͽs�4��a:�׸�N��H��߼�����X�(~p��0�V�|��)��\e'�����s��ݛ�����r�pG�s�T�K$��'�I�(Pdj׻Dc�hI��#+�ޚ���?�����{/�`�w��� �J��I���,���q^rv:�|��w{������ӣ�F��+8v��?�0J${�=��Rb��1K�60?c. %�ߞG��Y�ǀ�n9!m�{�~%�Ir�r�Ugˁ�'5fbD!5qE���]���G�Y���1��"�H��|l�@��fe��3�;����E�X}����kU$�y� ��'��u`݈)�6A��<ye�����\Z͂�{�[&�Ӛ�bP<��v`�!,b�uO��yy�AA� ���i֡C�eE	%�Y����
F@�9��S<<��%�d�w�T�F��;=:��K�N;��`�,���γ���&�2Q�~�����v.��t_)T��t� dS���b-���d9����ei�5�����0�	+ShrH"11��Ȩ���P�o�3�	B�H�� �[����E�?��2;�m	�&�#�t�4�ƻ�Ǫ��E�V��7@ķ���{���u�s���ܰAS͔T�` ���'�7�cP)�e��_:���0�w ?�{=5���[��~�HE�T|]-���f�-%]��c�|O�V����S���h�
���Q�č�Nr�_�k�q����ȯ��n�xY�aY�U�6cX�\�2�K�櫮��P�W�����ðl��Ț�P��<���3ۨ��N�r�ݿ"�|4�F0�#��/�+a�'!��vψ#?���i���M6L2P�m�8jPZ�ÿ�o""�_[��:�(2\`T$���ް���P�q)y�z���Y��N�r��\L=��M	�Z���N&���Z:^�M�
-h?�Ke�b�Ĭ�8w��f��z�*�_ĶB.z���S�^�N�5g�w'
VL���⾑r � DCPp�t-�<�&4�ˈ�[&�����:*�qH� �1=��@�����>�<�g�A��AYsi�=0X~m\�Q@E��iv��t��-\���Q�ȲU��g��a�a 3���~Q���M|B������^�� 
�]�([Q�<�v�0��O�GP|mmNg�����Ĳ��Y��"�W��H���<G�S��e=|m2�ތsa��'��)x���oٹ8QAa�����"�O�Nyp���݁��ݷ̋�Q��_��Q�S��J8��9���/i��p9L��-����0�@x�y�̳�9�<@�+E�7���S��wV���Ź�b�-�̫s)"AQ�a���>I.�KVH��K_ �;���b��~�n�7�J�h�M���]D�/�r|k�?L��%n��'���"���P�}��I���Q��?�-H���=�o=��lң��n��^��$|�/K(�I�k�*0���ϴi�����]��}���(x��D~-;���[�����a�����P�9{I=�(�`�)Y��qD z#&��YxC��W�Qs�ۘu�J�A�0L�||�thK��!Pz�Y��ng�ǣ.6�h�F�/�;�p:�߫h�P��Á���{.���"s3���S��[�)�����:���w�� W��Sa4�D[>��o�˄i
�
�|(#�ͼ��P	V�+�-^��y�$NLq�H9&�^��"�r�Ukݺ�bhyiܯ[5�/EuV�|O1�b�я��K����$j���Hҷ�P2�u���zx�ݛi8E�)���k����	Pr\�,t�K�C��������x���Źf���T���t��6�e��I�B�JN�T����;�Y�Ȓ�ƎlPE���UJ{�@�����H	�މu���6��e,��(9]5В��z*^U��t)ar�1*��ظ�P� -�VL���-Ɖ��r󛐠�>�bK/X��,�����H���C�H��[��9�Tc�D�
o��^sF����1DZ��5���l�.���p+��k�FFq�����r~\Pζ,���/�3.%�� 9����[؂�T�F�x`qY�,��>��A���"4~˄tO��m㒺�
�1��$��e�8����'aR�jS5�揾`@��0R(p�Tf������͊��0<h���P�/k����k��Z�3��v7��� gb�WB����wA��k򂈒E3i��~��bߴ:��.�#�*>&����g�1�FV���5'��InD���~�N�mq*3��
p���͏VK3Z�
����m���W���{ D�j��_�v	��Tk 	^��f {��������f����H���%�a����r8w�FI�b��V��F��05�+�&�����|J��m ����`�S�SX#�����#�f���s��0� cbq���paVh�����u?"��O� %����:ݱ���嵊��$}�1�]��8�)�ۖ��`/�
L�Uз�� n�dsѿ�9��QqX޸J�B��=�����l�%;֋pwB6��by��=/	�e��J�)�y����ك�_ŵP9;X�`��KE~��%O��j�������ϒ��m�z׵(5F�Z��q(Fn�x��?�1E�ZG��؎*wX�)�6�1v(��/&/ ��拽���2Zzk��̄�Na���M${�ސ)pY�Ξ�S��5��Ep�b0�pʜ~�gޛMԇ�f����_�AC�n*[Ƌ�n[�8�����9]���X!�7�*��1 ��c�')sÄY�Z���6���K`-CP"޿�qu��ϩ�	J.��Mq�ęoIlD�,�kK�)�����%<�*�i�a�iǕ:��3�jK!�/��k/r)x����r�0�^�&T貁N�;���IV0����D7%�=��؈Әa���~i�Uq��d�N�3H	9��G�Scĉ�k}gHF+�������8�����ޣ�1�/��������.Y��)��Æ˫
s� ӆ�E��;��5�^ȶ�����!l�pʊ$�"K�E����p�(�s/��7�Vp�"�8��~G6��!aG�i�+C�ɗ��=M�ᩩN�c�l�XL�ه��MV�{ r���ъu=�#���,z�!u��>`Ŭ�c�׹qI�}�U�No� IH!��;Y�9_o��lM0���Ja�ߧ!G��(/!O���W����GQ�
R���������^<�ZX�F�迾�����j@����>�h����[Uc>�����#�������[/�6ށ
�'b����Y/?O�7h_��w ��ÝL�4s�L�nf�X������*Zc�C���ku ����I��,�K#��Ԑ}�Hp�2#��L#꿏>f%�B=b �	"c(fns�� �6�-¤M�>�cY�W�#e���g0��J��k �Ch�^<����ܞ1epB ��<��(��nu�cjN|���`�y��߱A>�i �9����u���j|���6n%��1�)?E�� �ٟl�Ut�����?�2*���VX�Y��m�xp�g%�g��.�b�JUf���pj	�d
�ʵ����I����U\d����&��������c#��0�)�󞾥��bFP�ݷ`cdM3��S��rR�S��ϳCY�T/>kҙ�l?�oϩUI�H-�a&�d3h�s��њ�I�Z��	"f2ƿщ�!��5��G��&-P�N���d��I��.圀�O��~��:2޶�1I��v�^Fx:��[���O��!�q�NZ� }�h.�9F*X�@2�����/F΋�H�K��U�R,E#�1ps31���M�=��ﭾFS��D������_��̒N���;�:��XP�9B^���O��Mb��_ו�3�{:>�����e@(Z�w)�f��Z*�*��k�36XK�����$�߱Ͳ��j�̤I*������֒�b]5��$U%Y�)��#	�8�����70��/�-6]u�� ��M��M���.\%`�Nq��L�Հ󑷨����� ��Aa��U�Y��/��FL�m���J������^،z������j���5���흲�;y1Dh�N)-�ɗ�}F�����;Q7	�uɿ�)��'۱#{B�^j�>P�A�V� :�����F!���.�k��՚���2zy��gZ�a/�g4�dg��CD�!���YHF�^H�I�5����Cuh�_`�� 9&0r������-#3�����Z40���I�^��i��d�| �w����p�{R�[k{hY�G$6��'_��c5;W��9'E�bo��[M�D}#@5��}�8Z�I�O�4[�ZD�;����)�~���[�A�؏��$ aBl��=���M�����w�&HZ/ȁ+���-�q�W���"U�B ���'�Y��J�+`o5탺���}$�C�����g�%��� I����r�tū������9�������,�U4/�H��ҕ�I��1���1�{�3͡�����TC��j��k\�S���R��hH2�:bx)͂�QWd��aJ�C��
%��5/��O�S~�ⷼu�C-�n�a�¯+�H�a'c�����b5��_�7�T�����'OU���sl�3踹��q��b��:ܘ�n۸�����cjn���f���>7yG�*�E<&5[�c�e���p���~t�?�L���1r?,+�	m�-<[:�߽%�S�'�4��-Q�\B�ܥ�Y\n<��Y/Ʈ4:�R:HID�BgWD����W➎-�����a���C������+&��gZ��J�!o��3A䮘���N��?d���%�R��	�A7�i8膓^}*����3w{G����Jf�Ѹ<ز�ǡ���/�fg��4��Z�� ��t_���s/�\u�S��~��Z�!�X\a�4$B"��" z-��"+7+�D69�;���)�i�1���Sʢ�@��Q����T��0����p����$���_,��{�#�ȕ�WBw\�F����)�ե��Y���1��;�4S�����פ���H��u�n�K��n&�	��}p��Y���;͝p�:�UY���89�SIYMN��E��vX�F_��tK��+�l�H�ɡw��j����rI�h�R�?���wt�������:�)�X��i���̓ә���zG'E/��@D��z�㆕�9q�1�8�������68R�H8���?T�vG�}�pվ&R�X����`2Zb�g��ҡP���{\�������!J�D~�g�;��J�>!��`Q��T�e�b�,�U�rR��VtB��R��p�0�m�J2:���蛋���NZρ�%�J/���ke�Sf��Y�8��?�g#�Uy�,��r�S�h�\�A�@�@�]ێ��XT��ɝ��e�R�ч�:���~;:EM��
f(�!ˏM�{9��+O���O���`d��$��A�J�`~W����W��ǒ��c4�����yϑx�!��P�B���9��҇��)o�S������J'�cG|��^ξ����+�0ڼ)��)�w~a�S#��չt�j��e)O�r���vp�tivs23�y����|G��ҕ��?8�~�EpsVP�8y_Q��'B8U� {���]��� �R��`ϟ�bjpw�4���6�]��Z���΢��i0dr�JZ^>L��2�	ڜXW�\%�k�+r��9���Z����=�*3	/ � �Vf�9�q�L�r9��B��I�ݍ���hġ�n�E�H?�V�He�~�N󜳘Xե�5;�0<F��8�)�U��E�h��肀!�ė�2��2�ː�]ά[/%һ�(Z��j������ʴ���'T�2���_D�G�%k+���Nhg<��5Qlo����h���W˵ ��,���C۲V����Kx_�Y��2.A�p2F���꠰e`�8�|h�!���G�B�몕�
(�j���Ć"Pt��eͣ��h�u��P���]x�]ʒ������}�5�"�Sz��Z;� �b�⣇�P�6���l²�s�^z}��h�)ܶ�>��BX4D�U�u!����O���.4�P�:�5a��_����P!��)+��_�K��  �ɖ�3��1��=Ǽ�ñ��I�R�s�uHB�x�c6m:�S���.��17�p��7Tn->�B�]+��)}��)-�����/<RU���� 	S
U��Տ�4'S#�h�T��r4�DP�����MVp���Nrn�km<�<��+�K��]#�4�?�4�*���?�G�W�Γ_�e�{K�e�hL-�l~������=ҕ���2�Ξ��_߳�dn�w���TM=;=N�R�H��2��|S*�Ёo=�_�>���h_Ź�W���=���B9r$7�.��}��|,�P��)6!���᫢wD��Tɱ٢�D^g��CMSY�?�C���z���:i���ݵԂa* �|�$\���7kf�0�% -0^Ҩ��Bp����:sΟ���?ǜ޻9�M�21�h��J�%���R'�P�sy��8��*V�rm_��� �$4��%�o��z�X�`��"2Uқ�l{w)�O+�]w���C�C��&]��������):(m�}x�ɚM��������z}2�u��R�'��*�UK�� �5�M�(�KV���t-�Ņi�#�A�"�� U�+��@����f`r�;�6^�w�
0l�I��j8��qm�R�"t�� +����@��y�t���v����zN��(�6
h9�#��n��&�A��X���P�L��A~�����@�x�\��UJ��r���G1��2ui������]˜r��GW�U��o&=%O�%�C7R;qO���ȞaU���Ǭ��[������c;��a6W�ġs��b;hʜWS�����9H�&�2�Z�0��]Y��G�Hκ|��j	7}��ܶn\�8P�
!l�zO����_�tPh/��^����Z�o4r��3�A1z�7pn���7av�h��'��y�Y �e��j�]�"��l����?A%i)`"��ۊ~3uc���uz��ܑ?�
��zG�]��M�2��*(�ek.�dS��w�*�M���MϲrR�.J��n.�gAKX��8�0��I�ϾjW�\��h�ݣF�_ˊϴ��Q�FEi4�Ȗ�B��"n��&�5z�"�����-Y����@�/iެW�ΥF�A*V6���I��ӗ��2�B��D��T���T8
�F ��9/�<�ֶ�� eR�@;������q�9~�g� Z�I��0{���:[=��,S�z�(\H �M��-cAxb�*�DBլZ������$�M�2__b����nU�B7|����;iQ�;�#�;f����ƠxG�Blu��
�8�7s�c\��OA|	�m�/m��4Ǔӵ�<�&��B����%Kzfz�̌ ��A}�C�Z��h͑�/ v��=.�W__ZФ8q�d��	���M��A�Bl'+���RDF���9QTI:eW�z�	��r�.m�:�3���"���KNs���ˣ������.��
���x���iJ�ƺ�z&'�9�P��y$b��|�x�*b��������QGo�J{������O��\rÛ�˖-&�ű�ae�"�]@�2�=��UYWG������0(��z��z���B�*+��i �;�Rg��$�6����k.��ϴt�A\����q���hKb潫ѱ�d!= ��l!,���h�/g6���vr��1�s��`h<�Ϭ���Ը��������.&��cL%��6�	�����FCWX�2�~a�_6�|6'�jB�b��e�CJ��D�C��o�,U�x"R	s��tn���D��=�}hK�����,�y�τ'E�n��Na�e����!�_�����"w��v���jN�â|L�}-8��iPV���%}��.�2�-:sd���4����Y>݌5O�yH�î���]���X���̂�����Q�2h�?�Y%n�C���g�!cEII�����x�ֲ���'�~>���g��a&� h��G�|�CU�9�%��rN4̵9����.渴.psT�V���l�^�v[*�$zʚ'u7Lয়)�4��Z>���m��o���o���vƞ!������|���:�k��OFq���� ��C��GK��!
i��b��&q.c*�z�R�ch��������'�o+̹��>V��C)�N|͝�i�gYj�[�������Z�\��P��g ��s�d�@�!y�Sñ3��5��0�8?�C���3���V��!�7T$��4' �R��[��	O���o=�X�\�pb��b-��r���ⱳ(��4��~� ȭ��
^�Sqsg��[�lX��
Ίib�Xyn;���W@��6�w3?n>�����Z'�u_���,�&����>�+���U�*e���"�o0
�r'�r��_҉Z ]3ʺ
Lψ�B�o:{ ���{�+�2 Vf�����Y�*V����vB��u�X�B ��䅗_<�?�m�����
��ɫ��ؾ�ON�Q�9/d;b��37I6Xް{�����v�w�u��x�{dM��et���~�X�
���p�)\�
2q5Բs�o��AIN��US�b�;I\�U�đJ4���ax�܃X�_XLP���{����,\�+l��A/9n�(:D��5ua(ل]���4W ��wo�1B}��%Đf�ЦлU u0P�c2�6l����=I�nH��p��]�~>���
L6���g���J���;Dgp��npqy�� DO��Z�S�P�.D�D!Ve2��ٖ���C����Q���%"(�Ʀ9^�7J�����x&p��+/�6a(�X�xL�H:����Bߏ��/�yN���?9-JI:�� �)`s��"���
.�2�Ea�u���S��Ӫ��Z�@�}���'��䐌����̫�r�?OM���WJw�����G����AX��}�:���0�����L7�+w�������/�>D��a��d<Di�ya�h�����16�>�R���=��w������~i����0qR+_���n�:� �Y�=��a�꺨i���Δ
��%�D��p��?h��s���ܘM
���,sf�ʙ���O�2���Z+����aV��	����Q�(�'e��Th�&7�4L��1�2�ի*}��פ�yxg��� �1�zN��47db'��1����f��1Ú�r�������=��jgO(���a���lTզ����
0~4��X������Ѥg�'��Ĥe�y��:�?����TT�29ߑܙu��#s8�._��֓N�_IK�(��V�\�a8G����iF�YNlV�kۍQ M�>70�[u��Qai��J�ب�����[�@w�N�z�o%��$��ߍu�d\�C
����Cq�5ޕ����f����������֯3ݯX��#=�T9ʯa#t���������^�F��aM��a;���&�(�b����~[���魽�[k��x��{��f�BI@�̖��_�Y&�<K��2'�\�ZW�5{2ˠ�yF�<M!+�l�?�	��̋��C��Ttg,��y�\� 6ؗq�2�4s�>.�?�$�/���Z��mBi��a����z��5�c�uk2�-S�*�%M/�|u�3�e��bW���LT�m��"w�z�lJn�n	}U+����D�;2v �G�sA�A��T��3�l%��c��ٹ��}_>
����Q|�h���DQ�E���b����q0��k��M?|�'����e�B�B��b��,� M�Je巋��#
���[#�R�2�2�>�䬲I���1У9zJ;�\��E���3d��5ш��D�P�����C4hUUC�7G��T��J��� ��A�0g�������%����|g��8�RՁ��よ�]�p�Ҳhl�oT� eH�kO͝�@����If�5/��F�|W�Lu��"�*L$�S��5"����uϖ��P��D��Υ^}klp��TWMN�4y@L���vI�q�}�e��B|�;d�8�"3;$�㮻!l��m��$��1Qע�5�����)�������O���
��D<���Ɨ:_]R�$(L��!q�BH e���w�,h'-�}�qV�h;�����[qͧh�]&s㓭S��Gr�. ���](�pp�a8��	]� ��;�ׂt]�2�$�KkTt�X|��\E��tat���K��;��xm���YM%w��!@���A���,�r��K��ߢv/�d���H�>�}ȹ ��i%�=gfE`+?$9L/��� db����	~�Hr�X�t�5&�̜�#�~��Q���ą T��6��]������ϠOH��c׳�ڀY�!��o�\���1��U'��S�!p&Cu|8��H0	sm'�@oS�s��l&�*�,���m��ohf��)m,��K�������*�����	�ye ��X�/,��%�����P��@����8fN*��1z�u���wo�Gh�:Ii�ܺ�jW�Q(��,��BMu�/Ց1�Wvηu�A�w}`
_fOz�j>����d�D�)�l��3B�_d4U��w�P��
H����e�T��_p/3hZ�����.<��
�|s�>�3�0'��-7���♧����
%"��4O ��8���-�ݚ����	��ǵ��(yIO�����ɟT��'��V���ZM9���|�O�Ӥ�7H��#��>�=���P��x�^(,��xs�O�x�����[R$��;&�[��#JdϠ�؜y�Y�χH��5γ�R".F~{T=�z��}8O ���i��+Y��ek3��cKI*u�����B1En$���{8�N�3�)�<�&#cC�۰`��F��I�����!D3~��4v$R#��*9�Ň�o�Vϊ�E�\Gr>��x`�\��d�صrN�RibB�t�D���ĸ��'�v�b�Ԑ�������0<#�p�ߏ~��Q\J�K���IN��� �Ӗ�����y��Ċ7m&�:�?\��w�H�+�,�P�V�Ue+�q"R�)�m��S����V� �'�`��!�^CV.w!���7���q�/zG{©�zl+p�g�~�'���6�J����0F�g),��;p:� y�{�Y
B/�0d$�˸��GkԶ��<e����x>��{�	�3�:,@���?{Q���1��Ur+��S�0'�s��x[E���ǅ���!�Ƥ�kl�pB��
S�ƃ&�X�Yd��4;J �y����\A4���n��Օ��A�&۠��Ad���̩�~˛S����t�a-Z�������F�lU̙������AM%�6aBj�[kK��	_�˙�dd3��O������(E�,�!h`�.ö5�-��x��!Q[}< ����r�^7����T��$ޤxݻ���K�|�PlE6�P����bSısz�
��X��6��@�%f1I8����R���w����t�7�>�`t���~������{�*���7�K�@�n��J裭�8��A|��Ƥ��r�,���/��z�<&��ԭ��I�d�1H�����|�]XJ9�wlIR���eu\;����̲�o4r"~~_�=3��>�F�؏7Չz��P��s���Ց��3���9б�7�pl�Q�{\ߘ�HA�#��{ڨp|�V�[yo����A�/�����@X����@t�+��i��VJ������-�Le�� �p�lT�Z�)���N�bd��ԥS-��o�`�D�4[��zZǅ�Wc�V�ջ�ˢ��'ԙ'W�q9ȼ��ϏP�i
˞���E0��vo+�/ �:rI�#upU>�k7�d��=�y
�ΖC�l�J���P�2Ż�ط%����=��J�ֺ \�/2�+Z?H�Rv�1�m#�mM9*�M0ҝ�7ͨ��ܼ�.ץ�n�Sp�jz�`-t�?��H��u8���؛���Mb�Z@��RӨ�?d>ܺ��=u;���@ٻ.�� G��v����^ޫ�U��c�k�3@J�z��l#e�W��ԛ�g���6�w���V��=k������Ox ������!s��!�ʑ`��+ n�`�D��E�c�s@2�G#H��1:��˵�����H���m���lZ�;DB�w$��#?�
����3��B+�j;,��7�kl�[���$z��-N�������I7t(bk�e��
ba�<5�^FYz�#E��~}Eo�1��R�F�MN�b��#��M"��NR�Ȑ��.�=�%pB5�Z��Vt8d�X�d����s�KS���!���8e�/O>�^�xh��GE�V��B'�9u;]�3�*���O�6��^��o���9��;���9�"	ٽa�E��Fߗ���8֌�J����2��¾��A�ʷ��f���	�N*_>��߷�9J�;,�T��N���|���ݴ��l����@G���>����뵇�k^LM��ɶ�?�)�UH��*i�W���H����S�����@�R+��پW{Qpgv�'��؇ζ]�Y��EEC U�vR��|��	f����Ea���췈B�	�sȸ���5��Fv��-���0|��gP��1���u�l��e��D/K�|<+�qU�[�-��K�U��T$�C����[��gl<�D0=�_OݺJ~c�R����1�� Ѓ~q����.?i͎�n�NMg�%_�X��=�[�ʆ[LY��h�
"Slw#!����$�5���I2�.㿨�3h�7�����)
se<-�CNG"��
Y��T޺=��s_F~�qx����I��X��Y��/aԔ�7����pg�D��`z�d��&�pU	_!s��4gQ��;;U��/��Ѕ'���&0)(��h?������D�$��4~IEw!��f��Ǫ��$�Hw��\��F�ƽ�G���w h�v��NَW5o0�J7_J\�	4���z�������Ԋ��3�G�g��>���D
b�$��[��ik3�f[]��T��9e!ҀQ{��a>����D�2�4E&��ah��6���������5�)��[t��j�9��+	��A���}Fk�V!A%,b��| ����Қ�U	�;�fD�h�-#��k|�$vr��c��_�k��	_����h�"���-"Q��W-̚�yI�K��15z��Z�L�����G�x}$��N��H�\�����uJ��t^Jie�����qb-$���o�A��#��y����:��v([�G*��:ԅ@7�����8|�U�W��b0��c�"���@��i�(�)�b�k���j������Ԩ������n������C���]�J�XyO޶�w���w�^�o��su/q#�PӦ�l�xdM��<I�-����`�m�J��O�?h�����y����joc�s&f�{�0sp�3fuuwm1�v������`!t���M�qSis�+����JGg�\n��!��k�o��>�-G,�Ks��HGeI�G�{rvVb�3)�m�=�>��pXkۋ���i%�8�Ў��Ex�O�f����<8ޯS3�IXM��\�hYS4��:+	恢���JWY5�⎩��繁�|�iks�5hŕ�R�#H/��XI��b�[�����gc�>���UGL�pm#����i�p�8~<�Q�du*(��c��D\B]9��Jn�tn����]^��MS�-Խ���.�=�C�]b�i\_T��bڽ��;M��4�Ҷ%u�9�G����S�f��,`���͕8�=�PV�75��e����^���a ���I�h\	�qY��H�ʕ0�<����Ыy�{���gx!k��e@�;���H�z0�=g;�4�ƒ�"吚����x-��,3��!ΰzԅ�,��Q�$��H���E�2���ڣ����*�^�\���)����l�lħ��! A��ݹ��k���*�(G��$�ˁ�R�
_�x��o���^o�`?���1E*�Μ,j��9~z7�_��5�1
��N����Xk3��_��(�Et �dO\?Rp ̍��O!����L�91Lr��>�&�� q��S������񗍪h�.�=�`�T� Ǣ*�:�f��ja��?�`���PJ��.��9j\)������Z���l��rƻ��H�\�e�Z6C$#�69ES:T7u/�br5�����2���[).ﷀm�D/։�_I��r~Y��'�DDpL�Mio(�^�#�<�cA_E��d��y7�)�[���$X���K�V�! �L�Ma�T�����.��,a��ɐ��6D6��%|̬E��|�MrI�[xѼ����R�V6`�O3���|�E�$uA��v.�sq?��u��/꿛[E=6$C��c!�����U��/�X��O4���ͩ��˲�A��B�yo��m�E�ݖ�V�~��@�w�NN�� =-��7�"�	���#9�s�B!�9���?ӗ0��0�4|�Z�cg���+�j������ˣ��	��ڋ��֠�{�"��yz���QP���ߨ��6�j�Tz�����8��1�DT�\BqI0�v]���V��L��d��lО�����C�����ԈI	'%.�p��'F_/k5х�G��I��a������(�p����V�I,^�?}� �&;��FKU���F�%o�6���I���Yv՗5��)��l+�T���fW/�&!z9H~َ�l��s˪���;��M'd��D���� ��F �,הm��#@������|+�;��+�nż�H�G���ڧO���)��}.��ꭏq�ђW`b�CQ�GA�kV������:�U�e��a�C�{$X�� �!r����^A1|k�L��;U6�H��z��ј��Xb����M^���[L�МJ�p3�����q-���dː�x�dpK�Br�v�x���W<뾹�.W'��WC�űEP{f�ÿ�$bӸ@栩z��b���H���u#�p��a-5b���E�3�J��s��%�V��S�D���G���i/W�n#���{�8y�.�97�#��m?[R|l�F�|�L��?d��=�s����d����B[�	��ڐ�����͙g�Ϻ�+��~�A�f��/\�`�8�Ҝ����;æd����ǭQ�n-�s�K�2c�s]�knԿ��'�:^��D6�rp�99Ǳ-�nڴ���͟@ϫ����8��r�%"��0	l�TU��_D7->�J(�@<�\6��	�5�OO������P����D�ns��&^}�tx����7x�"(��Lq�h?i��V���X��^+�O��J}�0yЯs�x3�R�0�eqQg\�7��l�X]�oV�c��G<D��V�M�.a�E���4��A�� � S�m��s�`Y��r�"�ux�o&�/�W��b�kb_w�%'��"�|�4	0�}ѝX�����?{�����Nq1R�x��D���%���v}���ݱ-z��,�/ȯ?{��]��S���-)7��b`���|z+���+Ą�S��.Laս�\��Mȼu<k��[��� �IK�V,9)	/[ʠ�Uw��r������$t��Y��b�+I�b,��Ɵ݉��ƂC2⽓�P:&ϙ��S.��N��wG.3B:���D5!\*U`-�b���4�&ͣ�}��?�؊�@_���D��2����0;	�@p�������9i�g�c�5� ��JPJ
�Z	Aτ|��Ц IO�k�/�4�LX�w���OpW��n���5�$�
����[u�]�	�R���7vՎi����!�?ev�bc=LS���i�&�2�3��&{���x�1����z1@��$^�j�������A7��?]�=�^|�MB-�>?�RsM��&ð�u��i�vg؏]�4��z��|�����27��頉7�묋�|�?���\�+>G7X�t~ɤg���{�����Jr��y�9-C�#̗~T�|ۨR������,�KǷ�������0H,fH0p��o��R�x'�/F�5��WB�)�n�.��$ϒ��/�2�C�!Av�C��<��J��=���9��9���$ o[29�� ���o3�w�;O%�)�-�f{e)f�1�^���b�~�m�EQ{��bO���r.�0U�NT�ՠY��M����L�W1��	�cc	k%ua��m����X}���Ǆ���IHc36�A}�cdM���ѰX4D��T���ebuBHi�Yjy{��8V��J@��%ݞU.��b���o|Q�Ǆݖ��@����3����{����-��X(��v��JCF�4㩤q
��W~�@��ogBI}�.zcA�r�m���������.��'p	򯵶/��H�]b@	d�)�W�R|��.�\������pSS��ơ���'��	�#P;����ƕ[��'f-N�U~�>���!��
V�@l��DB�Н+�#XZ�V1\ �&��!ɛS1��U�/��R(W�DJ��KwJ]u�z�cb?Aی�n�)7I��*����^��Bz�����kц^��\k�R�x�����"T���˒4�,g�'�>��F���y�[�]Ҭf�V���=���D=�4M�/_N��@����h.w��܆u�ীd.A���\ 4��
�;��ڪ�' ����PD�ȎZ0l+ '��E�l�з���r�5�귇6�Ll����"r6���3=�
��:�a蚃���};���)NU��{�V2LC˛�t ��&;WW��枑��xK�D�L����G[�L8?��<}�iz�s|�*���k�~��BKml7��}ɸy�����̖R��d�K�+S���͔j�i��wS]v���|21�Lq<TH��W�(�sx��M�+Ɖ��5��a�� �k�V}�H����ԓ6AY֌Pb��KƘ}�/����R8�;
'`�$����s.d�f�o�����~Q�/|By4F���eC�2/���9������h�V�w��RH�\/Ow�3T��-7e���k��� �|d�Ǿ�=���ʆ��w�E�Z��zf���To��р�`k�'�8����~SoXM
���䖗��f�QOB�Dfwd$̨z�0�]귱k~�3�8�X� �%�F�HAm���]��'@M�[�����xY͔�9��
u�5��N�6�!����+,����k9�T��Zi��j��0�4`��L1�zX��Ĺ���}q��?��**U��ƪ�O���?��if��]`1@�#�]j��1�v�i���+p<S�1n �űv�#	� cc?��F��'�sJ*�g����K�?�1FA�@w��Na��=���]Ux��M:#&P������I�N�#֋@LGm(i+�����s�A�xe����	\���,��	eY�bE�Ǽ!���/P�`z����g��p��1r�5�C���w�oɉX����O��ф
c-U���@�zj��:��1,tW�ٓ����!��$�v$����N�@�Ƕ��^A�-Wm�t��Q�9 *����%7/m�YW�R��r]pe:��g��ˋz��fX���>�A>���1z����n/��|���z7��NKCz�X��-��.56�ږ�]8�[�����S_lDrA��Mh�ry�KX�����
�J�[t#O�_���!$f�s�#=9)�k�k1���@pD�y��J�˿9q�e��R2�Ǽ��}��W� �S��wh�bG=� ����c"�v%��Q?���� ��mY0�4��nzè��WN�qܿ�f`Yv��Cy�(48g?j� <�v�IV�#�Σ)S�e�y<�i�����2@�U��w�ʭ;������q�|����sZ�]���L��U�8Yj����yIR��6̍B�义AA�!{�>��?�f��VP̇$�F]bʯ(n
�l���#�D��W����|�������CM��FM�J%N�f�u�|��V9�;���6�X��Z��x������G��_�����ztѪ���l?�����
.��]�¹a� =�7�k#�$Zk�^Ue��Z�پ�B��Uv�n�m��??�|yQ���+Ҙʢ�u�:r�֢NQ���A[�yI�E�����#ĩp=W�0�*YT
.ը�|v���1���ZK^Ʀ�����`�>����nXR�4�t�FG�K�lw-1�}˜��pJ�%kY��i�����4y]��f|L݈������҆]-��H�5��eCL{ટ��L$��$��;�H��I�]0���d�}�<�B���s��|z�h�Zy����4L����)��uiS	�i���cQ�I]�C7�gE啫`�B�b"�LN�QWfA�<>D P�Џ���*K�躀�J� \������>���u�������ojs�PzR]�_NU���6��72�J�`��5@��'sF���0^4�]NL��ԓ�[{i�
`
����k;�g���l��j�����Qlc��k�oc6�oM���|w4���|�5Z�o�D������Bi��	�{�i_�& ka�'V��ҽ#�wz	�lZ��GDW��d�7R���{@�]��rjO>=wM�`�����]Ȫ:ga��]�j3�c��uC��p���!�� >�K}Xk�R�������E�ø���x�h����`��f���PcTS:g�$�z����o[��K���4�&R�Ɨ�{�`�� >�Re~5�yo�l"O��*&BΥ6w�g-��qH�<�J��<š��[V_�P�$OH�I�1&��n{ R�rz���~
�?��H�"��^��F�WuS�|�\K����OS�7o���0��	ڎ�#h�����/F��t�8G������^w���>����I��J�Q����> ]J���DM'��W�2���P����p�bu}Ϗ��o�J
��4=l �¸Sa~���;p��/�IE�]Ej���b-��;�Z�bI���9�.�oz2Ui
��.c<Lo���Ck�Q�ex����k�(t�jZVZd�	�f�턆6(���Ο*�z������$��"r��b�T��.���h�����4���W�Uk�8_z�0�H�w���5����F#��EƩ�>�������-�I��g�.!��nޮ����o�ɖ�T!:\;���S���Ŀ��J[j`�wD�	Q��1m\]S�N�n��EV���;�&���ǌ$78�bu��I �8�vF�e�^m���nl	�<�~hrF�UN˻t8ʯI���ğ��8�xF鍴�6�d��,�����5zW��3�yj���V��lr��󓀚L�j�	K�H��7��<	ꈏ��&���FZ�F�Gy��O�;Z�4�z�*�NI|�&�w.m'��;w����UY��^�~��zqo�]��<�Э��M�+�w�����s���[�J��f� G��w�����`��~�P�.�&V�uy�z��Є;�,�&"퐚F��d����Oc��Kb%��A2U����P�hx�W��c|v����E!4������V����A���ղ�~ĭ�p<����n�ծ�Yl�$F��ž�e5|@�6 ��@���|��w�X��}��JbԶ�R�YCH��*]3�V���.+2Qn�)���]�����6Z���؜V*L�l�� �B���K^H�1�\��D��%��"c'3;��|s'�ݩ\�N�ۀr�_��^AՃz��K���V~�2g*�L��*S�HSw.4�J/����և)�p��z ��
#�Z[c�Wn���7b��E�&16c���2E��hY�h�7��´��P+�f�	���ȿ1�1*ӊQ��7{(�I���ƅ�i���W[�4��5a�^"i��"J���R�-3�7����>?&OI�������^DY���!I�w.'ת;�Z�6���}0����_����Y�<�d`�
N�4�	�:���n��6S���=Rz�H�d�tKj�(��O�V4�H�NO{�-�$�j��T�-�g/#��%2��K6?"�hH�A5�9|f�q��$��D@�6��%N�#�Kr��T�`��5�l�D�)j��\VN�S�*���\�)cFx�������z��=����/͡�/Б��+�>�������f^���d�n���;���=ֵM��L��@tij狩��n��7�3v�]����"t��3����%����`[+�~�%ؓAx_�T������nh��H�N;���-�q��ނ-���1���ֈM*��q8G��4���F[)�G���nQ��r�Ci�_��_ɿ�ό��\%Ri6�"O6��FXF��3�P�x��ku�N��������گk���]��n7�ٚB�A��w�k���hć+�Bٌ�W�x�A��+T��-�oU�N4p�	�WM�5X6�5���j���sr�U�:o�7������g2@�J4�!pKZ��~��-��I���3�̃���f������`�^ݚ�ߖ���FA���!n��*v��t����6�>��!��P���,ҝ�rl�@4=R��[+l
����z6��l���; ���Ҽ��H���
!��렱N����\��+�TM:�۵A)+��gC���޹��1/Q*,���0�y�����|j4(��l�G���56���vW;B=s�_�����&l >�W�� 3���|lX�N�<�3������{�҃����w���X�\|G)��)�)�"q����u��CS/�@�� \�WC�L��V�����`Ϝ�m70^�+�V�D) �n#=�OK��o]���M  O�߳`TM�t;�M����®D2��J�<x�Eb!�'�s�ɬ-�wL�hn����1�rOgQ����f?������]�k�|����=��nU6^��� ���.hH���PT�Ԭ�sZ�iC`;�՛�*:D�'},w᠃m<_���b@p��+%�Ku�w[�Ĩϩzm��U ����K0Y^��e��^� ��l�D�ǥ�$�U���͛�H�v���-�H�w WT���Ү%������u�ڴx�gɓr�-2DD@�X�z��.�H�A�J%s)Ԋ��n� ��r2�JG��e���{����i襺� C��{~��M��W �}ȮY���H�j#I��)�oA��+7�1�\�Q,�96���<�1�H߽�6��tsC��Bj��f�hi;W�I�J%���:�k`��`q�ّ����i����)bW�[r�*b�){z���VW�^;��"&��f�fmG�����:�� �z|�5�?�F5���)`G�����)8�y�p^�`�� ��T�nQ���Q�8.9��$נ�Z�OT1�.y��������dB�3�����\���ׄ�q$Eʞ�_��*�`G���f����m����2��kd<Q���hm�Q�BgP� ��y�"��f�>
5�'��V��7Ω��V7��?y"�(����nI(�.��@K)i��ր�w�	���Kok��I��#�`����D���R����^�T$�`lLt�e�=<x�G/f�K_z^�1A���.h=����������KId|}��Iԓ��Z�p�c�v�'i�.��ހ]8OǪ�G�_-�����oEJYn煁��|ӹm��g7a�i���Vƈ�ILEe�xP{�*B&Kx��Z�P�HI�������H��l���y)�J������k\I�Z"�#@������k�e��A�fo�:�3i�<�<����·�����22�~���8�Ќ}�~d��i�싿�F���c^�w�n��H�n��E�A�y/�T�t�
µ;3f6�3��ȴ�����<��Ɇ�KQ�p��ۀ�t�o��% �~� Ԣֆ���xc�w�Ϙ{6�Ԅ~8Z��v�G�Ӵ�bLh���r��%���v'�����+��4
zV����Lb<_�ئ��Y�eg�G����1#�[�uj���C�'b�������� ��D��f����] E,�uj�,E�'!fZ�wK�ک`L⁰YE�;zހ�m]�O$6�k &�&@�<��r?<v]�ļ��qճ�|�g9N����|�c8�9`���K��鄘s ��l�v|���DDAH����ǰw��Inlz� �\�Z�$�=@X��ڈ��u<I ��LU��ܺ��_�7kJM��M�AU��	FL��+e�D�]�����K ���}���I��Ğ:3ˁ���N���q��WM���V6 .�*Uޓi����������a���U���u��C�,3�20�b����.�,�ru͞���TN��SQ�zi����;�I�a���#f�3[�#E@�:�h���%�E@�5�Cj�W��z��v@���nlǜ)D�~�ˤ��u���� "���� ek�wy�%�.
�l�o6�E����Κ60pZ��M����In��{��{B4�D�p� <:S�0@3\6�7Ω>���+ů�ͧ�S�5��8n:��%��2�Kƣ@:Α����	�1Gw�s�qE��D��>Q�d"��Mw'�Tdf�Z�W�yw���g�0��Czg|n��������w$���*��R@�u���q�&v��k;������������G�^.:M���A��������-�#�up>��zj�6"������/?'�-���F|��
r�[Ȍ��l�uώ�qlU!oV���]d_�}|1X����L�^�n���d�*A��[���Dx4e�NAA%��CBk�~�0�������a��(񄴊y�WRْ�koA����uPߵ=�� 6)�&ϝ��Tn�4:j���:�(85Ma�A�e�������zZ/����mL����KR�/�'��7�+#����0Q$G���q��
��d�{-�Qy�ZƇ|3�����2[w���گ�S�^#k���ɊLp$�~�?n���v��s~t�%Q}�EvR�Ck�\Z�14}G#u\�}�.Ȥ�ҳ����q80�|�e}DIXG�׿E��.fb_?�{�N7�g2��hG�C5���N�M�{G^��ӈh���ۆU+Q�-%F�ft\��d��ئ8�Z��0,>�z�TTY�"da�Z�"ߜ�%�
^F�~�P�j^ v���5+�{��!CXpOD�bݳ�Kl�I{�f��-����6�b�][��V�u�l)!��:�#��XI��'�Y���vA�K5���iϱB���;c!�1�]����5�r �T�n��`2w#}��)p�����~��i�Q���~cy�y=��.�G�GU�/���
S�Mo@�ӏ���)�����<@`}tC�{H#�;��^G�iS��~G��-w%S�F]�A=o`�>Cι�$XB'IU��dtVٵ����$�>f�`�PPo���D�Ĭ�� h�h#'ǐ��lȗ�l0���<��թ�󓂅b���W�����(E���UפSFHJ�}��!P�Z��<�J��J]���c΅y�%����Ыj�
�	��6ؒi���aKN�Q�,�0s���>4��"@ �2���ca���U��	���n(u+
OE�n!*l���b��}s��,nrA|9���8�/1��p�·-�>z� '���IM�\�̖ �>f~��u��1jC^s߈Sj���vօ�D]�K�&���/h7���b]���Z��T������l�����$��%qJ"m_D%�� hּ����{7yaz�ߥO/�å��я_��%�&zu������(����C�LB('�2���by���� $g�m�h(���B�=���֋�|P�֪ES�����U�u���+����gک� ]p�Y�;�}(�m�<@��S(w~�gU�0޿iO�c������kt�a�����|�sЌi)��U���ǐ�J�����#o<lX&����iz|�.���d,{(����9���bސ~ҋb�+�h���_�mʍ7�9�R�p�|<���MB%o�|[t��C����<s9C/�_���'�C>r��W?M5�D��őX>F:j�f��[`�}���0
��J�,s��^���u�@�{ؑ�����B�ĕ��FW�R5�+g�"��K����{'?����27�@��N t��N�KN�K���Dd���[�?n�m�+2�<�O%�Qc\����:��1��0�� ٢f<�@����t��jE�u��Oq)�F�dឳҹ�c;8Q���X�^�Y�7�$�.Yn�~B0P�PF̍��6�s.��x$B� @_�o|S���Pe�J3}o��C��"�~����O����&��|���8�eNv�C�G�W����#�i��I�얦��B���� ��Dl�<7G�����e����ڶ�܅�����	2)�!R�/�|�Ӷ��C2����h��w6b���9 S`� d� ڠ�K���s��c-��o�⿽Z���ȃ;�%���Y�\���6�w�H�D�ހ�����yA�Rfd�$�Z���@v�4�T��.�̆w�iPM��&[�Vے�Śl���Ԧ� ���\�s!����4�=���	7gDq�p�z���_�լ��.�胱�=z&�N�'�y��2�/lv�̆)]�ڐ��9rFIHv�R��^�7�w�%��"����j��4Szs�;��p�L~��t�C�������.c�+�]{����޲UJ�g�����7�v81>��:��y�ʓt�����8�������78�S��*
��� ���|q)��U��L�_��j뉸�j��Y�>"-��i�g��Q��/�%�hU��7|��(�
��*�n��-/�}Į'�	���y*�T�xa�=[�V��g~���ъu��Ո��Oh��r+�d�3{^�!�!caM{����
��Z�̚O�-�?�����z�c��/�h�<���Z�k�[ �;%�[���2	'��?�>���z���e�x����B�KAˎ�r�K���=���ǲZ��-֠9@�DT�d��%�(���6�7BșA���W�h�:6h��e�;U�.�_�f�)���	�tQ�?Uͦ��$T+ٶ(��v��m��ݸ��B�e��jܿ�� �}�ݺ��,�a��`�u�?'�*%� j�����8�4��P�.�Hq\����'钲��wU��J!��nb���q�z�(F����KЈkP�d�(h��I�.�q1�Q���z��.��z��U�/�X��`���|�a��:_�?�(�7&�����W�B@sF���T�O�����jK�z�
�O(Z=�������//'��z����`_)e�$.�ЌU~J������q3BQ����[��^�����d�(й�jGn���
5��A��Rd��gc�ڟ�o�X�Qy|�P�1Q�?��9eu���[9>�����7�$|1��?�#Un�'Џ]��|����Z�F� 1Vx��F9��Ξ���vqz��p�G�*��������:�uG���ՁI�XY�����C�J�WWp�O+�$<��F�TI\�{"��.΋��\���T��GO����(3�C
��؀������&��23;_�k��1�M����\/9���2�|H*�m��y��w��C�I%���<|<lg���n61��;q%hjM�+D���N��h՘�t[�>(2�GG���.�7��J�<�S9DD�l÷�f�}�7��:��?݅�%
����o|� ����y��i#A��H��}P����JT�d!r�	lTƞWy�KI�y�Osr��9�3�>�6Tq��r�Up����S�a���j_89m4k�V��(Y��U���Kq�2�G��|�hͨfĜ�z�RdG�c�.(��ӳG�q�T�}<<�%�JY*}���z����!���s~n�:<�ˈ��Q�eiWMt2�J��}%v"����6��1���/)�Y6�mD��Lr�)�f|��rKDf�:"��,���s{~�G�B0�T����=:ӥ��
�gx7ng6�7���I��#�w�#��'R�q���5� �ӞW�U�o�WE��t�SpE�!� Ԟ�I<
S��RZ��}!�����.k5��-����EU*/��d��҇yƇUg���Kk��i,t�/Ux�/�ίg%9h�܂RN8ٕ��5�E�	W�^u�.�y��dm�K{�5��WS{��ˤ(����Ŋ寀Cd����]̡ ����wᧂ�L�n�E��Z��a�<��C�s1����8���j|��q��ՠ�z��5�5씨�!�v�!�#\�wv��D����p��N�f�:4���P�s�*�B����y� �7й�����BX��)]���@�оRF�`��?a��(�������]B�_�î?�$������/dA�fc��fr�"'__�.�UT:�u��$
-�$^&-��	s0s��%���K/�����T�RM*���Dnh�e펌�U���n���0�ܗ��?W�/����ϫ��8�д��iU_ �G]�nVb6�E�(�����m�D��.�i�IM(\��	h����z�Ie��(�ӝaY�+b��R�4W��^D���	�����[�,�f���,�U�X���1������2v��Z=~�`�lq�C�ja�\��Oi�w������g�Dlsb'C^�]M��G�q;��%�C 댊�{y*�2b��W,V(g�<y���q��H�'��*ȁ�HI��<(��b>}��>o�e������o_v��LY̻�`O��qכٶ�����u��x���0�L�;z�?}�!���N�u�9����Z�G �/;d�PR�4jo	���i���$�*:{�:U(�8���ή�dyͽ{���������Ⱦ W�ha����r���V$��dL��Q~���=t�~�T�5P�S� /�v�v�˕�lK�ü%�d[�
E�g�W.����'�TZ��ľױ���������܍�x��i鏺eR�;�g&����]�8B#����j��R���yE������|n�=SO��Ms$߅K#��l�5Df��Y�x/Y�z1h��b��$�$��+���dɯl�٬{���'7_�mm[)�>�?���p�05����y5��ӿ�u�V����W������r3�1ʃ�F�k��w��Z:\�#�C�y2�|�����Q"+���{����/����b}3�e^�vu׵'��n	�X&]<82�����iNΔ�g��h*��#��&ٔ�VT�+�I�T���]�P�e�k�w�q戕ëD���,�t����-��X�cU���R�n��10幓R�Tn�K�'���}U!PND�q���{�Y��}	FHO����c+��K|�&|���۸$�?a��;S8 �����)XP�
$[n�^�}y����V�Ef{k�D���uڸ}XBJc��]X�90(�s� (�K\��?��+�K�޳�)��[3���شj%N�@��?6$&���:o�V}�6ұ��b!�6A&lL���)��l�����y�哘nJ�T+$~<5�ٙ����0���r�s����$yl��ʽ5��)��dA�T4f���`ㄊ���(d���ڷ���#���%�
?A�@��c�J�B��/�)vIl�Pl�cjV�;nv㾉�|��c0�ȇ�(D��#ռFv.0.�l��1Fm�z	Bf�6��e����Yd�}�ߜ}O�b�����j�1���9�A.=�'P�]��/Ş�E�<D���T��������M�9Y׆z/�����tC�+�*FC��F��D��������L��j����"���p��f����R��ebF�k�a��&ThP�]�$��ٵ$DѾ�	���&�)j.=���xt��f���4z�I+��aRr�炙�&�ϛ�����]�^a��-��矑|3�[�s�DH���"��[���[�e9����l�}��v�N�+%�hG��>�r���6"mI�i���;I��7���Ć:�wT�m�m�b�3Һ�^���6՝9*i?;Y��|�l�ȟ��/5�O���ꆒU��ɹ=�вI��Ĵ9�J]&�/鍁�h����ɱ?�z�����!�ѥ���[�ԍ$�	����o�z�es;%�ڗ�c���q��=~��,[/�微���?s؂�8�A�j����yM~N8�����0,���M�����(]�gց����l�3��5���~��䰦Ѝ�U��!�=4[af$.s>��\a����S��P���?�^�R��S3�A���d�]mz���9f�h�`s�~��F%��!�{u(�1J���UI�;�9�u˭�wI�6�?��e�LP�)`��2˩�t�Ém;���h�&$�����DK���7��C���@E�v�6���[��q��EF��=^Z�[e�?�o����R��}]X�=�%�iD�ᬒX8j��9Q��� 9:���X�񺼾��Y��&��P�3D%���,��*��S�K��R%�T:b�]\�p^����O1m��| O	����Z��aK6|u�.�����ő<��XB�i��m�;�����|4~?:6�sS�O����s��큧Q0[��~�qO�k���	9XŮ��d�цG� ���(���|>)(S�`���B^O�wQ��PGTVԕch��P�qH��1�~��hԷ�����H]�J��\��CG~�':0ß�V�_.}�fgxėݤr�f��'���U�ߓ*��~�EVb7��f/��4�uC��^Z	����C,?��&�b�����K�k;������w;?�X-7f�4v�,��� ��;��R:
6���z�K����@\������|֍Z2yv�6ΙT�qц)P�o2H�{!C���1a,9�I�:cnrq���/����i���|��F�����y�����%q&�L��~��-w����5瘿)U�"��5|�ڳ��UJ���a8�S��uU�(���s�5ݸW�����l��,��.d`��n��8@1��aw�[�e��qj�iBˣ��d4�ތ�l�3�G��0��,͠tҵ'�r�=�����}R������*���Bx;9�Ҭǰ�ݦ����n��P����E��ki���taTf����F��u���;W��'�8�s�BIk��Te�cE�Ł��¢rJ&/v��eyr�=���#su �J�~�h�r=���;�tz���懯�p����@SP��F�}��>����~���>by/���}$4\2�70:��WQ�k�G���@��s tm��_�\�;�4�y�LK-�*	F��� ��Sw�1p��p��#��(a�.���o����1�-�ݛ~��~�n2��H���FR��b�6��V�>/����r�.��z��qR��3�u�x��r�8Н�����+Z�X�7X\Z�$x�.��>٪ۅ�~a�_��_ �xMO�]�;.ڪϤ��y��M�ڗֆt��})p�}�$e)�
n�J�O��XW��
!GH����,�|LЅM�_�3$x;�Qk�^]�������3� ��g�.���@h����H[ݞ%M. Id{1�B�g���:�W��k�{X'$�����V���fJ��(.���j�p�����b���CǫgK��U����#�e�i�z����Z*����,��>A��;U�|z�����׫*�ŵٝ���+3N�)v�3$D��'G3���	��h/��6.\w��I��*]�X�z$8������|���f�qI��}e�p_�N�����ѝW ��(>M��:�ޒ����
P���l���= HH	�(���ɉ
�h_��3�N�y�?���E�苾�+e6��jd��hm���u�"T
kN�k���lxǿU޾�s�J㋺�:�;�q��UT�����s�>��eS�NHɤ��щ�N։���D�[5~��d��é��-�~��IB�r)�8�?� Ն�n�p�������Đ��� X��{����6�3��{�H�I�-�׫/�އn�˺rh�X3�R6����e��_HӲ�BPg2 �[�`%т����^g�P)�v�7@�D�귇ZQMZ��c0�:�����ڣ50?ޏ���'L�H�0J���3܁ܼ��k適����7+�=������$V��h��x�6}(�ZO��Rം
�C�Ā�r�rI�ı��y��և:0�E�i��
�����)̊�����OKR�ּ���|��k�_P�Ȗ��p@�"��:�_�<��I���-�}�kL�9.�N���P$._cߋ$�����y��g�ה��<����Y�S��c���y���7�$�v��8՜�RV�k����M�U#�R�*����cߚn��
��,)H�dir�І3_})
&8�/B�]�v��m��V��9���)mG&��f֤���У����F�A�K�C�D	ߨF��LL��K{���{B���h.#u���o:P���c�r�t��'���R�d2��Ab�Mt1����;��Y&�3>}֭�����4�����8]C���^Ǭ��bf �&I����8�0
�����̌���D;��$�̢�h\c띝�:ߞ&��
$���Jq�/�P}@�Q:��+�6�t��P�_�r�xO��1:�}�#��]*�]W�F�Qw-I�e'�Y9v��/��9�!�SjW���!�'�9*F���_�֑�����s�>��1�~�7�AO�3�^��Br+x��%,���s�,ի�6�r�j8���T��gU�+$l΃��0�%[Is�CR�Z����r���KhY�?e�0n� �"Ff@Jf����K�M���W����Wz�H��T�O�s�P���6?T����#�vM���Ǒ54���\U'Aľ�v����M�Ao��E��{6��y�[�,;���`Պ�������[�f�׿-�C�pS_��t�*��&�3�e�{�1��7�0���͇��R�其+�s�k�
6���Lz!�iE��[��l�ڶg���j��+��\jP�#-��E`��Q�N*���Pm��
S~�Fx����d͜�v��)N�qy� �k�-����&�v4����:���br�A���^'!�~x@�	4���<[si�U��Y|Wa���P,6�`�	9t`ʱ�{���t	���_�Y��
^N���P�Hň5g��]~#��2�eїD5Ff	;�Q���	��/��%����F���R��V�-�Q-�$3�xlb%$��2>h�Ki�6_�<X�Јc��n$�PW��I���E@����nᓳ����)I���p�6�z�S�ӯl�X|�`V�M�(F�2�x#n�e�]�����f	e��~t�G�ȶ�����T����`3�؝�r�dH���?4�>3bVm/z�d��xO[�g�@ԙ�S_�_@n������������Q��m�=M��N��\�JmfϷ.�&�a#Cӗ�� ��`���z�u���t,1�mq5��3��ǻ;����]B�@�S�ذ��V��B��}��%rNI�P��?��5/�
a�f��%+���VµfD�o�^[�� ie�D��yu��*%���4x2�P���Q.��h����+Mk�Ǝ��b�$w͠୽}ǋJZ�͜�{j�}]� ����x�*=��K����[�`�/t�ܯw��"#m�#{p|�c����?�ܨ�4�!hr&��eL�t�
�	H�I] ��ڕ���C'�ב��ޘ���S���HI�p[�Y�����JA��Eɮ[�����'i�GvzzA�AS�5�\e�J�~n��0�| ^��T5�4���_�1 U`�,������N�K���.�7v�J+��h�3�#r������D�4��I<\�0����������/�tc󫳘�y��a�H����ZЛzw�����c��Ꝫsl^2��ѷQL�� �����*Ǡ�΁��m$�Z�cc�P��������X*+!��'�{���0^�Z!Oc��ط� ���1��6�2=��J�\}���0�.\�~�G�ui�If2�!{'�t�zm�� /�d6��U�G�l�4"�\��T7��Ӕj{��J��ϗz+����>ݛ�IFld�s��/\�����)<o7�
��DHǞ���k��7iP�+�5�e��^���������Mxv�+�(X�$���:�@�XǫIMN?<`	��+	z:�N�)��S#��>��\��>��O��<`\'�;�bYT�������V�\�l����~KP���ѥ���sb���˦O�r�WIÖY�$��Q#�?��t��:���E��ǀoRL��v��Su"�K�R�S��x*�>ڶ���(�	 ���ɽzWy��y0�2�������h��o|�.�d���	�@r�F���x�r�OTR����+K��[ˏ�[�yH��!%��ؖC	�d��/�F�P@<$�����Wi^k�Up�� e���=f�f�t�]:�F��FB{�7���Z�2���"v�k��cMc�C�E�0'@T���S����k�T+��g�J����o��OҲO���Y���dC],���+b����w�@��o!w"�H����+�n6��=#�y5��ι>$}��3��)�'s4��@�<�2@�qRS�������E���|M���Sl�X��!ub
�I&��0�Nt.�F�n$��E=c�{M�������)�ԃ�?
�D�5$ozed%ESWn�Gw� �aj������q��	j{Ġ����H��o�3-�]�6)́j9��f/-^t}�����<G��a���'��d8��������/��.i��Z~%��*�����0[z����a5���`m;1��li��Xn�΃���5�O/��{���. �_�u���Gʱ����H��á�������d�a����0W�*�(����F���%��eO�I��5_b`�'��,X o�o��h�h}���f<���`�޹�!��cj7���!5T�H��jU |Ozv�����UU�+���!!|x��6O��s��C�N�}����'0i�^��Q�)oj�=�-��}��cMG�v�+;��Y��I�!\g��/�I�g?�%�J3��gь �97���*2�ޜ��)�lP���Siʹ�\;.�����?Y����Q����qD���p�3�������;F6ZW��g�4���Eԗ��>�Aª��2���W�M���&�7;�:EM��/�5M�����a�4����rn�,�l���`)h�j����
��[�"O��<
t�i��e1q2�-���dP����k��!ݦ����ܥ�u�Cw~�����>�ַT�Lq+%�l�5���G2f��IC�E��]S/qR$Yfw+gxר+�ʐX�  [�jq�^F���s��PdƼ��!y0Q��zd7����K��ԡ�-=�m<��^[��)!�c�m3�ZxS���k��|��ϋ���uQ��`SNuEFWK�,&䍭T�>%���z�����k�Az3���O�I�.�ٓ������^,b�x¨��>��׭�4)�����L�cȸ��
1@_ D���_��4:$�{�M������}��&]�k�۔s������Тi���־"n��}9[�_@f�.�*�Џv�
��1��ɉ�e��7�c{L�;9������F8JuV�w�KS3��6� v�$yAT#F�_��rm<< h���
�	5m���-S���é(!JY,v�)B}�/2>���{7r�a^�����C~�W2�~���-.Y�]��K��>g���#ws��0�a�IM����iO��:���)jò<]yּ�Ċ|yX0V�ls!l���~?}�2 �KC���9P�Z�K2_P�r�ʲ}�+I�����A#�+�ng;���4�;��)���!���F�6��%RX��tL�L\��/g*�*�{[7��~�~pD�B����Sva��x?|�<iXH�l�Z�b9N+��ԯ�jq��K��*8h��C����ۓ-&R�b{e�'ď;�u_,�!��%��+ި�7u%L����㋄��o�c�_�B�  ����%4T�*QV^�D��l��-�Wև���.�t=����!�ǉ��*�p�۵�UиL��'�.$�[\����y�W5%9)�4����La�����uƐŘ�5b1�����O��Vvd�F�)�=0���0~;�vA.��z�yw��z3T��Ȃ���:��&o�]�*�bX�*�?�u�誊��b�7Y"���U	s���b
^d5��/(F}�0��,� �x�[[6���A��Do�1w[+7�k�����a��	�����6G.'7������m�v�D�^�֋���,����9>���F�[��v�>H伫���zF{��~�F��fQ+���&e[�MPZ�j�	��>مO��� �D<�9y*�u�Wk�̑����ϮMKϐd,�[R/�d�Ɇ��R����my�����f��=��o�����ᛙ�� �x���' ���YzF�
�-��Zԇ���VB��l&Gd:�jt��Xo!u���H[��J��?C�A��h��Z^�$cT>�P�+%=�_����=W���w�
(���F\�m y�gN$�>INy�;��M'=�����i���j����P���JQZ���ʰ9A%�ȓ��"`�I��'��fg+�kr����y�'_��B���)��-Ц�)�L�� ���t^g��E�ҒL=��YU����S4����,[����;���nэ����!��h��u�LLxc�l�f��T���,�]:��T:y|{�s��娨 2�������B�������X8֭2D�Qx'Π\ N��ǜx(7�W,d/� �<peFM&���2#0OJ[���bڈ]�]<2г-�:�q'	���Q�uYn���w j�j�~�c��������dY"6��E��H�̂i�l�v>��ٖٹC#�K���9��%ډ�{��sj�_�h�vd�pq�-�<#�ԁRX_�Y�1�RR��޳3��Tu	��Th�E��ƚ.Sf_\U�Z�c���6�x�(?�,�a6�����P|�u����ޜ�����#�����Lj�k�,����_�מ&�-S��%��*{�F��)A�'�'�d���m��շE��,�s<��n;��&@|ᗲ���S����ؗe�۝1��G�$�e���j>%�ç����S��O1�')C��^��V�o�t[x5���/��` �<)��QV?	���oe�u�������aR�քD~�h�X����_l�?�"Lj?���#�`�g�M�C�9��۫��T77��~�#;��&Q+�6��f[�w��r�s��� ���7i���5������ �{0z�h�|	�D�q^���4?�z_��6��R���
�d�ء����WI_��y�h�tnhC,�aH ��~�:q{) �)6�I�~|k��7�=��L�6A��ď[�G�1OT���ɉǲ�z���	Ԯ���W����r?�Ӧ����Y�V%6����BA�LE:����,EwmE���[?x���O�S�]]0�0�
���+�����|��࡭�#!�
�[a~�$�A^s(r>m���ͪtm�(�JO��ȝ�`�2��|���O����1���-9�m�j�ڕ�a�\��� ��q��<����gmn���D�:��%�����o��)h4L�B��E�a������䋰����g���G���q�xI�w;�y晀�_�[K�&�-��]��Ȣ�	i�c��EQ-!k~��]k�˸#�U%�����e����)cR�wSu�^��%]6�zc���=� 3�gF�|%��
M���[�c�Ѣ-+��h�Wf�	��S`7��	�gxF��sP�j�b���I8�qچ��܌�Ο���3��A˰���Ĕ��r��B�2�b~n�i��ųn��B2zp�äO�Y���o5B6X�u|o\��IH!��{'�f�����-�����(��W�	|a��[Q$�p�
Skg�QR�DężUND&��@�+�O�uL�ê�2�ԳT˥������F�C�'P񪢥�/�FEvX1RS+��|݊�?_'�`)@�,�E���K�����[�����p���\�1���:NX�Z�������)�Rr֪~n}�[���1�~y�ۃ�;.�[���B���r�S�Ly�ћ�P��#� 9$��5�80wF�"�=��BV�B�<�s�4ARP�~�����d�Y~'΂ށ�u�ᩥ�Ll|֕�M�Bצ�|��R�A-$�J�fPW�bk5��1{�W�C]������\�⏫mmBY�ʬmd��[s�|W�3[0��tp��DM�w'ui�J�>����iK*d��(�����{dd�ϳ,��ݴr��m���� UNx��/}��ij����W�aD����,2��A�)fD��;ݩbؗ��TL�����{jwNE��ͦ��*;���0_T�-���X��w��#<J�
�=���VF �5��\�eV:ӻ���2v�΂��˺�*�[xw�li�k�һi�2>���3�[3AL�~x������[�t��_��*����,�{�"`�%���#!��>c-��\�w��++�'�O�[t�g�qs�˿����H���z�]k�k;gn�V����tK�s�h�ݱ<�u�B˹�l��~5�p�U��
F��Ji�	Cu؍����[��J}������x0�AJ'����(m2���Ua:�@�>����iο����ͻ������ܲ�2 �0��J���wݸ�r�]Bōe�"�s�iDpd��N�@9j(Lk��O��[�LR r�{��zM��4��	`���+T��=>��TV�[��0L����	.��X ��-��g۴����-����w���	\�D�&�qm�r��X*�M��:����s��n��DI�8�^�c�#����Ol�6@�#���P��@�H<���8�V�9�,�����J�2)I�C�4���e��� �i�b^2���|�#���у��hcD|P��:.- |70��D��]����$
�t�닒�ªhԬ!����E?�jٔYg䭬�bZ���P�J@^5\��^s���տwM��$D�T��:��|�WFÏa�ˎO0a^2#+6�`T�,9����f^����eETͻ��N3b����P�2q�v��k��D嚰v��f��x�ێ�c�) ��z/NR�{��Ϫ�������� @���K|�-$��id��iE��_�y�e���!�gI�~�	TH��#~]�b�4t�� �7���Q`��N�ݨ�'a��*��@#��Mts$�h�aX-]T��B*pE"�.�5Ŀ���	Ѕ�Ln�L�?���M�'����5�#�BhݦG����5�m��9E7}�o��Dګ���jlB�
��{� �za�g3K߹��Б�sh�k1a�Zy�ڱk����{�Q;�V�ּ���I#��t���@��1ՑN,��qn$���2�C����o�y�q��D��D�w�!��̬��n(�\��ʝ���u���~��&:��mj0����\�JZ֟7�3ޘ����@�(����:���uL��ɺrJC��Q*!\l�9]IN��2��\49s^6��\��V�N/��|��_�����^����XZ:gQX��khg�`�X��>;��U[!$�@�Ւs#��u1�7�܀��m^Kլ��iZ����lf���o�[9���ڪ��bo�f�u�HxŜ��і���m�����XK)��k�ߦ&�(�ad�T��?SV<�Z�`���i���'��h~UQ��yl�u�L�Bi�XD&z+� A65rRi �%㙹�#r���ŧ1�5ˀSM�z@l�d�X��~�?̇n�7������'(Aoy���Ȫ З�?����G��f
suTQ���6�R�;_�e��¨k(]��A�[p�N�ۿ�DCJ�3�����H`�̫�x�Ab��J�2����d�DsQwՏ���^�ٳ�����ў�6ݠv;D�qv�戧 �x3 ���")W�©J�5c��"��B� X�!!��ׅK�`N��/���s
7H<h��<6�����j��D��8ń3mAt�UN��P8��P�ڝ rs���òR�S�Qk�P�C-��f��X�V��^�u��p�;1q>�O���G7e�&v�5tv.��H*
���6��y\�����b���vu��LH�>7��,���\̚�����z���`���ה5�A�
�F�_���U��b�ڈR̕Qh����>�DO�)����9��W��Hח�˙Fؚ���J����B.�f,���3x��3���&pb$Mw���c���(r�a�����o��񰞣��&�V�&��y�و���g�f�|ʊ�~H���0)�eg�dw�m���K{P�5w3�&ޖ{�a�~<�����d�<��H�F�r��g�rm���W�"w���[G�!L����'�[���@��
.�z<��Bf�}�=�I���13~]ƥBu4�jo�_Ƨ���x����*{�����if?��t��(�3��?�i����?�Z��4�����\}�rw��b�1,�&��RL�/�r�L�T��co-
|=��m��͏����V��l��"o�kvݹ*v��F��ۢ?(F�D�%����X߿M�~p��"�֦�����]�"<d[��[ܩ����]�_t_z�u]#\9�Sb���Ar� g��cpk�8zHjr�=����}��L:8N�^e*+�5J�F�(n�4YE��\����p��\}R�o.G�q�5�9B��[�	,�؄�B���%�Z����C9�� 4�����Kf�"wT�=����K�q�.%�0V��IWǡ?��ȜUPXǥaY¦�Ew�mCH�+b��WK�1�����R�#�(�9ɔ��e�5�{ַޟ�<XU��?w�{���V0FP>�b�`w%�:���ҫ�+���?6�o#�l�MKb;��B�YHr6B���V͜���gj��m�[Y.i�c�!����j�Y���
29ёiq��Q���u$�y���.�-D�r�<q�g�/IC6x̺F��#�%|
�W�d��:p-�r��0���,�3�-u�i��o! ������O��a�9
G���6�������gw�冀��r>J	�V�;��DQ���VeGnO���J�ƃh�m���u�^$���\��%�)!�N=��hxy�y�Y���G�-��iTR0T�O��X�9��N��$�wޟ��䬥*7sBe�T��D7�����)�6�f��3G��qY`���P��*�"��%=�,��i�2��5	H]�B����0n�n�y�3�'|9"���]�����7*�F�%a�X�л �
�E��m�+�vk��+�3�Ҹy�ß����N�/��[��kC��=�zhv��i���~No>��l ���1~-�2�M$ ��.W��!tg�t7���/���,�_��|D5W�na���{�&Թ`�mI>ˋ"�����b�(����IXVx��g���愑�λ���%+���r�,��'��y�&�?�h���_f*� R8�p��-� h_�_�&�B[��N��I��Ŭ2�0��1�*�Qm�38}u]`�$�VHE�2�#?����Z�.�R�p'�Q;���~�:�?��̼����l���덌UI��s�?t�<���À�-�8$�%8E���+��� �[��W�=�VW��� �o"3�̈�צ�\����̞P�ۃ/�U��Y�<�\�)^��{"y-]Ҋ
��������"� n� �)Q�Wx�1�u���Ś>ex�w#{���8��C���`�6��Y�>�I����S �
,E�`�V�� �X�ٜo$[�	�x��4ci	,�JXIY(ʍ�Csv�N):N�t����y���vJ�&�xU�uM�m�t�c˒��������jF@ GT��1Q���Zb#��Fݭ��N������$�mT���?h�o��Ev����w=Z���rA�I�P{x�����-��ui��l�{���G�x��!��ҨF�8�?�*4���;�P�����*�>��"����Ҽs��� c���$/Z�aĴU�|wM~�2*N~n�a!�*�CB`��)�C�:�tzj����U8+܇�����������$�(91(�����2�1(4X�Nؠ��泊�5KjX��}Hl���9ڈ�o��!};��6�ʄ�J�jD��`��49�"R5|c��e���� C�`/fz�V�PÇ?�Fnb�ޒ\��6\����y�!tI�������};��h8C��#�
jJ�f��mq3�}uU��oR��0��B�.Cb1ζ& d#��}�C�9��(�EUP�YM9� �kV��R�ޠ��?�@�(��jŝ�n�D�լ}A)�M�8$s� q(D
�z�-��u���{�u�i~\(���n�o�����ڞ��5J3�|���cSk�[�����x�/�2͙�d���3o�=��*�a�o7���U���+�O+yRƿM¨�@R5P:%Зh����E{ly�*&�5�|�{v'�ޏ���D�S�4D��G/G�.��A {�(����%�y�j=s��_��Gi�$ƟN.�P�+���3*�.�yHJ�
��.��I�4�s}�S߃�ɖ�-���BZ��Q����p�"�U�~��G��@��RT�g�zڪ҄t�3v�+�"ك��[�>�%i ��Z����V!F�o��A�Y��,&��Ya�H���hLȥ7腭~«.;Yխ���5Bb��\k>��D���x��*g����E�C��Cx�B�]d�ɟ�h�ލ�⯬�g
�Ol�vSn	ʲ�����s'N������G�0H�{]�Cy�M�9�J���
��e���.܂������Q��6�>>�Ci=2S�����\�l�U� !@i�����ܴ�"�ٻ(�~��C�E�:���H�\P_%�4ֵ�Kzz/�����U6v�9�辫���C^PdF��P�Z��/�RA�)%su���r�@*�����nn�+	H:��./i� �K��L��M;wC��[�nKxj��Dh-��M('�>#�i����EE���H�� <�F�B����;6����j��^�N�LO�����OP���ꆴ���"��N�Ӿy�Xq+Jj�4]�-��N����{!��;��9�hH0I�l֫o����\���0��@t ���a�\�#Q3��֚{!��~��������a|r��R�6ٻ�����������\��ɰ
���漢��!@Xe�ّ�w���3�����W�}����C�����U~e�T6����lK����ה��V�6G؟�\�Pg�J#Ao[��U���H2Y�;�>�jK �x@0�U�Wj�$g�^�ð�� pd�sߒB1�a������B��a��WQ4��Ř[r%�:)��5��hq�bQ44��z,��%8H�E)Q.��Ժ����;���l^ӑcBt3d �[z]��J�$����������k.D�ڱ!�7��b��P�3t��-�([��1�P�����@��a1���IT�}�=9���,�:���6St\��,)�4�̤FY~��Y���B������Y�����W5�� �r�����d�u���W��M�\~���.��7z	ʹ�Eҗ�9/��N��@�Ft)�D�Wi^�4�����{Ådv@�_�RNNw���˶d�nS��k :��X=*�rU��z/�s'3ɘV�R�Y���U�߹3St~��a5ZH��qn�4�H����0�wB}煪/�O�!�YG�x}��x����~��`z�I.4�O��W���������5��S��3��r393�;� ��+���d+M+�!{����i��e�1�<��)fa1K����B���|��("�q0�nÍ叹b:/+G��f��O�>3�J}E [��h���rO�y�g�o��f/��.0�׶b�C�w�u6r�Z_s�v�����t�`~��#,�D��4�"��v��?��f_��`L�� ��D	��%vRbn8��i��Hbx�3c��B�D�����(]8�Xn�u4���O�ߟU*����J=�;���0�k�K����ϭ�J?��U3	��bA�Uڿ�5�����Y�x��#tS���$U��N���&̈́F�2q�r�tڶv�A9�'�Zv�����0(�.��gk�w�d ��&S�[�S\�P<1�+	��lr�X�7|�B���~I�K=��������u���o���X�
��ـ��6�Υbt?�fI�\��@=�P2�o��񀖁����鸅���Φ!N��T���JBX���m[�[S�������e�]gݘ3�ħa�bݵ�=�)�%����`�Nj�ȋ�����{5��!�C�����l}_ӤeP�&�\�Y��Nv�^z�`LX�Y����i@�N�@=�U���X�=�v�E�7/�g�1��?�soɏk�Z�7���?y ,b���{�]|IQh7��k����{�":���T,�]Ο�bM�H���y=�\�"���-�R%�VJ�����JN���3�a�%?�)K�XK��}X�����Wx~M��S�s�нƉ��u)xŖ�1�s�3��w?�v�C%��̶�{�&c�>�V�M�@Bɹ?�`���%9�L_(0���Z���������X�I��v���V@����m�-�&�@2���B�(��_�����
��'���A�tf���pR��G���,�9[�m[{\��]��Xh��<���Q�<l��@AAB������͖���ݑHD�3�>�z����۝��gw�D�=��SK0�G�Yw$߀
G��C�4����Iϖ^�^�Fz��oO3�UѤk4�)��XZ ���`��d�q!��%k*k��*�r�t��zz��i�H��R	VN˪Qf�4n�/8m	ђR;��"C��	�W�E����3��Ϫ��j\DǷ��&��{��x����d�?�ȵVP��/�����ɹ�Y$��I�4��b�N�X�FU����):�;�iI�l�/c?b��ؽ�z���e��1��;��]�,D�2|�8/��@�.��Q�>�l�9"��*��"+ �����=i8���[$��t%�)N�.{Ꭵe���:�����&�P�̺V۠gJ#~��[ў�0+>n�Z�K��G��V>��Q4�x�+�J�YR�]��˟GxF�-w�e��(�Z���=�ΗO{���.̲HB/�2P#�^�GͿM��2^\���F��~��L(�29��cS./C���	%��%�P�ol�
8�-���:��$q���8��F ����X��V*_����>����d�n���:!ҌE�;��νf�+�0%~�1��^����@'�n�5����C��x�C�"\ۥ1��/�� ��"|ǩ*H$��Ο�������a���!�J�.�yv�K����N|w�9�P(�^�M�N�ʲyK�]QZ�6�>N��4%o����X*K�ϔ�������&5��K�A��+c7
x�t����Pt�LTZ&
BG8f��!ݗ��]���|�9�gM����@)?L�x�S���z�]mӟP~��%���&/40�
-Y��`%��8�[}[6Ð��s��V�S&�1�-:�GItm��a��&�`4�mG�P��]d����:����jV�zy #7�޼<%�ə��q�-��q^E=/g���_��������DqaR�`w:�V�CKM�~�sr�Ƨ��q3��(�Q��SʗS��m�*l�M? Ǒ
�#s�/$���M1 ����5k.A�~���JQ.�4�K-w}��S0���#�F�a�{;�ѽF��gkKM@&�5���d���]�{rh#�F����@�Y1���-�Е���6/	��T��(y�ЫǞC�ϧ�&k�3M{��$p��KN%a�Yt��:���!�):����罽Iﭵ��k2�P����?���T�li���{0��ŝ7���*?���Ҕ|m՟�u�چYv���0t�4�"r(����|��Ya9�c	�rF����~��Kyׇ)���	���n���e�^���밧��\t���"t�����+!x��
X|4Mj�x(��"�2���2 ���8u<���=c=������w�:�۞OW��0O�
1��iC�IgM>�N6^��YC�<�K^	=�Y���S�l+����5���%�M�h�#��m�/5�T�H1u���)�N�=�l۔��,��a��?�5���awh�A��[&�
�]�9�|W���3�� �oH���y�]��Eǅ��@+�b�'P�R̥��݄����Ӽy�UE0;��j$���ӑ�ҋ���I����������&������~���=�P�^��!�=�K���t�Ek��
P���
&4VD�^E�At7hO�S�=���GY\kA(�Q�V��e�h�}��O:�}���J�@���KX���L=�$�G���Y�m4i��n��|8�Sz��@�SR;Z��i�u�10e���>��aQ��3�1�q�2�Axg��|��?t耺�^����^K~�U�&]����z���
5�\Y|�=*!���㾺���J;=�GǸ?V�P��=�40-��E8K|c2���%�bj�a'���L���LdI�Q�W�5��#~B[Q:���8
i��󇼃��_��u�3mǭn�O��'���>�~2��Q�X媿M�kr0w��F�WS��ʽ���B��
�2��~vF���<-.t;>+��{���7(�`�my�b�
CB�m��яhU3�̲P2����[T�y���Xi��dZ�� �m��v�
�t���`w[�b���)�g �DZL���t�i����yKs���	� O�
�nOO�c���Ô�nk.D���5�+�}��`��5B�V��d	��nq}��|�M
��H�v���GM
���LOX��,$�K)h�
=�l�ߦ�t4ΰ"�Flr-	�%?����|��5J�9���c���&#:c�$�B�Nܣ�����1;�l(�l:�������8�O�7h���J�O�������fF�����z=�%�PN.�M�G�AtV"ҽ�T�5?���63a��Z#ǚ�+&,�-I ��3�H�zO����9��X����G.�OS-�NǄ��f��IwCũ@,�o���9�[��gg@��hM���t�_�B!�|�8�,O��{'�7A��nJP�J��]�7N|���|M$�]5�*1*������bõ��-o9~��ⓏC�${J��Bp8���3��<���vѸ��P��h��H�W�{bݰ�O#�E��!��Ur��B"\�c���QU?���qF��,Δ�K��D�N��/#�ͧ=��w%�U��=ڍ��$�p�V�#�����b�ځO�켤V�Qt��ǆB̵$������ 2<p#	���;)�U�K��:�,Tgw��0k�s��~����5���s[�o[��uľ�Y�37*{lI�]w�����y������j�M�<�N�A�x�<C(t��h�a��lc��Ed3EP�(�U$�EO�a�����AJV߃na�D�����*�{�A?�s`�1n�������&����54���e=�]�:v��Dl <s�D&ކ����H
Z.5H(��&�2���4y ���sw��_o�W��u|.����m��wM��j�:�)
֦��E��w,���t�Z��E��9F�)@�� ױ�v���|��}��L�*�Z�D_vʳ9���eK�y�"�9���/YoX�ñ�e-!�8�+��� ��pp,��!�s��o����)���-�Sc�vg)ݓ-���[lƗ�p{9/(���2��?Nl���5�8�����P&�L	qPۼ�7˂�Y_'<��.�aH$@\�Z�b�@>'�O��ʔ�P��7�� ,���u.��Խ����� q_��
�gU����B/�Рz=����6���(N�̊]����<� ~6m�� ���B-5/Vs@��e����u��ѩ:����bねC��@ܘkB�j��[9�I���_p���aQ�B:9���^�� �"1��%�<Rz��%��ύ��܉�;�W|w�'�k��i0`Q��$�*!�ԁ�,f��8����l�© ;ӷ��8T�u�f�����r[#��5[w��(aO.B <�e��ͩ����1�۬�Ѕ
v��E��3�g.�@0'�U��W�Xv�DN#�<�Ş-�<[� zC1xή�y��`�n��qDK�7P��oW��04~�L�ż?�b
�+9�SK�a�(��сݕ~ڵ_("����$S��(��wi���mtm������3,�hF�)CR�� 5xv:���" �u_sF�S�Z���$��ݬ=��':��_��eNv���NZV�>��D�Uܲ�c!��DГ��kv��>����jL$S.,F�����2=6�jw��}b�$�&Mu,q"�}��yC#k���"��c0��$��Mb鱤X��9�)����<i&<Ut��^�F	�����,_cp���r E���ܿ���T�,*��Ǵ�i�����~0��b��>�\�>��P�蝤82�.���1S���J@���ن�u�d�q���ƞ^��$����nr��8#��v���<�n��2�K���ބ��ɢ�����0��#�0 -4R�KqS�J6�;<�Jb�M�A+b~Z*�H*�5_s�fa6u�M��9)鍒S�b�«Dq�P��*D0o!�\P�Iz�Q�P��1�"����4C$�*\AL%M��K@\�����vсq�r����t`+x�\��^�J=��~2�����\J���� ��,��R//���j�g�3�h5��|���#O���S���x��j�|��m`�^�}�:��]�^�9�퇿��A���B���V%c<;�|J�@���t2��m��Y�u�G�����R�.mYn��:���3�y�����U:o!vG0�Oj>u����B����@�N�6�Ge�2F���=�?�N�J_2�ނM�׆�63.� �7E����n�Kc<��3�@u����D��\�o�ڒ�@Ѿt (����&�<ϒ^��f�Z��n�x�[�k�(��;4{�����%��r�@��\���S�Y1���y��C�i��xUo���2	�k"x���-X$ϲ��+��i�a�S����A.����M���>�R2vؽ�}�۾�hc^TJg�vUze���ަ������È(<,�|/+�G�j��m�F ��x�~��
7)�!ũ�m���|\.����3@�|n}M��m��`������6TY���#�E���W���J���pj���,}*��|
R��I�9T���������9���̥OZ��Kre�����r=�g��A���rƣ��}��S�C��
V�L<�6��s�;�8mJڹO�@J���Ql)~*�C�����y�2�ϱ���j>i�iܩD郧������
�ǂX|f�:{�Nz��>����~�D�$K^zi"�\ R�E���.��	Rl�A�%b�*6����?-��������<��~)Jx,�׵!�	��x���+�>q$�v�bsb��	ph(jh�37/_ѝ��#x���BC�|�j0�0��ǅ�xcq`Y(V��%����j�5�J�}1����MD��B���j[�l>ĠP�����tb���Uv��2�N��EFp�AW� �1M,s�<�@��lZ�>E�up:�@�����o->���&��/��{�3I�>G���g��^#c��v�R��(q�G���Jϳ��W������?���Y+?�����83S�Br��(�$�c�/C����@,���aƁ��j����Lgۗc��"��)ҮA��o�D��ο^��k��2�p�P��ԆR厮dg�,J���J�V[��0yr��0�a��8�1g����y��A8�gU��Y��@�<�Z�(�:@���l�њDC�j"pP���P���a�+���^+���y ��-#날o�#ʧ4%���A�X�.	�`S-%�Kϭˆ�4<엨Vj�ar�X <
���{��8�h^����9ŞhP�L�b��zm�LMc�V��%K!��&�5	#���I�ؖ��,\��N<ܗ2��ܠ������5���o�}�>x+j��7����,2�u�fh�)i��yK�^YY	EF��M	2�[AG���pde���m>݃�*:?^0����M����0��f!�bA*;���nbZ����݋�6L�ѭ�;�ƨ�,j�R� ��R��9(�5%�/�SGm�%��̀�u�&{<R��h?h��k�I�w�<�������)�f�$�qvsI>3+^�+>����G�ƍ���������G�������pw�|��]F?�'AH�%�v�"�RV�_��,�sKyBJ��.�]_���a۴��9�9+������{��/�����%�W�$���l�o�0�R�[����n�� ���#4�s�eO�o�K)n��F@�N�ng�q��χ�b;��)X
`��8,��c��z,�]#� E��������D-�q�#���;��yE���������ZS��/6�U�̹̘�O�܏���۩,��u���%��S>��B}��#��8���������������L��m���k�wk�y����:��0M&kƙ���INg��!��� �Y6� ͊5��m'$�-V�	�H(�l���y�ԟ�:��95���ď��(��\�.i��3\>�qG%d0�>5�6��h�%��\I0��d\����'�c�K��դm�<E�X�'0d��d�%� A:���P�ä��8��%�i�������o'��}rS�o�5˄1�����
/hr������/*�ʍx�L`Q�1!ow٘�r��M�nt.���+�෉����rbn���lk��� О�H�����@x�1�55�{D��Urg ��Q��<�D�~���Q��)�����U
�#�R,MA�	�0�G�>*Ҍ��9
:A˘]�I�Ӎ��0E�5���KM��w_6�Xq��k��'��"ɔF��㗽��Yet�`����q��������#*W�{_�"C*��w����j���d-ǐ�O����@�[T)�c�]�.3��^D�a�� ��B:�*����Ed%J=���Ũ�r���+�Y�S��dI�0ܦ�=��q�;h�a�{�,۶]�'Pi�82ŨĎ�D���$��>�m���5x�m1���cB�)P-�tM�]F��޼^�׌�i�Ͱ��6���N��4
ζ�r .Gh�g�>�ć[��J�ˍ���@܀�yEm*58�d����jU���0�}��0���{���yv֓,��h��{�̇
Hv.h�Q?4������ۤ�������q6�Hy_��7v%� 	w?Su�̩w΂e��ZQ�[����_ W9V�{�9L��A4K��<z�����w�a=�Il����ǆ�'��y���wq|����}�@"�YƮ3#�.���˝x�����RYY�d�e���3���rYui	��@Ak"ٓE`��{�#�
�U�vv�,��p�$C��n��5/�%�S��}k�%6<��� ��@=Y�p)�{���SsR�9*E���Ͳ��c[E�o�{��d Y�����k�N���F���H�7TR������}Ѷ���]��,z����^���zP*9�9�L���e��Hj���P{�T:ժb�"N��г| �(�>���^j��رy��(P'S|G[�IGD��C�5�����E ����OĀ5ՙY9�a���l��JJ X`nx5�a�͇��n&l�@���=%�?��Ȏ�����F�+@��~,�s�'x�q���+�����e>��/VA�˪���z��*����Q�T,8X{s8=�v�6lR��(�Sl��Ҏ�� ]��@fۊ�ڋԷ'�5#ʓ��_h�����R��S4L��H��/��A�G?;������f�C�b&{�c�`�i�6���srgJf�x�=Ru+��,	[�:j�c:� ��KǤxʭ������R�o�BtB��_NQb��<Vf~��L;������(��_��pm� �� T���JP�C��R�S��AF���Ek]O�fl�4���/2�CSخ@x��*n��W��������ii"x�����)]���s"���	�=���9�s������\�zF���P��o�H�BX]S�N�ˉqa@��!�-<Eu�8�s��ȩ& b@g��3�n�vQC�I��{����Ǡv���������Fx&�g��
p:�a#������s����V�wD#�|l�� DF�ٌڹ)��(k�/���R�A��1�N��ND�@�K�CqԚ�$.&3����*�!W�S]�[��~�|���dm�qJ*��0V�84W�Դ�S:�Q�h�2$��!�
�B���c���[ڋ���<�F����a�a\UT
i����y螷�/���� ����c#^%�~Na8����2�#7j��_g�^�Q㓂�݂8�'7@`�a�kN��{D8W�r�T�[s�B��{�������U����}�i�O���{���4��͆bu7��˜Yw��Ӳ>E���C4��i�t-�R�f�=�x+�dԈא��#��ګ����L��h�\��h��y�J����~��]���k�)�t�c����EџW�-5�W�a����юh.΂JY���� ��-��c6���n\�SYm�$yq��j���YݏB�!�,�$z7H��CR��3@M�_�{��Q-��Iaz���w�<�+S�L�="���!,���H���������WsrBcʁ��[z�;��ͨ�e��Z��do41}�lF���DIȞ벓Hn��>�{����T�.a�*���mu A��@�m�zh5kI��8���z����!�����&3>r��<7��g.Z%u���W��t�<+��X�K�'��bb���SpsP�S���(?i�i��/�e|xࣟ�D.�����Y�m���W�֚�i
�~�Q��^��%���$��Rw���t �W����xb��qNΐpTȳ��A�1�������u�
�ڪ|i�`��Eӎ�փ�����Ⱦ�e�`G��P���N/�0�z�
p� �j��o�1��]r��o���8mY�@	ڝ�P��ªK鐀a��0�9���/v��2�g�ǧM���k*��t���''��)wV��86���m��m�NI�建}�[r��3������<(��N@`Tzɩ��u>Ճz�B���&S|��W5n����i�-�t^Z'kD��UrJ���� @�B�X's�N��L��K
J��x�tU���J[U2$ ?��ٝ����!6����M'X�K:�ljP��٥��(	��1YU����.���K�26�����tF�
!�jYR����|Xr�̄-:rq%NE��~���K&4��ql�Jc��M^���5�H!։:�����- ��g�d3��r4ɓ|�G����y����_SC	Y<����ꖤz�65�+��W���C��j��Ͼ�~dU�*( G�\'��
�[$��]��B�3����L�b,*�B̻s.T�ل�A(+uRSG�AoO�rm:G~Z�?�CB��rE�
`�e��}$���pml@���F1�W�����)���-�=���}{�m�>C�=`k�����{�����ƚ�N?�uwP�a���%t���-�-kX�I;�x�����uZ����ݪ+�����9�W���BҢ�H.đ����Y_˩Η�Om��O�a��Qe8��m�UT��1�l���O���S_�x��N]:�<DO������<O�#KqjO��E�����2&iRw'����:�5y.���~p���1�U�L��(��RG
��
�:�2}��0���$̊��|<���l��T��M�^]�0O�PeE���KS���:�E��As��������k��#.L��P�_d�o��*�õ�x"��!:�h�.�rNCZT�Z{�lK�5f�c�D����l�-��U(�������6�҅x���z?X/�4��A��$��)g4��MZ�S��y��2v,�o�{D)����V��B�#����nJ���;��� GK�����{e�t��F;G�D�ɎrD�M&���w�y}���d��k���Ha�4z�)�N��O)W���邐�[�@u��?[�;����6S�ƙ7��e��l�Mm:�3(U�Q��w������r(�d>�8��XcOi[	~���+-��x�m(1�)H����ś8͸��dA�8���5�cP�­br�Õc��5;�B:am�zK���v������<B��-B2��R�j�ti�p�X;u�4i����|�b�t�� s�ٵ���{��!��!����/	];*S�3�͉J�LE�zP���?Ċ,5���E����ߪ?B=z�� =��o���)���4	@�`��S��9���SyI~Q̀�x��� �@:��0����7
/� �A�݊��.��w+�y�՛�:���b�yf)qo�I� Qm�����sy�+�������+�DN
w�v)�w�کUBYq�=�fcfӀ��O�.��^��!�%F�ؾݗg	S�voj�G>[�^c�寔�Ɖ�$��,�, ��zjۗ/���?�i�!�\d!��B.6y�Y����v=����oЍ#�������1o+��|{�k��q�	�D�-j���\g5����5��m�N��+�@���>�a�ָ���9N;X]wZ_�̀
�4i��
����h,����4w�9��|���J��n:=07Ϋ��c�L#ǟ����F��o2S��"0 �o���ڬ�952�1�[����
=�ŵ�W�T.?�6�7P\�xF�\�p�e��IΕ�Ibƿ�D��M�U�Q�iќD�;�W�1��Cބ���ר�r_(��b^�N`��h޸�<=F�&6����}#u�sFj_�����26�6����&Kŕ����e[���0v�L[�篊n���u�a9G�!��e��"6�%6��N��2�u���}<��d�SJ4�BQ�<�T��ب�\����++J���#��Fi������NeN���jf���}�b����-ｅȂ�a	�0>����ϲ?��k�G@R��9���
s-�p�<>ǖ?�_��0�-n23�N���~"�iYSL��U��6)�5@���{�2�%g���,���'���c����G>�aR�۳'%'?�\ۻ��Sb��Ntg|1>h���~���=|��3#��
s��n�D��oۣ$M�`B�r,ҭr@%u��f�ub)}T���eO��b>SH�m<��h*�̹T�S��,�.@�vY��~�/Oi���V��c�G�����n��إ&��ɼ�dw����|5x5�/�J*u�Jی_��O������:"�.��b�yR���ͻgR��P�Wk�1�����L�V��o(^��;a�mU(�q����MG@�S}�=��L���05�U+��Z6����h�W�0�һ����u��X��) H�۹�*p��m���P��1*g$�Z�@@��keAB	�u��;>�[�ǸA�q����=���Qc���
�`���}�$,�Z�<'����:���,I��zJQ�C���L��w�'*Ar�Ó�G9$�Q����acS�u�*Z��p@�-����&�GZ��*�V��z�<=�=���-	<���E���{׿v�"EI��]�1	"���߇�\������PgVvo�ux>�O���T�bl��u�Q(�n��#U#�O�3��I��{�KR�OT&��u�$9���e���� -W��ڕ�1�S�
��v;�5�'F�L�o�ߢ�L�!����pR:�H��<��^��
I�SrY�<����:pYz'�B��6�lG��Jt�[��˹�Yړ�� �7󬂮�a��ť}�
{ڼ�b��8S�$�!��T���O��a��) ��u�kx�`�� ��o���Q7j[eQ7L ��E7���6wy�2nl�g �fo�I��m$2N�qe�:���"�=�β�u'=#E���Eu`�n~}�d�#�0���M�'&�:�SZ��K���؝/}'Ɖs���M�A�v��p9��?�����UJYWSv�9�@�`q=�S¢5 �����(t���W��O�=E�&c�>Xg	2���B��kG������иbh��vѪbSIc�I���o����1�d�"��d�cV��"�$��ZO.����\Ck��^)\��Z	c��zu����#���E��.��sg�>;�`���0�E�9
',��S�)��׌��MS�-��|�%Q�3�A�瑯��7���E���Q�p〵�C67�)��[�iV�#OBb��L}^�73�U'���%BU�b�#��ӆEؘ�\��
/�$�q��ڕ40L*��ɾ1�̗	�Dm!��֔��~ڍ����Ⱦ�,)Y_e�CV���$����-U ����fo2s4�$cKm��xq#�:�����n�G�n��["�$I5���K�8T��T�bAߩ~�>V��X��0Q�
��n����^A>�$DYk0�Ð�Հ{�ؠu����YDǡ=���W]�Q�3��Yj�wQ��)2�nxb_�L_gG�A={�ȑ������9�P�m���_�[+��B�~�Nhe��=�������v;� �7���RZ��:uL�'p���O�l�9QJ3Ã7&%�&o֑H���ș�;}2�i�CMu�� ���)qcÇ
�X	m+���UW)A믖dl7�f�6g�rOb�����0(����YJc��M���{�4��~v?Or6�B���y^�q�I{H�/�9+-<���J���ei��O��K��s������W�+Uw%0W�dU��j|ԋf�9lm�i�^N�>V�c�S�Y�ϋ��`�T.Dq�*i� ��w7�cG�n�3\������ãd�Y �Z�W�T����;Ss+L�3Xw�dsm��%��ٴ��n���?J��:_�d��iGt�D�`o���ֲ���2�R�$� ����?V=��^r.gg��l���dWI�{��֖mmy6� j|$�j�eX�]gUwL光N��靭feuW�EV"��Ġ�
��}���{�^tت3���wNr¦l���}�ئ=��:lvA���%�8q�CB�V�A!����U���E\�,��t�f��Jk�;�j��7�[tG:0��&��̝��o幽UKh�:u!f�w�B&Yy.X��hI���!�����4��֕I���@p�"���%2r�=��.��vR�W/��K�*Ck� �
��EϢYXib�m)�� L:�
�@R���p1:����m��bPU�:v�0��I��	!NrJ�O�^ÄDmOB��Y�w��Rx5HxG?ä4���R�0U���џ�zH}�d�St����A.��\�<-��t����:o��
x�0'��0�QA[Z:�c%�HR��4X�=�5S ������L
�N�9l}w�)������B����]��y����J�Et4&)6m��߫N�C�Ise
t �`�S��������� _���?��>�"��F�#"�y�����fR�o�s��x�;��E�
'��3o��T���Y zx�@�,�-��Xݛ(@aZ�:OC](V-��_=UI�-b8�J���9Hݳ<�f �g�FN"	xr՜���t�Ե�W�q�v�����	�Q�t�ĝ�q	NS�5(#
� �.���F����EA��o�dR܎�=J�v<0hKT�>���+���줘;I�O�dΥ��Q��s�n��Q���g�����K���V#�?�u�	�߉8��_�e-T�H���x�.�WJ Û����W\wS�?䴽�׍w�"�?�O$���4�%�d�?ԲT���D�� F�;�٢_� �&�oN�#\��a���{�m�����?�J�3L���x�N*U��Gi��p�`����߹��d*��r2F�3k�2�?;��q��f��"���W��<�H�XC�7��6��h1������r_"��
�2��7QL�Kk��U��k�D�r�H8��}Jp�yq	
�)YU�,S̼Z	��M@�=p5�+��T� =;6�N�ɴ�Ҩ���b���Ć�&U��w����f�#�׆y��� ��eX�Qbs3{��I�������o�M8A��\�\�Ȕ�R�Q�/�sX�hXĽ�@1�F<�����ܼ��y�Y$g0b�y�P�~�u�~l>����b��tva��u==%)�
F>��{g�(B�m�e�r�s��K93B�w�̱8m�q��m����V�Q�u�bM
�32cn��1~�W{�Bs�7��P7r�p�R��޿��=ϗ��Ћ�����W~RH�LS9�����"�A�1���GCd�5γ���~�ˇ�:��B�(W	���t%r�o�F%a7s�~�U9G�3�\#��J'�N ��smɜ��D�x���p��̀f8sR��4�(��E*���bϵ
Y�VK����>H���n��.(1�"��{tYA&:��X��~ެ�!+�c�,�L����l!�-��=v'0�<GF)��f3��zYr-O����Q5�!%�N�"�B�]��;oē��K���ĉnKR(���x6�n���F���.���®�i�4Y d��G�ͤ�rF�큛;���:���A�X��b�3\���Fy�������>�Yi���Lp�)�;�_�W�9PWC�`/,8�N/G���fuc���H.��(eG���B�����OF�y3he��ǚ$����L�f�QHT�υ��~p�|��k��'8�k,\���4�|�z���4�ԧ���hX�6�ީ�~Un��y?̟�Ae�+�H���Ŧp^K��$:X��0���T��ɱ�ъB�)&�+�>#��1RUhcp�a�r�tu���p���AYRZ�ga�N$�h�.��v^�wv��L_�*�Y"�<��#�E��6�ӲZ��|<��Z~�< Z�EG��TQq���+P��-VQ���%9�@�I��� ��c	n�(`���R ��0�ނȐ�f�-�4j'�6����e����@K�r񆨖����WDy>|�E>�
�b�Q�J+|�~�m�o{������	���Y�(��b;|zP�	w���?�n+H'+W���M1��_��{]E�ϖ����l+��	���0Bv:$P6o^='�@�}qb�GD�{QY"�<�n�jY=�����T�5��{���*���5p J2���Z8SQy?��)Ed�y��lmd,j%�&p7=r��X޽��\���ŀρݪR�i�"R ��s!~�x���
�|cZT5Z��ԁg-$7�}όё�'�?c`h�.�k�Q�.�ٺ�-��׶�L�;+�V:���>�#ߵMt��_I��56��@�}�	�����	ƭ�}]�!�0�A�^e|C6A��_���Z��<rh�n$`����SM�e���/�9~��\��T ��FK5�Kc�(3�^]F�{F��p�X�d=��Pa0�Lo�?�=1v���\Un�FBh��3��Ef��4�saw�v\��|��\��Nqy\`v�����n�v3��;?����}SIu�W 䧷2�Åכ�i�h⛐\ѩ�1SK���F _T��\Rf�j�zC��M�|����}�K�� ���l���8�����2����3:����� ,�Y�p��6O���Fs�1�7�ܡ���cG8�H~+�� m�S�k:���m��k-#���+��uE�-[�AU_\'��h?G�^�OVH�Pk��sY�Z���ʅ�6g�岋X���p����᾵O�z(�#���0�ʂH�q�\���j-�5e���q��&�nEPe�ȁJ���6Ke�D��l�ɰ�¶��8<�������J��Ĺ�-Pv$������b�,�����ƤW.��=?g�����C�O�8]�G���K�U�
��R���=���ŲL�Xj�G��GG���}1u;�vZjMDS�n���.i�V�;���O��u�A��q:q��\����Zss�덓����O
�\����2��/��m��	P:5+�W���kvᾲ�uL�A�"�g���j#�������6���9�ϊ4�]`�I��E�R/.8�!5�9u�Zv(�����|"�+'��"��%���ȷd�f����gf䤝�ݠ��>�"V+�)�}����EJHǾ�Y7Y�iA��-���H�E;z���n�E�}�R���=N���$mu�\~޴#�/�X]�j�7��_�8�n��}0��r�������ì��#[J'�x�'g����|����+�d��*�o�5XH�x_{+x�;]������f3�O=Lk=V�=�&Q~�ݒPR�87�\ 2><z��B�H	�}d�T���+�<}��
����	\U���=��]$��ς�-�d����Y����B���+�|��7����}c�~|ш3nBK���wCGY��`_@�.� dR�]ky�N��L`Q�M]GX�1zdA9
Rt/ ���*�'�����վs���8b�5���4��xI�F~N$}�h��`�|Vz�rnuB�n|]�b�)�\�/�sf_*��別�4�z'�wX�L����X[��HcG�쎏�/~O)n{��<��q��I��2��e��.�'���+�Q~�At�	Ѱ�������C��()��A���
��=c�HKe��R|2ْr0���lrϚ?�!tʕp���[?0P_']��_���L��Ba�1���Gvrj�oK�c|�2aԏ@�U�$E����0�fq�Q������ ���*v���ļ�S����Pw��JW8?4/�����a�ΤnPݠ.E0z�8�Fhm�6�Gg�P�D3���<�6�a��h,�g>���/ �n�xG���o�ѹ׮�iT�Ҏ���ZZz@�\T��Ar��bL���dn��.r�"R���$`�������w���h��Q���A��*h(/@8�����̻���J��#\�Iҷ�.��c���V�!�� �%��&��q'��E޸�V���KW�)I������������֭�o�|�B�M J}�<3��x�� �#���(&@�������JAXMP����" R�m|L�L��JX �b&^m	�
�z�`���X����(n��?�Ւ�dd��`�B��t'a�rt�����!�T˳��I2��45_��@��ka,�j|%�0�)>C�Q�L&[kM�)�yuÕ��������G4��fs�y�/�hv��ף#L��Jv):��Su��>?��j�����Z�k3\A�j�Ç/�)Un.D��;񵞟r�tli(* n'I[�bR|��5�aI'��1'j���z�Y�W�����Uf�qv��������p�����M&(YV\KCG���	wʠ	Q��c���"�*���I4B��^?�`u1O��,M KU�n���,���Zr���3�띾��#2�L�iŷ�6�H�m��K�n]���p�u8+\�*J
�[�#�#� C��ղ�O��CPY�>"yk}��J\M������>����v�h�R�;˫��#�"�F
Ի��Ĉ`z/�i����=�
/�4��/�R�N��M$�����q2�UU�����ҫ���< rL��������hW:������u�~@�<��������'��S��:vL,�n��N4�ાd����-ɓX���E��p�`�o�\o5+Bb� - �:���R�(	����JϠ��ķMu�&�iO2�wh_�4􌦨���\A:�/Q��3��c�^�f�z�WbU=�)X��'�����i��L��"������)��(��T�C�P����v�	���8��Ӟ�e��U`�x�+CtQ�j���<�����FB�
���&M{��Ir��b��=<������C%�	��,�2�wu�u��J������엇sÂܺɅ,�n��Qh��E�Nt�����10�����4��VaX�0�-���'f���$t}�Ȯ~T�淈�����2�]T�����xK���lJ3�VrirI����3���a�mЀ>���`^��;��,�ۆ��RR�C��l�G�c���P�cd)&�� �z4	{��ʐ%=J�K�i�k���k��#�!?#tL5��ኃ>�Q�%&���i�/U�$�h�YU\Ke��1td��IP�8��q�7��8Z�l�y'#�-)��V�������~Y�?�/ԑ�|u_*�h�e/'a�Ӗ��͸�@�am��U���h����G�P�[������LT￳��@>����0��:wD��kA��5��\�95<$�����&d0���5����}�[A5��lF��?��,��n���J�@}!P&�FwW���$'a��~����2�Ӵ���Ld��SCE���"Yu瀇�?_��V�R�����WiD��
����I�����ϐ,���Hª6,�3�C;�O�6�M���U��ڟ�U1�$!e�R����n^E'��頨���n��8��Ƞ��_t|��J�&��;��`c7�f��$L	�]q�t1S�K����r+Z�R�M˴�:�%�U����ШFa��Q0c�!��S��mݲJQ�~��cM@3���1�XV���b�jR��h�F\5�:�Y�_ ����J��uO�|�.�3���fK+:����e7x�諠o_`�[x�Ֆ Xg}e���B����W����q,f�����iJ/�����V٠���9u�8u	u8ڕCt2�W]q�YF@ݤ���Wdw{]Ju�S����IY�5֒��}d��XP��Q��Q��B��՝Ӿ�Cj*ez@/6Y�b5���fτWn��ϐ�m�p1l�� u<]Y9�L-k��(�Z��L���8� �r��H|+�����C�'�5yƪ�wK�i���-�1�9��$�=S�a����%S�'�s���5��7e�6�*$��tCؼ��v;�*8fTP�|���_��k硋��2\c8%P ޶�]\����(杠)0�[�l�$>�|^�o�#��Vv;�r��>t���?]:;�lK̎GTR-��W��ښz�YF^Uy?{��a��xI�#@�]��;[8�"�ۍ>�l(���`�`�c���ou`,qK��J���w8�֤9�n�\�ICEi5�p?�^�k���y�L�Z6l���)nG���g�f�8S�|s㨛��]�0�[��ѵw��3�6�p�1�]qS}].M���ZF��6���Rg)��e?ׂ/K]vq��f�]����w�$�7�}U�����f��������烝 �"�{q�X����(�e��_5H���}JH�����≊��ڻ��}9x�F��zj`a⋏�GȊ���Y=L[��#�p$f�#�ס�6R�<��jy"��5�GS�QV6"���Av�J�1��>pB`��	��sZS�������C�F���:���z��w�aMn��g��Oh'e�m�*�(̠�l��<�����G��{WW���(�������v���螒�}����H́(k�(��Z��b&�/.A_?��Xf0��ʲ�]_O��O���
�����VAyi� ��YBF�����f���eTm��}���C����� Oi�ѣ��~N�y�k���e9?of��5UЩҩ��C�S�y�g*���91����lf�b��2w�R��}�3"��P(��wXj=uJr/�>գQ����:Y>�z�3���5���Lz��>�o�ϲ�9��� 2�S:?����Y�P[�M�Q�Ϙ������%)�[6X]R6M�At���6_J�be�l
>uU^wit��XW�Oh f���9�Z�V���mʔ�T\����5�Cw7��3�Tۂ@��W��.Jj��!���{��>���_���Q�
�؃�fH��D����iv݆�b��M�4��gЉȲ�"DԲ��)N/<�B4���B�r4������}u��gV6�kM�$�F�&d�ߺιL� ��]j�,h�%����ݨa��!OHn�z�K(���5����3�7h�[o�*<���)M����:�X��`!I4p� �� ��=t}/k�Eמ$-=�.s���O�&�c͕� ηN���'cNO������x&���|���i��Xf���H>1���*��$�&n!=�{[��N��s�©�D�����/m��Bc��$�)�|,���S��f1�؟c�;�����?�:� [����^I�_���� :E����r�_[�@�e�3��+RKF����j���~D��r��9s��j��,�p�Ԥ�G�*y����:훆� /�nϫ�zj��`�ip�9c��RQ-@� �ծ.�
�Ӽ��~O.3��"s=�8�)�_ �k�Dp����4-�߱�S�cBrg�fv:�w'����c�q�q.�4Q 2�$a��y��0��qt��˅yh����c{�e�����1#H�3'bh�^s* �Ԭ����X�4Ηj��hl��H\֔.�Y�|"2�U��cs�H��f�`�ݰ��X�w$�E2��� �F�3zB���Q�\�UyW3p�N�r_Xi|�&���h2��F �α�.H���}����ޱ�%]L�K�G)e������K��3>������J2 �j^�;����ڈ�{`]
nн��@4�蛚��$_�P�~��u�s<>~�C�a�K>P�:!l�
1㆞�'�8*?N�{�X�!>�%!@I�)�"s\~ Q��65"8^H1G��,C�Z"�D��$Y_.� 7�#�p[�C�]"Yui�+LSඋ��;�`�����9�d�*n`�%C���#��E:6��T������'�ڙ�9��ޯ�jh��[�z<�6S����:*"U@�!�"�޲d�b�`{k\(PJt��OIqa�m�lEI�M�B2z��'*�d;���<HњYݫ=@�i��`6�8"�
���8n���4���DIA��ZŠ�K�Ӂ#����`�U�`�Mѹyv�̡��=�/��!d.я|���5�?Ȓڬ�w�c9K6�*{ ���U���ߪ��}��r��}�����������"I�awX\�jkΌL����O���XaHm��P�'y1y�-�� �^���Rb�����w�Ve�d�� �H�:�h��	���fO�G^Ăx��v�����c�i��F5.�8��:�l<&u���%b���Y"J䀦�����*��kN'�{F~y���'���J����!%�\׏Sη�![��x� ��N�U��!���n�X�������Z�.�u�"��G��2[���f&�˭]+�N���FA�s���a�i�Sݠ�����cٳa.$f��tO7ڔ82�s�7Z
�J����6μ�.�}�%�:�n�ǯ#�l�7}��O�!��[kk�Y>����4B�d~�����q=9���Q�a3�i_@%@���W�j�K�p�ߍo7Do�y9�0`��k\}f:}�))m�F��s3_�W
cg�I^�J\�|鉡��59�0��+Z|@dv)d��ܘ�J�*s�x��*K�o
�,o��n�$����������V���b\���<��u�o�����,0�uh�<��t�w�n�����@>�Y�[Q#�[�y�,�?�{�&V���"7�����"��$�V�o3=�L��2ĘwW8R��z5�s��e��O�� s�yX�2k�j���ޘ\�9g]�$_�Bޕ]~Ų��/��l���#?m�P�#?�=Cm�<�x��1���
��|�Z\�:��&��#}�� �l�S���$�P�ƉU�_�v����J@~��gI!����?
J�T���->)w����s�w�s]�D=(�s�t+�G$C��*\���d�u^�fz�^@�p�.)�L�O�j	6�*���q������(���k����qp9�h��Cw��e:D�Lq+{�ӗ�̸W?���W�Y�w	�������u!$�%<~��Y_Y�W���o�]`�r�U���볿�V5u�B�,v Ϭ��YL�8���E�l&k����C�7񁄞5p/� �$f��	84>��p9<5u�h�z0H�V�dO�,vX��0��_ɧh��^՞���&$�ye��-+�S�ճ���SD~�-�06�z��ߣ�ŜU�� ��}tAjs�,��3�N:�4�P�s�8u�����5>��	��"ܒr�� =��<�3����MQm�X�0���ν��P	��
��}-��r#�U����FZ�5.=n������ZY9�E'po��˛�Tљ��ݼGD������_�Wov�Ĕ�Tn@{�2`�ǈ�,LW�z�U��y����;��j��U��Z�f��c�8V�+�/eV8���n�fj���;+K��7��)������N��||�]��;)܌ǌlWu�5�ݔ�Y�qV��Ck�.��ɛ��4�r��уh̑�)j�9�'!/�5��W���c�(�xy��zk s��C&�2%��A�m���M�M�> �RW����G�X5��ϣ`Kۦ�b��ݮ������B�~<3X�鵥��7���wx�������9D_�`u�~!v�G�
���Ѕ��[��voI~�36]��#��VH�@F���9��w���ܰ�����Pw�@�o���`
�UZx����Z�~m^�&�>W ��+�!�W�Ir,q�Xx@��C�����"�vN�6���qP?yVJ#/?A	s�iD^x����S�)C�#&c����;(�Q{6+�i��Pe,�~�0�o3$WI["�˹ՀȬE��|�B59�=�]�c�@X�E?��<R�k[ao�Ka�O����)����=��y�X��ǘ�*�!� ��ݾ��5���S~�	N��ࣖ������8�z'������U�u��z8}���f�����tP9�p��ݫX�73�5z;#G�T<��L��, ��ʓ��*!V'����?F��#���;�cV�����,������?�'��۶��}%Xe!�`pc�'~wE�q�5��3�(S�X$h���Kx�ۍ$���|L������]�����o[O���!�	ּU����i�+�%��T"�Nw|�*� ���vY����F�'2�E7��̪ˬ7�RYz�}ԕ�L�FR��#��^���^�^q�p!)����hK��GN����h�G�s����nǯ C�����_Q{X��>FLB$��($jД.�m��1}�c����=!��&n"n��/�@�5�;�y�N�$�lIO$���#w��2�
(Ҥ��a�T~�,9�U)�q�<�kFB`������`�S�qp��������6�\��8�����&��F=�)�R��\��9Z���~�u��/�_�����J��n���e���&���b�B��{�|�s8ĕ�z�9����>m����Ӑ��*�6 ^3D�F���r$��i���Ko[_~��Z�[:�0��L�/�5~��s(�������q�� 2i>�L��� 䚩�Qs�E��Z)%ѻ��t�r8���^��hn� #�����
�j*�[���~���)�e&��$JÒ4�J�e��e��~�^�^����^��*�9p�� �Ƽ{H[zx#�����1���!@��)/h$?��\�Y<�3&�F$��x~3k�%XJ�h4�a�ʴ��ݱW�.H�ٴ��?Oǝ��+���D�d*Z���Ⱥ�BO.�k�m>L=e��G�;��pQw/�P��6m�p$Y�9�u��@�x��F�a��5��b��f(�Fd7F��f��sh�9��aCW�i���ry��+Os�I�M�v�'���*T�]Z��=�ܓ#x�[v>7#�a�,֝FE+l}����-�Ka
m3�s�"a��Wͤ��?f��Q��;�9�����m��zr�O6�O`�D���;Q���x�9<;�<+����L����qG�t�rD��lX��q�e3�-J%6��0�uUXj�J�n��Z�%ރ=�X8�ů%z�PuX$�R����������$:ψ]��;(����r�PΧ�2n�Ҭy���%�li�t������������V�����KI<�Zm���&+Y�u����=��]i���B�g��`����i�r���|:z�-!��J.k�N�����Ơ�É9�������Jv�� �t����=	�3{��ŴQ$g��X��$��]�X���>p+�X\������JGxmA~�j��j�?|ۉ�ľ{��p3,x���F˩�o��ĳ�D�1`�F<,a�t-C3��=�|���aނ���t�W�J��X�m�ּ�,FĲ�n
�5�gi���� ��z��r��ű�b$��=��xK�Jx#�v�%^кHLȨ��zwN�E�F�����E����u0n����y3530] 	�.�_�d[q�������^tڐ:e���e��8"�<ڂ��4@O 2�EW|�����]�>?�V�x��!+������T�5��4�d��!�B��`{G�=Ww�^��#Z�
����Vg���@���`S�h.&���(4B��^��D��H�3�u�1����J�J�F)��'��_F����v���/�'��T	�9��Mk���h,���B�p��˴
� �t�������:�Y�âA%����j�����g7���REE�=�<���l���\@-��9�]		H�/'�
;�h�,����b&�Π�u��r�� 5T�촠_�]�s<���3��?��K������E�I��)��ߚi�N�hl���5�~���5,Y\�*���w2���WЃ=����Ş� ��j�����d�j����IM��,�=YL� t0�2��nQw��bG�W��P�� ӫ��B�;i?�z�WE���TG�A��[������8�3�M�8�~�3]��w ��!\��-�BFE����+n}��A�}��(J3zY�V@��3��T\l%��#K	z�YRh$�����Y��F;��d�a�_�ڥФp�VUꔃx��iZ�^��8'j7��/meD�	��_��Y�Z�k����<��H<l;9g��^35N</|��)��φ�	_����I��z�h�է�JSV�v��e2ˀ�N,{ߞ۬�x����l�߅��"�5�\TB]`�H��XӰ�#R,����������صf������[s��l�������۹j?�ѩMs��	hƲ6�)��h�����N���U&�Qi�6�����&�>̼CNL���r�Y�7+��$j�Wh(�Gpb5��-��i�
��d�[�a�&G��Tf�0�Dn��F�0��P�Q���H����6��:�Ψbo���K�@���Xwt���g��Ŕ�4Kv2%�i�=�Xw��X����=��2��e�(ΩF�v�xJ0�⤾�L�����v��^�HXp!�����þp�7u��ŀ�2'���#%)aH�;"Gz�� ��~!g� ^�3�j�� Ѻ'e���_�E+��w��fv���+�~�,4=B�^�f,���kѥ=|��Z�&̉��^R�j���S�zm���v\S񣠠���a�j9P<p��E�q��<��u�v#��ɱ�
v�BgS}�˾��T�'R��OւS�A���}6���ٹ���m39�,1��ϗp*���lm�]��Jo�+[A�#y���N��=��6��Lm޴��,�LQU]�0�<�䔵���JF���-��U� ��Q��H��Fç*p�x:��n���@IĞ)���WL����ۯ�{�)�"��|~��gҊu�tȇ-5}�]q�v�_�v��n��1�l7��2lQ�B��N�wp�x������V�����j|���IV����^N��W�{ �QU2���t{NlԿ���5�,��کW�& 7�GQ�����,��:�t�i�	���GΦ^�����v����=׳.|Ŷ-��.)\���5�B�rnMrl'�3j�{���I6
���~A�����C$g�xX�[EM����_�u�
"�а��K����VQ�`�6�A��^��dz��"u��Rhi2�y#jsH���Ǒ%��n���l���٤A���_`�܋Ӫ*��IL-�W�8�
�$̓�2�chP?7�3[�ӟ	��~Ëld���9�Hu��{�5�M�+<�#Y��5��Y�YRFF��ؘHJWn2ޅ�!н/l+tgۃ��8Un�R t�m�۵ߵ�f00��O]�$�������;�\ܤi�DlQ@9Ga5dݫ�-~W�2�$8�����|8�Q{��=���2$������?T|"�����Mp�e|�\�� ɏY����
V��C$����̾� �=Pf�Z�z��|�뤱�*�d�6w��p��|�Ũ�:�e�U)߭�;~0_b�p��m�c��m8/���N�-�������<������c�N��w>/�|�g����Z/J[��T��|��Y�/���ެ|����o�D�� ��$�<��~՞z�M��Ŕ�M]�P>�����]����Yn𨻨�&6Ѝ�ƾ�nP{<���z�� J:s6%;oʡ������8�1��#^/�Z��i�S��o���cI&�m�Ֆ�^O�r�V$�\y���ƫ)�B?��ZE*}ҬM�����.����/�<;��Q쐴¼�}��3�>����^{����戄� +0P`�=ۺV��7���5��A����a�k�y�շ@_j��q�8�k���7�t�j���n����gY\��/������T���	L7��]��
qt���1K�C�� � ��!����I�#��f����^Q-�_W�R��(�{�3-9ͥUډ6�(ٮ,P��&>k]H����,������$�,e�
C���"��~+�#�-0R�
��_(�ݚW���f������%
$0�g8��k���aG�P�����f�|���ɉ�>���;�+�}2�ò���gD1��E��2�QIr������
Ӿ�P%P-�������-}t$�-�&�������Q��P���숪v�Ն�S)n:� ��X:�U*bD��� pLY��R��`�r�mW��B�ɮSa�k6_�,?���}tk�p	M�dbJ��˜��n�@��T
��]"����d�*���O�6�g��|��Q�ȅ[��*�Kd\�і����ԝ,����=�����E��$�/HU�V2�.�f7 ��Ǧsh��<XB��j+[E��U�o����֊���+�?`�ڑm�'c�����mc,����SS�]�tDb�R��/fΠ��k�U�|ngڽ��e^�eMTVo]Ci�%Ŕ�k7���A�(�cV%k���UlS����0I�ǵ$��U7�=f4w������+�}|ۋJ�x�ϲ�]X��6��͝�e��,Ȃ�A�z���:9W	�'�x�)T���7�OĄ9�Yn{&	<���.�k<ygҙ�dGe�@�8���-����U�s��H�͇.}R�#�_c���fHzKgn�c��.$���%O���@�3��c�,B�c�J̎�Ϭ�4�g�ys���F󶌑����q��������wa�C�&�Ӿ�~�z��zb��|tT���+�<M�`ø2iL��Ĩ�Uq����vaS��)�A+߿�R��H�~?G�z/?�Z�΢?ZV��ID��K�q��$jvHh�L����z�I�%���F��F���O<�$�����!$��m9�c�۽�O>FB���щ�w� Ttw�d�_�G�Ƴ���M� Z�4�S'��:�Kv��m*i���n��z�u$�-�ҵE�4ƨo�Y1��C��V4��;pZR����Q|���v��YwV�)�i+��J3_�QK�_u�J�u���n��Z+o��XHm?�e�d������j~�� �i�\�p��c��-��Fqcx���'�����;,�,\P�3�0<$�!�4o����7�ⰱ�v!��d&l,�cV!\g/��ݑ$�Q��[��9���P�����y6XO4lu�j{C=���@v�0��̘�M��%ԯ]��U�x��I+[L��C�����^
�ƩLU�w�����
!�1�X}���A����M��N�C�"�o2����qF�s_Ng�D1 .\i�`0�G�҇ Nd��CEu;��U�	$b�p��f�L|��������d������u���l�	��L��7z�]�@�a�ad�/�^R��kp�{�a��ptL��:2Ey��u�xN;�r ,��p�b7�6��(�,L�^�{�CŔy�o;�A�#��x-�2���s38�ْju2g�LI�B�.�Z<9�tp$R�(ܓ���Ț9��=O�Qq�c���ߗshC �KG� H��)G׶�`Mg6�K�uP�Őn����).`��e��;�$�z[��32�6��<�fԴ��d
R��p._�y����`���_��!2ѮgJ�O�l�p��TH�Av�t�oӗ�`Y������V`��:��	@S*�E���<*�uSe)�7G*tZ1�	w����-c-�.�e5���配�#B�*��V/��0!b��z@�/q4�[�{Mx ��]�kSƗ���Y۞]H�-�ň����F�oʭ��*6�9("'4�L9���Oн�5�T���	��� �B#�ݗ���_@A�N�tu�t���Mr�GjxQ���x<�P��3�ؒ��J��	r�3��)=�`ಞ��uS}�^�|1���v@@�q�h�����c"�; ���쫞TV� ��|z��u�)5���V�3�~�̱�b�:e�dh�p�A���|Y��Z�'>��2C�v&��+[/e����b���x�8�2��R8����2��M�L�%�i+��)�X���w�e�2���Zk(ק0���[ZA���K�����5���lMg}w�ڞ�X�0��:�K\3l�D=�����Y�=�\��fEX�=��%��qcX�p���Q�Ȱk$��:�,�����kr��C/y�@U^�ֿ�s��o�t4���ޑ�/�zo��E!�%�h4r:e�d��X�Gif�]F��F�|��1t������A���!�.'�GJ�,��k�T%,��0s{�dI\�X@?��#�^4p'I��"�ɇr.QȐ=�w���fj��J\��2}����>Qm�P�����>��2��ʿ{�(�5ے���=���/#߰#��y���E��De�{�_٤�������X��2��x�\E�K�Ұ4vlCP?�֬[���JQ���v��N���%3JK���Q�f�!�z�7Qt��`eDH�a �|�v�
�OFC�N��I�q�D(�`h��%�֍v���iTi}/t趦S��E(/���˾RCI�6�}��$�wTt.��
���Gm	жWD�Y��}N�����1�U�:����E�ɾ?q��w'��n�2+��9�ܓ,s��x����4)���	@�`XO��C�
0�C�����kˇj�C�x�����aρ��1���=L=����q�P�ߚ�lh�9�T`rO5���R_⦊��W�7i�C�ƭ���8;I�.�3�����h�uFi�gO��`�5*N�IZU
R&��O��M\/�Z��� 9��
�|���%�- 6�	Y�[o�eH���ˋi��%�a��u�KF�͡��U�ζ�dh�L��G���yv��ȏ���:��`x5OL�������Я��'z�1
�r�NS!~�����i��V7���@g����	��^����J^����3Z�V�\s2�޳S�T��U�>�Rbj�b�H�X"]7=�w���Ux�O4zU����7q��c*�Ue,���v���~�n�i��	�6$#��#��ڻ6
(veh��oP�����;ze&�#��|�5h7��~���|Q�D�.g�W6�� �s��p�T����_/8X��y-4�ղ�=!u��t�=��(���T���znrp%w�Y��������X8|��v���\1�FO�W��F>"$�%���6罗}���c4�"��_G/)���nQ5���Eg�BOM��ec�J�&�e�����|w���8�����+�A\�5��dd�5�Ө �+���fpx �\ŏ܃�j-V�Pg�<�V8ռ�
=�B~��Q0����������r42��sxA�y,�fp
iٸ[�uQ���9J�@Q�3jL�M���G�TF��4���][�P��M��q���'=��I� ����s\�������m�@��P��ɑ5��9Ղ�͂O^W���<��i�&!(��̉��OJ}����Ș��'��MʟP���,H�����Z�q?ό?Y�p|�I�k1�>XV$�%O~
���g�>	3}9��rTJ�:�9���}IF�q�P��`'�!���W3�#<tK� �׮�E�$�}X��=�Y�%�"7:��2�U4����o	�=hy�;(D�@#Et|>C��[%S���ŭA%������'��B;F$c͌�I.�"�dh�"�W&w딞瞸�]@��`�(�UZ��� �t�֥ Qy�o�CG_�oE��=�Q�D�Lv/3��XZ�T���'�V�4���u%��)nt�j�l	�K�H��_武"ݴ�K����T[���=Њ$_+_K+��� )C�nH�IA_��0�8h��%WR����"�c ��MtԱ<�C- ������i�P�N��=UA�<��V�M�~��I���O����quGWA�ہ�3��}`�?gI�x�|�{ ��c"��$ᔣ� e��t�{���k�I�]7�h�-��~��,b9ͭT��j�[��-J�&9�DK�Ip��4����+Y�z�&.,�xOŸ;j�Z�~1r. �`�/�(k�>2iprI��Hln6p��H�T'�ikg�L]6��PD���>�)3������R1��dC
%��=/9�]�馕o��N9�:���C����U?f���)�iaDW�m�@�qL��$R��ǜ���� �~σ�<�7t"P�'��H��N�{S��.հ�]�����i���D��$�6�VT6�I��)"�+�be�ƯTD�pQeq�^�:�� �:����5�"J�Z���o 6~B3�ҽ���qɿ"\4���Or�z;�RF5�J˛,�-�M#}.X��Rx�,��<���������F��2��q�bg��y�y@���=M\T,"�Raj���K�s���X�hH��yk�5�E�{��-���Q�6S�Ĉ󯀨��(i�<(�}( [���&!�5}�hi峷�H��WH,?�ں�����ײ����"�\4c������/pQ����B�� �i[L��0�r�gqg��).��{g[�ձ�ؾن�3q#���vKA�%
�.y����O�P���gA8(�Ν&�������*�n�"6��7�/:,�k���O��cr1��d��$���5��?��KD$e�-��׃<�w\ݾ�bp!�I�\�b�4a���0�5 RgR�0V�]N|�E�̉3�%Rԋo���J���t�!�K���2hH|��2���L��I��y�'����;�����������h��" �Lش�6 䌪��ZG&Z`2����<n�c�d�܎�v� Ηv����}ɸg~~}M�kj�c/�5c�r�e�9�pf��~P˅�P��u ��	Rg�c�(q��ЪvWo��u1��/vȃ>�~�IjJ<u�^�L�X�K��"�?�|��ʞ��7���ؐ;���.r�y�ஹ"����;�T[ƗuRl�g
m�N
���[o��F0�f�5�'�>��~ǀa���)-�p��c�b�"�9/7b'	�>�N�C"�+�7z�ԛ�K"g�E�fX�è�V�A:�=���|f$i����q�Q�R����f�k�K��Bc����W�?̆�\�O��ޣ��gw�j*��)G��Ja����2V��2�\f�Ɠ|�r���Y�/ƴ�s);��e0��K�����L_����o���� Yݳ,Q ?�U���x�a�qA��\��I'�\��n�Hn����t��ϲDk^�@��פ��%�<�0)�?TG�YRMû�Y�Kd���u���ͤ��]I��E��j�¾=rR=�*�d%M������j:ŗ7����o�5��@�+����ea-D!&�?��eӭ�����ܯj�o�W����c��5��s���b�m���a�T�f�ٷ��.�E�!�:��4m&�e4p=BH�?��t�����a����2�2���2C�����k��j�j��+_�ۺ��������c�tWfh1�/!N;��c�h6f���"��#٨d���}3YA�O3����k�5:�1>���O��.��ͻ�z��$�Nj�8���s�����j�t�W5����ed���;h���r�sy�E��Ex~�/���|}(���="#��D2��R� `��LAl����C�ǟԈ��n٩���7��W���{R��Q^�=2Ϩ~���aB��P��?U��ۢu����B��z�']���tJ�rDrl�[uL�Dr偑�k���f�
�,[9͞N�	��%��.��yP}d*]��N:�v`�^Y
�;w��b�;Ra��x���	�]K�(�Ah:�]<�t#���2�&dNQA��@ƴ�{�d�p��۷>G�"��,z眛���v��#޸GB�3=*����)���1�#S��u����|M���O fƳ���]7
u�%>\c@n�U��7ܾP�d0���
_vp���W/}AYa�t�����?=�lE1��ߴX������ծR?~$�x#4�`�ܼtMX��l��{�am2�:
w��-:y�����)Ry��ޠf"�J��B�I��$.ҷ!]o,|M�=���e��y)��*��l�S_?.�`mC�I\��s@6C}�I�����:�yM�X^�:*�x�?��S۵z¦}�wD0w��D���m�#I٤��ΤD����A%z�O&��9��J���Ϋa�X����qeL4L)�.čK�8��>[ km�����E���(g�xs�3^\N�hq�)Y6P?�����!ĉ0,�Ie�֙���e���N!�T���ME�NMAT^��j��VR)~����\��쭪�"�����ϐ���x�y���p1c�t�Ł�#�?i�r���?��Z�of�\E�埜��֟uJ�Ħ��Wj�U�s�E_]�y�U��L�v�J�M���_�_�����=o�FzQ6�����|��k���Eۑ�I�q�bU�֤�^nZ@	��e{�@�cU���?��������V�\�PEELȽ#��+k��C�g�z5���)KE;4���M2�'����E�m�E5�+b"g��ϝ��;�4�5)dK��2���lc6����f�������;4	�aM�"�y9�iV���5t=��?	��3,�|��&xJF9�L\��ڹ�Ƣ�n�� 䔉�Ӭ6������\��A��@�Y��L.�H���"<�$p��~�
���]#��m��yyap9K��BB��26�n�����=!�Ф�cR=��������؊C'a-����*���~J2�U�6H�Z���ٟ{��F͑5��� sg!���I�n?�2 �8����5-�����~�������#�[hov��Ɨ�6���$�Q�̿ޮz'�>�@��+�h��H���`��Ȑ�M2���;���<#0�sAPu�"�'m�ű8RC���2�CP���0D_?	��ndk͎�����a;�1no:Ů0~(����A�l��8\���/��NKX7q�J��P{E�ь�1V�5�G.AGo��%�QE;�����a<
?��L����L3 ������]!����jff��Yz��s���i3��b�3M_�=:�S��h1��-{����p ����:ɕ�It�N���t2a�R9�l
��	B±xk|��Z݉����"m}G�p�E9]�����Ő�H|k{�����I+�����3@����G|�t]j�)^��`��ё�R�p1������-�I=^�L�;3���% �Un�D���b�mDp�-�mVI�e�O�O���`m/��&B����2��8/l�]z~�D��~��J�@yK��P��u`�{L�cD��	3pу��Ԣ�o�AԅC"�0p2Lm�fJi�g2����W^��d}�Y~e�"=j������[LL��r�Kt2�lق[^�T$�[�`!]D�Z+5�} �9�`2�N��R_�Cc� >֪��?Q�x&��x1n�? E�8���ec�J� ^o�@:�?�R.��$)�L�E@/��С�-��<C�CPo�T���R��jP��|���ȧ�d9�22�W�P3榮���6��'P��?
�u�Nρ	��� ��L�`1����F�;Ѣ�:Vb���ȝ_���ȡ?��7c�{�5dChzи�e��fhl.�ɦ{o�o���!2�L��S�ľ>����W�Ioz�~�Wb�d�`�B#�M��k���R��@n�W��
��Ǡ��>�n��a�	WW�[U���RѕN�����$�>��6�߿2v��m�+�88�t�t��BDt�ַ7��"��v�j���r��Q O9%I�r��c��w*Pu^�ߞXC[6���L���j1p�� B�	��D���y@DM���Kz)�=Q�3�Â�Z7S�<�0�͏oVV��"��ɫ����E��ӱ��!�T�A4�D�v;*��ؕC�P.r�m��z���b��~�
h��p�4�g�4%�>[��{��g����5"���V��o��o"!�bCE�rT�۶�	�!Jkɼ�k^��
Ǫ�q�4�L)&��AH��Oz �O�6�&�i��]&$��1�^��W�t�S-a6V>��Thmjk��^i��[>��BBb���FQ�B�����F�-���3'��l�)SQ�P���}H�)�R���,�w�|�<oܖ��M���.����=:�d�VU��Ir�T$�#�p���n����A�%��K�⌇�(��9���@���('i���D/|����Dɥ�V�-�7��մv:��������"'��`d�tK�B�p�"��i���P�W�X"&�hm�-~4я�;�w����V�Ǵ����f�nk�u��)ۉj�dC���ቸr�.Z˃����#!�-p�1Ǘ5:ӝ�L�]d�7D�3
wD�,0���cy�2�*>̲��Qi*=����RB��P��BLk��6o/CZ*`�!r�@�rB����{r�RCD��u��n.��R�6����<����EC��u���Im_�[U���t�&����<j��MR�p;u�s��IFfd� p	��u'J:�G��{G2ڪ�e<\�p�fB�d<����������?�/LȀ�׈Ud���+��Ml .|��^�PNh���� s'ꮨ�|���!M:��ž�M�
Um�x�o�
���<����3���T�`l����q�B��k&��9E3����]4XC`~>Y9�B��9�|��o������q-;��æ7M��@�_����RF��^5���U��K��g�H{>���Ю��w�;+�a�'Z�m��
��
Z�ʳ(���'X��2h�4�M�}�T�����^���� �GC�������X1i7Z @�Vy\+��U]#�@��1�)��Lr��YM��^��d��G5����'V�Q#��Ҩ�HaebF/6��<�r�S'���.V����,h�ag1|�
D*U|{����ZNWa�Tp�8=Т��n~v]�h,Q�q���v�c�ZO�\��ˢ�"�4J���hM�����y��S��eޫ=N�pp|���F��}b �/A������K�L�3�jAh�'�ܥ��b���'�~�!�	�g?�Use<���0<{��7*!��	-���Q:C��J�o}��߄*r����h￰��(��'�v���\���At���v?����(qq_�A�]�Z�2{�$U���ep�F	��N�n3������o�._ ;>��e����uw|ltn*E�N��5C
Ֆ� \>t�'Z��WHb�/�F��i��B8�� ]�XC�ݨ�z�<:���Bgв+[G��j�k�Ƞ���{�4�L`w��U��h>?MQ�G-~GW��t�#-��8��i���ō�Z�=�`�@�l�P!��YF�5*��3���OVF�Ǚ��$�}�����$l=�����ݒO���ɋ&��gKd��DBɅ�'���x�G�	YA���w�v�z�u���0}I�l�O��&�-S�3(bׇ� 7i��=�<�_���cɱ�����m���7q�4�BŃ����<x�ȸ7�v�`kI��I0�܏�`�h�:�g��A�rv2>��d$�\:,k�>=�Φ����4��ǯ���W�QKS54�R�k�]�Y��z�>3�J�6l4��������s-�yS����M_<�I������&F-W�?��sg������0:�Ϝ2��������(�:`S]����)P5x'�r��C�0��I!y�d�.ߣ������չϚ����Ӛo���QJ�\&�b�cӀΫ�
�mb�9i\?�
�R��w��w�2�+�H9�B���C��p�q;HJ�@9A%M)���_c���k�����ū?�?�s0�u��ʼ��R���G+W
�f���1�K1�v*{�8�M���!��Ht=n��ɑQ�%3c����@��!�Rѭc
<�)�j@��OB�vt{�n��ꛤ]bP*8���κvdb$�L�͛-�50?�˦�N I����j�hI������{�ܖd,�G�̞��i=i�8�x
�m�̿��h�<���;Gjhu����r�~l��2P�׿�<H�lg��Q<�2�;=gxո����
�~B��0X�&�Tn�����˼����L~4��5J��S2�Ԟ�C�O�n�ַ�>CW�*OP�YJ¡|�$�h�7B �:�EO�b��]�i��޺���"�L1f̠x��jd�{���|t����� �R�0'�&+:V���Eߴ�\������P�+��Ey�mȋ*�c��5�%܉ F��C��H7�`��4�������^v�1��%B��w���λ`-�KV��Y�$��i�e@�P����@���<���!�9z��B��~	|̗ԭ�x����)������e��.��Ԓ���Ix�_E{�3l��.�wzE�Wj��^`I������� �:�_O*�wtUeC��Vu�3	�7kܣ!�������g(uZe.3�H�:�뗥c��0_�o2��;z���`v�t�������f��Ǻ���n�o�|��W�P�Y]��K�(8l`���?������}��P}�V;fK���x^'�mWFU��AU.z���[0=9����exNղ��W?.��EYK�W#�G}�[b���@�9���qp��@Ku��FU�8(Q	��:a3��������E$���T��:3?��Ϫ�ti�T7
�U�z{�c��e�R �IG%�En�M|��ᑮ�þ�_���
�`�7#j8��Y*�M-��T�*�EX �8�$�g3Q�c��n)����z�F���A�H|�Q9O���^�_S��х}K�UH$���Pܗ{�/ݳ
��D��!Ǡ�e���J���5m��-�o�{5S|"���l݈ ������.>�͈���xz2��up��`����#��B�ط1P�4�y��pz#�B7"�dM̈�ۍ�f�����aOa�e�P:�Y7M�j���Kh!m �%]�W�6�|�*= \Sn#�H�����+{���u��S���J�
�h�l�f<��G��6��HkD�\�/|~�o��)a�������X*��,�U��0��TGl����̨FGo���{��	��ވU·k���5��x:�. W��������1�$�טv�>h��QA��WA�0WP���ስ1�����K)7�95��ZZ���C��sx�Dhʫ�TJ`F�U�����r�{/0�6i�m��>�n[�h�6���!��Eh4%���o�m�ʆ�#/��6�F���^�+~>�˱LPk�6s���+�)�	�3�+O����Y�De���V? ��yԓa�(��,Pԉ����C�	�e��m�SX,�v�L��"���Q(������#�,U�2��j�!��A��P�6�	��Y�9@	�n�l�I�Jmô�ٌO��b�o p=��RM�m,#�c��T���p	�4���/%��Ak`�	ϛ��dGmp�e��z�Sz�ɏ�~F6��wb�{��xĖ	&u��ZT0-�,{�p�9B��>B�UN1ϝ���w�DW��@*8�Z%a�EGg��%�M�Q��o$�Qm"��!i�!@��K*X�e��{�zV�"�3~�6���5Ӂr|�l��'�ƀ���$i�g>@Γ/��w )��:�,�n�u�����S�3�M�`�ӱ�xOؕ�����������d���o���&���lvk��c�3t�ɾ\PGQ�Ѓ�QO� �W� }�iGk��I1a0-S\�h��ez�,���x�,�s���9�L_#<��,���k؎�=P�{V����8����G�� ��M�F9�GV��N�T����߄5Y�A��sl���P9sf˒��/��gXF|<f���v_���O,��~*`	�ܓ�x	xfx/הa�<���rc�a���xӔ|���Q��������h蚸�J�z�Z�)�@�Ku��'��N*rz�oc�6�M�	�RI�;8��:��>C�{>.��J������c�mq+x��k8��j�[���,]ti=m%��E�Y׆��,��W�4ُO�M��@�5#j��&�r������n?�.T[�,3�3U<��yu ^E�d�����&�� �l}��B�IQ�2��-�{NY���Y�ԳeBp#��:܍��\�7[k��G�kw��2�����/d�(2J�e�;�L.���gd���APgi]-��������rŌ":��%�e28� q����Q�*�f_���;�n�^�]��Eك����z����cɧ�nCÇ;�y��cY�h���>,�nLא�;� ��ޫ�l��x�R�q�%?Ry�MLP�?]1M�@mM���=��`O�zQY+&|����؞�N��gi����W,(����|t���p��Ғ�Y���D�N�7��K���DA�S=��(�ڱl�}��8��/d�X`�L�9Կ`}��H!4��w@���>^�-��H�D���B��cLfr:���vU��➶D��rC`Ȑ���z��-u��u���e�#] ��48) �"IxNI'��7�
���5*�*��;Sg4�����{ځ���;9?	 '��ܣ0h1�ÝGWc������)[tu�'3���������tS�=�We�a�]�'�[�'R��^�.�Y��49��#A���N���11Y�Y}�I
����4�Z��r�D�!z/�V�̅z�`fْ��[�?�/g+z�*ݳI���s�{���>t��	=���K��O�$J��8��ߛp��[��WN��N��-g;�hp��eݛV�Xo���%��/�g�}�|y�g�^�K.��|�L2�hP^���O�'<y���1Q3"z3&
�|�
���(�}<�Q�Op�JɽHf�,��ؿ-�����%< j|�n�K#�S���^���ѕ�ӯ��
>�;f��8
%��v�w�.�`�����Ȅ~�Er��B����U�b�\g����������׼�I��oQ���)��43X����}�?��v����i�st?�̖��<؇�n����_/K59ؗQm4�ׂڸe�	�����[$�ig�5�(*80{d(�@Mx�vU�dc�6Knҍ*/l�,���^ґ����h�r�bg��9���F1U����UR�u�D��;{�Z�D'��sMw����JJv57�e�ż��*�Ԗ�ŘY]��n��P�Rj�h?���&�!�ܖ�P����_�eV��(,��Zw���Z���% �51b}����_#U��]	�1ʮ��য়>�/���@�Pc��ϡϳv1�0������HY�'!�c��[�}i�Bɛ��dΨnZ�U�nbQ"��Y�\v}�d���9�x�|�C�Ϸ��s�`TlJ9@���	��v3����	�ʤ��l���N�����<k�S�;��'׌UiB���ufʄ�J�8�D\dPb�V�g�����m���_>3�S�Y��8���	Ē�:�D���UX��������O����� O±��
&�ù~\T{ڧ�,�-��q 8KD��ѓ0�Jh�u:x�"V؋N�x,D�ҩ~��d9��C�@�~#�РZ)��D^E%p�ʴ����<>���RtP�]��p+<C�0:�Uղ�3(]d	i�S6�8'�mXbU5�Ct���t\�N�F}|]�̡��E\4�h44��>�s?��;�K�z�"r��ĤLW���sl
��qm�
3�s�h�oS���3Z�!Jc�q���_�����B��O�d[��)p��ɹ��i=�y��P��?��p�������k�V\�IE�� ~A��D�Po��"�)��~�*K��۠�����8�R8�_�Z�f[p�i(W?W�#�Aep){V�F��ƛ� ��8�lL��m˚��Mlধ��;�q���'&[��c�~�S�@}K�ų�[nN��ζ!1����4�Mq9!1�ö1k�O����#א�`k�M#*<RƂ�3�Ӭ�\�������}��uɍ>0C ��r\�Fب���g�k>Yu�yB��2��SWI����U��}��˞v������P��68�8B��ۻ0��܏���B'(_��l�纂��Q5�r�o�
���] �[27Y��L�l��ZC����?]Td������=�\��+҅%�Ҷ@Y�_�|����K�,��#�&�� �� �j�
4F9@i3Z��FD��՛�ZP(��n��gZZ�$�~�T[��$�d�㸋^�p;���;�|.hȄu�w���肑��Xm�3��H#�a��#P�V�����Q��k�F��Z�.��Zl��p<�Zc?��؛�$v�����0���I�	Σ��&9�E�Y)S�c"eSP��]J?�ʊ�Rzg��l��ۯ��4y���H�W����ύ�<��qP�iP�`f�&`{���w���*�k�n���:΅�G;����X��>��U����
m�-�����9�AP�q=&�cC.8P2�N����j�Ȍ3
d�1�E��Ү���E�Y�aH34�.0$adޓ��TO�\���~��__L��ę}��>ȍ���<����a��9`S/�n�[J����=�'��S����
2�x���Up��o�ϲ��X<��������O{$���p�w�^��dyi1��Օ.!#8������WL=�I�����G�ې쥄p�����1�׀�d�Q^��1�	Y�jF�[�[{To|��&>�C�����?A����q���E���Rj��gh��L�,f0� 0�K>#A�q[+^T��V�P�.�Jr���9�9u�"�{^�@��:��M17^��.c��bV��u郺[o�wm�K�2\\q��ί8��t���!�� �;O3�G��(*κi`�
p�w�a)��0�-�A��M�� ��%V���kD��M�q�~iut'Da�f�o���Y0U�v��P$��0�������9��x�bi��-����U��H�S�qGd�-�$�y��y�T����Z��j���6*|��	�g��ߕa.��j�-ߛ�`���@U�2&���rS�\_�"8>Xl�ݪ�H��8,��<J���X�%=�Z���m�L�g�S)z��hfˉU9�9��I^����P�d�����.��у�ܾt�����9�2�{��U�1����r���vѮ�M���iƞ��\�%���k����|/�Ɗ�jܒ%"`"����5r����T��M�X�f��|e���)I�j���`�Jwn��@�2|��1a�:y	i�˩n`�|v�UE0����N����"��,ޝ��$�l��#���]f��^H��(+ݪ��2O�,��<q�����Fŵ�����>�<����>�Y�`�ߕ���yAi��|���1ݦ������mg���"���
�_���jq�aV93�}��uTe97a�$ݰ'�����,`/.����7#����twY�NV�Zoz]�F0������8��?yt��ީ,�.�+����D��jt�=�
��>k���$VOg��J"��z��Z���� �@�R�9�5�K�N�N%��Ҥ�,�[~�x�d��m��E%t��Ȏ����ϛ�
JKt�/��44F<QnB�6rn��U�����o���YI`ٯ���2?7<0"+co����Su��`͔��9��S�˺FZ{�>w���Y��E�Pa"smK����/�����+ƍ(��*pѷQ�mՉ����Q)�R����� m5B��V���Iݺ���DY9
�E;&���m���?_�p������ +��9�2��YI?�;-���į[��ً:�a����[>Sd��7#�sc8� io�XBv�D���;g<�\��c�K��rOQ��Zi�,A��hMt�k��z-�x�*}Τ�̆@ВL�L��'��
��9a�����^I8�Zދr鷃Ju�Z!E��D�{'bf�{s�_���
.~xg�h�
����:��i5C^�>]�=�QB�o3\i��
��`B�I���Y82�a�Xs�~�\�&K�# y1^޻��%rcMr}�������?u���x0>���>���
��-����Pm7IV}����C��9��/������i`�(<����� *W	��W���Bxb�?{%�kV4Q;BS"w&���_8\�^EK��W�Ɍ���p(�ӏ�>x5?�,�7�Ug�Q5bϑqA�v%rul̷V�$�@xp�"�%<'���n
��s�q�޿��"
����e����4�/&�<��a!�"�zLr|%�C��^�����'N�Q >���#��L�h�#�`�a���Z�:9άgh(mX�q��h�u6j�\�`�lW�o���I�{�]Θ(�B���U�%�׺�XE/�_��oMa�����D��ؘ��n܁�r\��ٖ#V�d�A���@�x{�#��e, `��OkFT¸g�U�G�θ[J�D�zKO�6�{]���wr�m���sX�JPw����D�>_)�z𴿒I���}QmsY.PېT����K��ާ���m6�tm��g7+,��_�I^���#1ݱ7zm*�Y�/z��33-xT���r�6��%�� [2%��Ԃ
�Q1��l�CǱ�;���}h$�2�����@
�����Be�}pK←2ן�=�6^��P~����I��r%�f���J׊B�<*d�>�W4H��2��^�!*"]�Xa���ajၑ���쉠-\�M9t�p12��ǖ�ܵ6W��,�L�+�}m�#z�7& I�^�j}	]UHn>��Qުv�d�_Ꙓ
OG(r�MCk�ڱ_���;i�|��LI�܌��h@p�>��0]M�O�	G���\z0<�����o�B��
�l��H�"hˡ�ԥ��j�h]i��Nji�(��zsC�[�Zg?�o��r�|%��E�7�Hh$����f
�=y|�O�".�{���PK�u�Q�6q�#��Iǵ��@l��|H��wJ�[PB�g��I�^�3`��]�pf3 ���&���V�3�-R�@��s���c�38�>l�{K}{c�N�"м*S���-��Ǭ\T���-6f�VܵZ���{'��\�}@����t����9�a�;�{���؞���cKC�E�i}��@��D��y��_R�ƯU��zuW�/Iݦ�l�5�6z�	���o�+v���������WN�z5�4��	)��gg���O/W�N]D�sm��cQ�cI��wѽ5���������L�tU�o
r]S��Լo�����~,�RB>m���&o55 Si�[����4�w�)xfӛ�O'��e��@omD�Qj�����qNU�y��U�uN��>E�[H�3B��<�9�_̟���N�mT�{ڥ�ȍNbF���߷�!ynE�;�J�s��YE��s�]D�C3�.���7��E��K./����NS��h�}K݂�AРQL���|�}ۥ�"J��n7j��x���\��D�������}(���������Ks�y��hY�Џ����«�ϭ9|�k������XZ����0���v�.�j���:'=�#���TsJ��;���;�K�*��vu"d4���WW��5��B<R�)� �?�s���[���|'��XrV\/���$@�n����E�!�q���~�] [6�,��K':�^I��AƖo-/Lэ����5�q"�R�]IB"ȓ����b�?�H��>�iM�K�{cw6'!��qڿЂ�p��	׋�~ѐ*4ZH�)���1\P���e�Ύ�bP�x k�����)Hu�I�pF6p%L�c@��r��B�M���3�!L���Z�wE�OA�W�t���x�%&Qf�hʘNP:�V�Ԁs��(�W������8���ͻ�71�'5���B�i����*�J��9��D_H����tP"D̄�>a��r�@���Hv����\��:��YK8y��Kt&p$��P�0�k�=����%Yd�:�).ƅ-V��)SS@C9ͷ1�RB�"q�.�2rµ�oW��??��U�L�]�S�������h��b�g�N�h��G[���a�9J�[2Gbe'�s����)ȼ`�JDy��E�^�}�!ۅ�H��wM�� ���\΅�<��7�lQ	;���ۘ0}ՍN�͟�ڜYSo�jřG�C��rTN�J�yЍ����{x¹S��yX�x� �$^ܫ�4�������l�~��~ Q��֪T�CBl��1,�s��B��Z�+�ڟ: �߽����"Y�4��B��j�Krog�94-[�7�
�y���U{ðB�6��H�ݗw��_oVMڗ9`�Џ�M.bW��' ���#��oW��ռIyH��^��r*yHXJ/��VF/��Y����4?���i�+�o���m>���*Q��y��@O&����;-J�GX���.���v�dE�QNś��#��>=w �fx�����OO�dP"U�~�Y`��a����S��2'YP����C����QD��M�X���Ar�`�1�T���t~l��!�%�F����6�ֲ3%�q~Lθ�Ш�NV[&L��މ'LL��F�&�?�u_U����m�rg��ɋ�Uw�o�ހ�}�a8V��aM�:�lf
��t����葃�_r�c+�̤� O�����"�nό��[��KG�	���W�ЁZ���v1�����ٱ}NS������i��9���W|%���)�&G�71s���^��M��o�Tܛ���)	P���C�J��醗xuW����VHU���)��ٰ��׏E;.�yǿ�]2g�,x.�_A;��y̶���Cߢ�iI����L�`���_�����`P!��J\`�߳F��?�M���AOb����{~ e?l�?�p�46jjS���iPmLTIp��)-�Ǖ�]jP�K��#�S�����	��.��{�U5!�ӱ 	ڌ���P�7fo�U�m���	��L�s����)_�_Wj�ԧռ��T���Ʌp��A�OD.���}�3�����\�ens���6!�t��bDK�7O���ϥ�������$���E��	��6�[�ssԏRo�#+e�����c�dو$Q��8�|��x�����Rn~LЭ�EWu�l����k��+��M.�*�1I�s��tuN����G'El�5X�6
JA#��d:����.�J��N�g�YNY��ƍ�j�г���o&���do�,b�W�%vX��N�,�X���MזO��%Ep�F�.R�Djr2q���\u��Tk�?�����WZ�9�L�]� ����3G��rN��2�0��F�Fc�b}<Ц8�����Bf�a)ZC4K,�|�8/ՐGN	�~�)�<��!��>����Bȃf���7�� 	�Y'%����f30�8�sn��f	���d�1y��.�(�wT���{��y8	��j�����.FBN����<#��' +;@��Ż��h�A�_����g�UO��R{-;��,8���Egmz<�^�����·^8p�k�e���G�2{���.CN�g8��B8��9��\�a�T���)�PЫ��$�B�I��w׺,9���u��Ղ4�g�0�4��ﰾ*3r
���ke*���w9�i�.Z�$仈�f|��_��d�d��C�e�{d��S�[p	�q�� "Y�ju����>��S) uJ��'����'��Kvr���k7�ۯ�2OVB}z8�-7�$�.�f���z�/��lÝ���󀀡m�ܢ4Ѯ�?�� �d<��Եu��~�'�����ι��$z�6
�3���џ-�j�r�+��`�-��m�I�|���T��<'f��3(b��{��%~�q'��i;��G�� �����P��-�퀶Oó�"i�=<eu��ݣҨ��OH2�zY��Ѷ|"�Hiz��
YQ�P�t{y<{����	�T���S?*l�	��ceP� �XG`Ñc8ΐ���[U,u�T�	L1�)���p�r�6��=��F���\�*:����iGm�&ƣa�*z��<iD��N��	ۥ�6¾�Ak���n#��YTW}]~7=��R�S�Sx��O��Gv��̣fY����k��B�ܽ��p+��w!��I@��� �����T��)}�o/I�R"�-����ׯ��f�K�J��p!�E���)��@�f�}?Xg=?��������Jj!��$�V���JV?�R��.��;��^�
��߇1!	���6�f�jM}tf��-��˅5����`����,N(�|{��v˾��8؁l�Lᶳ��I���(�_<Ʋp�1�<�vۮ�k�xy�^�����a��쇔ۙ����,����c�@�ڏm2Cs��M�J�/��į�~��yc�i�|����yɯ����/�Xo1}���l�@Z}�'�^6DPʵM7Jt���8���{O��;�.=�������2����t�9�knC���T>L^Ru�:P�����6���0?V�;�Ī�vd~ݏ{U������.���3W����l����v���|>�?j�k���.w�-4��K������ɺ�-��.  ���5�ר%1�������TH����o�YE�sɧ�P�J��j��c��� a����=�� ���U"��C��ۖ+�&{�(A|��`˄'�a"�%�A��ДFn��C��%0����"Yץv��vBN���ت�6����Yr��4��GJ��9�7ZՕP7��Fn�Op�
��a�{��QBh�C���~�!��v^5@V�}�]��wuY?4�homd���SdJ�w��"�D1���p|���Ii�E�X��a~ʾ�� �
�Z8|N���|��܃Sz_�k8�6��.�n�}������N�R9p�`����l��.#�0:�r~#��x:ia�+a_�<��qf�2��Q�#�Ӣ�xee�r��	�kPS1.���[�9{��XB�������bV�>D3���||��'�$\zLT���hz�f"���d�s�V�eޞ����[q�}+����� �����-p����W���<Nngr�Ը3���������vlϡC�6V-`�g�Y�K8�f��W�A��n w"M}�&&�r,�&Q�$�Wt�$L���c�(���k4	�#�Н`�z�l�,˩H��f���x��\��B���sDz�<ojz�6�@|�����8� �?Ԁa������6��;E�(�Ș�D�>�sZI�(I;q��r�'��2�o�-����֮)K";�����s����Q-h,�d�ѡ�U�)U&*:��D�1�#zd�����ig���!8 ط�֙��_:�����[}�" ����hH�8����u�?�d�}�Զ�ȫݲ�â�M�4Q3^��l۾��ɔ&O-T]�VA�.`��2f�'���]gU�4,d���}��������B�26�~�Խ��ÿ}A�y���F��M��v�jҮ���a��*���4=O��u��(c?���2,zG��x�)�~�bg�d���T�jZ���\�S��YtW��ٻN��s�ﻪ[� ���)=8���q��Ts\Z����Mn�9���G�*�e��Ⱦ����A�S�g���a�a�ՐG�������9]�i+�W��I6zE��Ot�D���a���j��	d�#��z��5M��TH��#���g�j8Z
�ڻ(z���*+�`��������G��  ��
��ԑ	vi��-��2!�:��#���>�����dbt�Q���;��J��r���=��5P�~=�[���64�&*r�M�|%AB�@UC���g�{A�M{��h���u�m�!�J���v�q0����D�v9�-�/�3��@��}�ac���x�U
r��{;��uMN��lY��'��t�!G'��ϰ�]�CA����i�Mm�%�p�DXPh��>^g�o�O��N�v/��1
*�͢�K�e�G��~]w.y�<nT B��]Z�A�(�����"ٵ_�ǿ��	 �cl�P$C}�X��\��te&;d��vĕ�!�(̻͆�X΃ ��fN��"I$u�i
0����g�||َ2t�z_-�tێ`sbW��}\;)��	��8�-e�	�Z���P���<i:�2>��窳�\��8M��ݮk�o��l$:Wݡ��᭎h�z�T�s��<FL�MQo�.Z��Ӛ&�Y̤�T����B6N���ߡ����������{Sj|a+���`�K�G�+% �/�oi�H�Kޙ.u)���Hr�#U]�A}���) ���E
u�>D���dwS��%���&V��8Ut;��z�	���*}�H3�7	ak��c��4>4h}�s���uKW6���x[�	���z���#>~�6�lK��#�¯��~��&�
:ѫ`�Q�gu&Q���gܦѷK�ҚR!Q�Y+߈ܐ�vTi]���N:�1�H�����	6{I���&��� ,��d7_�da�(��»-�%�췡W�>�Vw�/�܅��}S,ԹK��j�Z<<�ۏP���4<�u��'B��a�9�?N�ɋ�A��C�3�(۠�;t��(��zn�+�k���X8���*�R��\ ���	q���j���7;IdL�ּmg��z����T��)����ҩ,��TaB�ע\(����Z@k}Zg��̉�p�-�ʕ�Έ\�A^T}�=���������CHK(����}������cӿN�KDG���yH��fu�t���_W��z'�⬓e���=-��p�L����8�8�[iH(��}�3Q�x�S�6��
n�+�$�,�-��g��b�� �)��=��� )c��Tfg��,f����ܿ譸�;c�
�=/� �d��`�ϧ�����}O榧^X�VFwFʦӲne.����J\�[�f��r�+��Ѯt_&w�h�e �ƻT"��	c�j� }�%}��߉����tՙa㺑�K����p�73���̆p㎀pn�������R{Y�?>1����3B\���FV�ܥ�'�ᒝ��v�������?ֆ���Ԉ3�]{��~x�3�6V��5G�n�T3�? ���1��$F=[lYn��j�|+TgL�D�ZV��"�}��;�6_O`�ǎ@��%[����7!�r s��X�}ʘПv�wP�g[�sN�f�ǧU����*؋M;�Q� ��9_�I.�$ɩ� *��V]�w��=��M��[�dd���L�mQM���5}�u����A�@�ӆ�|�V�����Jxl.�/9�Ӟ��mi�޴��Z1�Ox���y�Y-*�h�C���͘�����"+�{c'�j*w���)����n���V��>B1
�,f��;��	�j�*��
�m/\��Ej��;i���d���z����B�}Ъ�����6��}�w�I��c�=��e%m�-Z����P»y3uy��B`�m�6iG�Ч�=�"Q������|�.l+6�Sa[2\�&P �9����>����׵���W$������N/������v)�I�3l0޺���
��ԅ�\_�7�e���{s�2߹��T{��К�e��%�����;c�N9��j�V=<�ݬY����l��w�c"��=�q<%�dW�_#��Ջ$���`�#%G۬�zv/��Ӯ�p�&������ex��)ߌ�7b���z�����<�&�{��>�a�bk|ۤ����V/jV����(�)���ժ8 �4a�1}s��0	:�]�9D�f�`}z��^�Z���>��v�,�l^���M7�Y8]�ٹo�w�S��3<K��[��9�azuT���/�G����F������.Łÿ���� �c�����ޭ��϶�(.}"�Μ��Q��v|�r�{ۆc۸200���}���q���CL%'�F����P�B���$5NK�_�>�����Ӟ���F�|B�V�\�N��B�+��/[m�%L�,�IE� �c�xm�%8?HS��!�#Fj���u�c�����{��T;*�FR�/��f�Sջa�E׭��������&�l�"V�DN��#&�g,�\׃�����r=�[��/8�$��T���R��?�����@�j�S.�엲�Nk���0��]�e�I����a�"B���	[�j���>�X`1k�g���.���h�=W�hևY3��G��>�K�������8�(x����+tΝ��
-G�HC���U9����)�}��DM=�8��	6Wx����ckTB����Rh��v��>����X�uc��3_��ea{j=6�x�rg$��whP�hha�^4��2x�$oYq�*�n{��NDl��i1p4��;	?:j�o+z�܊�h��=�MZ���V.�Kʌ�{�3��I���%�`7���_��8P6Hz\O�3kv��W�)�.!��s�:Z������p;�s���p5fKE-g蟖WJ�_����\1�D�YM�i �DĎ��^C^m��_o�QqV�c�㲞F/�Z(c|Ȯ���zsX>$���SԘs[`�Z
�g�0o����ܻ��l+�� �	�_M ����4��i1`ϊ�a��X�X���upe��z~x��HL�!5(a��n���j��^���G*�lۭ�2��g7�q�|�f��U�� [ͿpqqJ�l0{��e���vDU@�������f"�햣���8��8� @�H��d����;C���E�(~�������\����2-��K�-vC w�S(��������Py��a��ox�6ʫ�̣��*g��	a�܊�S���D8�bA���P�Ar�Նި���%	�F{�����9x�<��ʏJf/�\΍*u�po�'ĩ�P\^����u��� �~ڂ�	�x�4�^%�~�%���J�bۉ���s�h�o)�Y��e0ߙkS�{���Lt�|~oS9�H��T[S���xl��h��"���=5����<�
%�K:���9[��;�u���a���+��U��Y�y�z���}�n���[�9�~S�Zx߽���B���W��(��W̰�����hS�~K�������w&7��A3}�\�u�<�XP�Q0@���RU	��b�a.�J� A�W�ya��a5�ׂB�l{֧]'KH�f]�F4�(�i���R֥�i�䃩���wWM�e��x�=�0������耞n�Ƅ 8O�%��}�sZ���|,U,��H��s�<ɹ�3w��(�˿����!�����휲o*��qV.�䃺�E���:�X.<��[��Ͳ9,�G��7i�ȃMw�D��3�9kF/~Z��k�o��\��m���Y�V3)	T4��y��%V��+���~��z׌��Tu��j�wऌ�hū2)7���9�V���Ī�Q�]��ˡ'��s]κ<���Q�wqw�\*��Wȥ��I��0��EHB�n�ώ+� �>'�KJܨ^���3�p��Ĳ����%�n��1B-�ۈ����,� �6]3����$�de��ǅ�V*A�Cg'�a�깧j�Ku�4���-���c� �z�٢<U.y��O���5A8:B��F��ų��:\QD�a�1iZ�*vҧ�R0���4iI��71��n\ �<�\_$� ��JɔC^Y� �����5jQT��4Q���2H�cs`���Y�t�+�_�$��M��'M��:����Mf�8�`ybDbX�*�ߪ!�oh�i5��������3��@w@�)S"���qlP���-ͻap����ϊ�Gd����&���+Z2�	�J���r��qӮ�1F���+FF��7���O<yL��z���� 4�`���5X2f��B�5�%����bP5 �Ks���<�
��G��r��~׬ld��ê��2
��"�a�SS�Z~8���k�3����
Qum��|��ó9���x�l ws(���a0�R��.�ys],��r���*���ny�Ї�4 �r�,�Ǵ�z�a�+����Xe����)��2w�a;tJ�����ca�B�e�e����U���vf^t�Ԫp���ҥ�fH������q�5�c+쒛���6/��O=d%е�hO��d&��I��ւý�4%���i�r �iS3�(�/٠ ��0Pa=�����)lyxu,��sVA)�j?L\l=9�wA�=���#�Gj��cDrk��,��4����c�@�=���*t[epQX�L]������ޑ���%�%3��	�Q�h���ט�3::�ßR�����ۋm� �t�M����qFk�_e0w*2]�)t�c^���]��[��� O�L��8��p���/ӡށdPyޘk2X<�����1[��j���` ]��#%�� ��&}`���!���J�S��xU]5nD��W1�*x�����j���y��3��_���{Ӡ�;�G����J���q��Ř�F�q^4�<�����I�l�u�[���N�g��{��$[�ݨ�q�g�N[�����t̟<�D��\��[`k�c��H����4J���*��U�9����D�k��Mŗ���K��m�=��a�Eis�Q�3E�$;�hH{�=Y��dl���뺍B:�"�/M��&�K�����O��5�Q�;NMs�G��p��V1	<��r�U�]�*�y&=>��׬��N��W=%A��w����宒�Ap&0g����}�\��c�9�J�Õ�q������-�^�"u�?� $�d�{<w�� �شn-�,?�]@�u�j�������i� \N�ON3{�۴���#S�챃=Rg%�D�|`&r����X��4Jmy�&o�Ees~�о�l<}�{}�S�V��o5_�wE+�	��O��|����O��(�"qc��?2q �����Ŝ%�D́����8I���.jC䯐M^��L^C�@w�kCO������C:���f�r£.���M��MOC�K�WWd�WČ\��%K`kѕ|t�P�'(a�*��S�I�a�Z�BYo�ɸ�m3�R��Bpg���5!�fl��!�hp�5��n�E:���f)��2KDw�mL�]���T�_�ca��3{c*�}s.OT�S�焓,��[u�@��(�Y:"��2�EBq0GJ���9��,��"����rG���9;��:���ܥ��b*Ll.�tI��B���V��sd��"�Q�Jx��̆��������,k�C��"�x�Ǻ���'����ۼ�ϯ$�X�3��=D*�h�	���hw�P�����E�=2�oD�������7�+:��n}ևQ�G��Fɋ������W}>��L�B�o�l�}���WA�7Ru9�`rm�;��yS��������.��/+��� m��VLs�_�����>��}���}�L�ȳH����w ��AkSZv=\�ܴ���F!y,��c�4��h����+�M�0,\�MH��1W�a'��3�|�W@f�b�Z��������/Y͔ܫ~����{F��U�g��:p�E,� =e����L:�q���az^��:��О����ȿ<�aAw��ó��-��q^�[�����="�_7TX$m�4q�	��s6I��>R��h���rU��z�U���c�=�*��C���i���C�S��SOU��Dl�rv���#�	aA���f*�qA�Q�o�.�\��:c*��J#T�M�1�&�D!�u�h0��8��2ޗSЬ�y�,E�`{��N�.d~A9�|�'7��2��F�o����:\z���CƑ$��AyKL�_��ޏ({���쪢687�G����)�3݋��0U����[*驣4�V�:gq� ��OS.��
��m*�n�U�(��S:,*�����s��c0}o��F78#�ݒ����z�J�:�JC�.�<X�T�W��
8�'��5�f�օ��t�K�c�s�flp�l."h�?ꃛZ֌���c����:l��;~�d���?w��7Q��-�znq�m�4�q��p^�>F�[yA�xn'{�+B�K~�#'TkA%
E��o-�ty8�u����}��Qh_�z�<�r���<A'n.ѻ!Nr*AŚ;·ip�!tq�w�i6�9K�c�k��L�~�+#В^��y�ΐ��w��Ƀ�WyB���ߎf��V�B���ymGI�6���FG��W<F����f+I��������" ~L�ϓ|��r].n��e�<zW����MXt�ۥV���kLG��0H��u����M�ݐ�ǵ�"�ˎ��c5^�剎99�,߰K"�c��ͮ�TX(d�o
,��;sL4���,8 �� �HS�O~YGCQk�_�e/<4���@�b� ����k�~����۵p�nj�O~�����~��!���9*�A������)P�_�{����
���K	j�y��ֈ��nO~�c��Ag����r�������	ː�N*��.��*�I..���OϬ���+<(������KUWN��ȃ%0��OAhϿj�L;C��d0�y�o�7ҹ;��*�>G��}��.��m����%���t�AE6���]oK��ϟ�Lߗ���ZX�O ���#��=�n�����Iѫn�{�WS��a�iL�-��OKW>r������ڔ��F�[>�~���.HTS*��$�y�KHq�*z �o�5�〾��|@����kIfM�3D��Vi2	۸�R������ M�����ZR��P-{��xސ9R�R���H����V�p���}���8���'�땾�53�Gl�7^��X�`,�)��S�0���z$���vESHc�I��1w��
����ICi��Ϻͪj�/}�I
B�Y}�F�TyT`u��U�LeJO7������9*Ĉ��O�.��+�}�c?h�p��� A��cm~̅�W3��o�}c�jt����J�ٛhj�I���l�{���P����3TuN�,�LD���S`��
!Y�Y�A#Ǵ	�(E�-U�b߾m{��0�D�Z���K�{�e�%^ c+0u/��t�m9�����F�x��f��q�j8N�_���1+�/j�N^�6�~����v���qb��~��/���0%:L�s��ңfS9ߖ�Q��Tٱ�K�L~����~�6�fb/1���E��w�����ѡG7�K�r����x��̭�5��R&1�޶�|��[Ʉh��AEY�����
k���Uc��*ފ.�Tt��=��'M��s,�e��3��HJuZ��E��t:bjdu��!�V�+:t�A,�Cǅ�畾��n�ϟc-Kd������w���c&�&^P��V"!�U�6�,�L u�@;%b�O���� ���0��HN>my8�R�]V��Mi*j�YA��yȭ�Y6Hd�}8��89�V��I�AÑ@C��4k���"4��#!��<f���z%��s�`ҝs�����n �0R��=�\��d�sn�J�a6�]?%�>ka��]7� �w!�C0�f2��V�v�7 �����}�W,�c�D2�͖��Ш��Y�����u`nI��z�(��R{�i&��?C^�\���eA;�_����_{���i
�h�2��~���*CMjǤ��+ù>$�dN>�[�p?�s�A0rm	�0^H�E�eM�W.{��GUi������P��`g�h����R�B(�${Ƨ[�W�����レ$<�֮�>�1�9{}@W��St��3���jN&��*k�������s6��
Wj�dpi]RU�%��x�vB��j���f2�(3(���Ɏ�Yp��MtzG�l�7d�i�uװ!�~Q��C��'H�ptr�s��OD/������Ϥz�Rٙ��~'E�zЀ9?�	'.Y�\l������6a�����\ֺ�]�)��s	z�{��c��RP-��P{$#!]؁���Q+�u;Hc+��j�orsě�%E���H)քU�F)B������j�G �3e���Lr[�;�S���}��;ٸ ̎^[(B�M5�9�Z/�s��7Z]n�w�zf������@�!��I� T~�(<㖖��kDo<?yd̥}E�����<����n��S=b�|
�ɰj5pd��%rb��F�� W��?k??�'(�S=���5���<ND�
���l_�9��:S����Q�S�����5/Я�ܥ7tI�(��~"�g+2�WB��qل�tm2֥��:�O���#e�Yn�?�,�J�ƾ'����]��K
汏 ˄��=�Wϖj��Ě���ʞ�� ����%��l?L�4��Z�V����٪��jd�
_�Y���O}�^B��]0���rF���]Is s���[p5Qsq"F����Ϯ��������m�����^y��4
�A�o��$�,���,�+����8ԡe@:�@&f�i	Kz���xD�4s�#���=��L�z���^α��X�tA�ĖZ!A퀑���vF��a��u�fU�7��8���*wf6.��_��x�h��R�C�9W)�&ʓ����C-P�b����ã������,Gpa��YEm�	'��Z��~���Q�'�0h�[��.��Eϣ��Z�7w��r�'K��sޤ�y���"��83Gk*����<�PEjY����ަJ�ﳥ�c���R{�P\y�&L�ި�G��1�(��Z!'�8��E�� �XnO;`������o�� {" �x�΋3�F�)��u�E��Ւ�Z�.�Հ�
���_�h�ե�
�g�v��\U�!zF�(��UQ&�� ��^�������.��#�}�jK�uf_9F12���]y��
-T�A�*<B�O��4���+׹�\��"w����	�������EG��ʘ�ڽC�����o^����!�KmgEMV�@\��ټ!λ�vʽk����?�c!RTugTO�������"��5�P�J{b���d"��=�a�mb}�C	������ћ}�`UtN���$���ec :�H;YT&�N|�mn�?��@#�c|#-�S��Q�-�]��{k�
�:���k�|=[�F�F.T�W�bm�?ճ�UK�L':���08M�ӣX�	���Q��Q<�S���M��v�"Q�GO�/U��ռ�9��K�!�GX�l
P�H��+G����z���l���~?��GrfF�'X#�F�j��OHr 'f,���vy������]B�d,	z|G�/�N����`Hb�HG���J��U�Y��{{��w@Zx�#�,H�:�<�̵F � �����k���bB�a�)���\ԣͬ-k��K�#X��虯�������5��r͹d��.��T�V�;o6�f@��WF@'�](O�o�/�KH%V�x�^�(��u�+�+U�*AO�;���m�U��'AS��dp2{u�=I|��O(��M�{ә��r8x/.�Gb��l3�4�Gr�݅ :����"���u�G�P�/g����n,:�GM��G�w)��z�2vY* ����Dp--C�!�W��ԫ�s�EGn� S�3E� Oڬ�?	<Wy��p).�!^9������mf�Xy��l'���叄^�������Ev����mn*��"�L/��>���ԃ��u)+�c;�7Yd:�$���i500t� XR3X�ķ\śx�g���e��,�5r �ŇZ���ah�c�G�+�%�k�����Ws!�Ic=y��FT�bɬ��))4��M�h�x�z=���Yw~�U���(����?�_nO-���t���GH3qDm��q�Z>"�QC����H8~�׵�Jm��*�[��Ib��,�����-��TTKM��3�^}I��d��7���rl*q�47Z��嫃��ͭ��c�H���e�S�`�o�>Fm���"������
+OJ���Tig��:Gw[C��ԪJK�d���?� UCy�憬�?����0;�����������&,��1&�r����

t�S����/jY(��~����۵��P�p^i�t.Kb���)�w�>�}-�e��j>C�nn�<�*������>x�R��Y�ET�1�?�A��`�F�iGk3[�p�]eF��|I�sb�C����LX�9}m���Ty�_�)s��TXy��L��ML�N�o$�e�#'f��^:Ο;Гю���k��!��yW`qbx- )y%~n粹Q��Ӹ�f��SGK�ןxR"������Ӑ��B�l������Y��%���)J#f��)w��r����A�)�w�*�OR�%+auĥ����96����Ǝ�����op�a�Dto	(��*���>r�=u�Npr��	�<��e�(�!ڌaS�A�n�U�Yy�G:�֑�DsK��SLIa�s}&��CmI��_%E������H_T�ՃnTReL��/���Z[;�� ���;�t��g�0���Dp���^�'s�m��N�(շ]���"2�0}�k�2�h����[Н�9����#J!ނ�]!���C��x�S0kG,���#�fwƜ{�v�v��_J �&F��+TxSC�b�0����c�N������5�Q² �Mף�ĉw��z�K�	���G�pĬb[���O/�L3ޘV�e�q�	i�Ou�i�<� <}��߬�Z�X�����U@jn<�jhQ;Y�4�T��p��cd�x����ٝ�  �C)�/����y��~��Jf7H}�U���*ޅ7�H�M}���.��l�}ݭ���8<L��.��n��G.�9���-�9���gs�ѝ�l�:��f�e,<��д�C�Q����crY�ƨ�r�"���
CV�����x���N�Ǳ$�S��F��8C���)���u�������Aޕ/ǹK?�Su*`�����dh�f=��
@Ri�x$��v��|z�;�r5�S���Ӱ(<*n�é.lY�R,!�P�6�Q4l���S�!�|�z)a��j{{��E���p�ڐ1�n����6�ڱ��
�=�x �qm�]o�?��)WU=��1�"�"+��3K3/n��2�B��8s�F{D�дdg]�T�J�)�����}Âw��"\V>e�$�pN�?����{���W��S����wL��U�����������X�"��(��p/w��s[I>T��~� q�ĉ(���m�If�@����;�C���oj6KO��5����P�U ����VH4�*���D�ug"���K>@F%����"a�⼀�̏zBgЌ�`IBo���n ��<q�#x;��on�
�`�f���$��j�#"���N�$瘱Sɣ}onٿ�[����ǃ�gl��[�qm7����w��3�6����s3������a�V�}k)�f&H���R���U��dZ��$#	�e襦��_[h�H��/�����j�́�V�K�b�� 2����6����BM��d��LT5�� W���h��Ƣ�Hg&C�����n�Ɠ`ܸ|yǱmP�.橮;m^{t8�Pv-=�D���f�����Q+Z͸����<+#�Y/�y�u&�M?�Ri�/�2{YaRU&�w�y�$0��� =1&qrV�ض�FA\ ��X�Z��K,C^�R��Y����O/5����o�g�C d�H�[�鑻�NNf�w��� ��"|�F�'��R���K>�$yo���*�ۺ6�JeKn��m�k��Hx���ؽ��,A��˫�����L罹nv,vC�%j�g��f�moL��|��}Թ�},��OO#Q/ln�X6IC��#-����"���#,?ҕ��Y�8��s���Cl�{�e5_g��v�H� ����YM+������&��|�N�'�f/�(�aǔ��K[(��ℇsL$m�mL�`�4�;��k���o���w����z�h��i"��D��᚞R���'�h�� V=�<j�[Ýj.���B��w��ț����EY� "��5r���<�9ܓ?3��w�?IX��B��l�T�����d�����{�������H\za�%�b����8Ҟ%�"���JF�a���ђB�z
��Q�b�h���ffa)$��R^X��Q���p8�au ��������JK*�� =�|�%���Y����|�.$av@	�K��y�� C�Q��J��1b��մ7�*�HhCPǈ��f�.���$_ʥ/���2U���2�<ɞ���ϝ��G�#D��C%��Ѽ)P���S�Vد�@�w��i��KL�x��,e�~�q����*\K>oB�ap���p. �y֏�~��Q�h�<�_H�k�6�ъ�L�!u�U��)!j�7aVs����5*|gOO��Ԥ��:��OnُT�ɢ
cF+�8Z������;ԛ�T�]s��, Q��Q�0�����x�6���D��M��*��g�@���"�����gXd ��.����4�Y�=�h�E͓
��.��,�F����	����E�YGգe�(-֗�l�.��o2|�GXz�L�����l�Y��\�D����CM|��Ua�cY[`�l�(���-;��43'������/�t:��u}�O��W|m��"�y"��.���h}����<��n��sp��iĴ�'�P��u�ށRc���F7,ݗKd�qD��c�0�+�H��[2@�Ⱚd� �X�>���!ϞUv��g�r5܀�������Ԙ�縯롶�8��帨����K�ruS�/���mFJ�G����.��I���g:Y��<�

�}yW &�|)��!��'�T�b�#�h�=q��j�UCj])u����2��(�Eю���X3��t�3kU�f�R� �I��J�jni�&��&C�
�o"T��7߻�CH=��5�F=nH 5S�2x�I�t�I6�{��nYJɍRx�F`Y�aCOi��;y���LY��a2�Ϩ�f>rH{]Q��䗣a��t}pDV��*�(�, \��`�[��l��/m��l2���=)_��X^�V�T9�DX�	l:�Qz5O� �8O��h�9���^)�#��Fp	�̹^5��39^�y�0�єQ�z?6]�{��5T��=J7��M����0�� )L �����ZS��$��`�t)Iֈ�uRI��:�G�iq�/C-[�������r�̷b��:�7�k���s�x��c�9�����f~]NB�D��d��N +�2Ǯ��hK��tҹ�8��ag�R��ЄxO7d��܄�~lz�ИڰH�k��4�Js*bT�"�4�� �}@A,��[��|�_���ƺp(�Ѽ�8k�0��ɜ=)�<�s`b͚�k�Y祫U���S�z�i����z�x/�|2}KZ�Z��<Z�P��1�p9c>Z��qK��"����6��L1lW�;c��ˢ�����ڑ�n���! &z�<�G�1 �9f��!{��|�$�t_�l_��Ғ� �:O��K?�Q�~	��]�[AMY�d�Y]2nbT��JzɨRH| �s��o�8����y�õW|	K���na�FzE��8�����]��n�/Kf3f=x��)�#�
�4���a��
v$~��54a�%��=��%��.�w
MA��j��G���䈥�!��_�]T 
1��CIA1�(�k(H^�$����ʤ��h1�f@B�/qAhuLqS�V\�L��Fx�P*}\�g��q�Ԋm���,��ݡ���(Z�\c�y�Q�3~����U�h�5�D)��_��G��A.��XL�J1�r��)�п��T�]�a�	�h���=߈C�ܛ����ж*1.�������Q�4�j�t�P�}Ǎ��I�#����qZ;�����?ο��F���87r�A�Jk��̢��91�� \IU�t�'J��8R�u�_ #���f "|�3/O�����(��|��%��H���n�UX��� ��YԔI5���c4��`Y�G�r��M0:~h3�f6���R��T�+�2��9#y�`�Y�@5a��{��3���x�mm�0O|�"ތ�����F7_G/!��4��R����Ra���Y��6\��m��5=�׆H$8�f�B7-�DMJ[xE�{W�[t��ʙLMĈdG=(8}�]VP,_��_uK���l���Y�裷����R�/X!7&J����EC�����{�Y�=n�1<�X��f9�F�z��Y����W_J�k$�)��5�Mn셡#���S�DCW�%�����m::ꑨg9Ʌ�Q}���4ф��v�{d��{M�8�5�;�74h2��Бֆ�5��3݅��P����+���k4���BwKFC��&���e��w���$�����c޳�2d����<�JDI�=U`��"�S"��IIX����ڍ2���߶�����PZ|w�T�Z���̆iN��ĥ���vcIA��pa���� �-��U�u��ι3��U'�]�J�v����/:��$� l�O�R���=�D�&Lt|�S����@C���Rhky$������2�4�쾧��atN������xX��H`z�n	�S�����=n�>^�i �+4���D�^�-6b[\&7�XB#TP\��
��8fN�4>ePju?.e$D���W���ua*��u|�s/wyO�����=�n0�D���`�˕2��������K��b��/��y���ȅuO�Pkb&L��,������j9ns"FK�Fe^��MAk�$���/��&��J��T�#�a9me�kJ�N��5�3x#����K�G����	^T��Y�_���*�X��!yv��*>�?A4-����<�V^�Zt=���|�&KT�Ջ.`�=٧�S�_�0�|g�}Q@5��ǥ�'r,Re�	(B��E���E������X�8��V_��ӳg6GI+��s�=J��>�P�\���\|�0�PS���(:��Sؠ�z*>�3恗����B�j��]N9��L�tܷs��(~��KoD��l-���Ju��$=����>�ؒO%͔��Y��=�I���vHp�{�p8�c���Ӻ[/�0�����4����ȕѷ�ޫٞO	��.�����Ƽ�l�����w`Ħa���<o���üP������_B?�߬åX.5�c�i�W��$9���$�?j���X��˥����J�|?c"8�6+q�A%m"� ?�汒�6vz��f���Oa��.s�J�F���p������A5�]��P�	��l%r2^v����rv��ի	)r��]�Nە��h�N7���H��=�N�D���K�.,���CdL��x��6iq����Ki��4��#h��
�Q����n���"��������Jqȝ��W��	2�K����/�E�}'�ۚbs˛2 �v�hWs&5��G�SK
6�*�K`�he�u �9Ǧ�n�q4i�U���E�PƷ����,w�,>��ILi�9��nN�&�{�����⻿�m����|⩴�h�L�o�t�١�u�5x �b���zfy���1	��U���ѡ��u�)�X�A���UXS�T��7�g9�rC�E�{v����f�
bk�޺q%�z��R��\��gC���l�.D��NJ��$�9��ڜ��3g�©�7��T(�~P,F�5{���#� �P'��8�6��4y!����U�N��i7Zlh�,��_=�I6�l/�y����|0��o!D�_�1������>=���}.��{�	�?$������x���ܵq�����L�����+��S�$�:����1g�zZ�ͤ?�\�(�̍,��_H�;}�,���d�R��d¨�p�eni��ky��='? %���8ON=+���Y��;�BK�)�l���h�B�-�٪���u��n�b���7��J���B��;����p�L�2^����T}�\GC|ʑ7���H��Tpu}{��9�`��/��%&���.���#f'm�`��%>��]����vG�q�EA���v8'=�:ǂEG�m�C��Q�f�����腒[�"[�e`mF�m�=y�2�E/��CTʽ����<�Ԧ<�t�,f���z�v�9.B1�t�%m�=����po��"�؅Dj$��
��_�����EUڽ���!�MՐA�0x���$Q�Ӈ�rF�(���z-}�0�ϒn��c�[
Q���V�mA����A�١�.�}+�fv��"�4���i�4�;%�����|�ӫ!_�t��~>���������`�;������Z0T��0��Q&c��h�]���^F��c/��/A����/�JJ|�"Æ���w��?U-&x*?��}�����~Cҧ���s�$c�Sz��F�׻���:W|�Q���VZ�dT��$P�%��<�ktV�W&�V $2m=�9��&�(+���B�� �aR�v�,�7C�x��R�G@��E3��9b��c(�j�����g���nu싸:� <c�uv�Ff6!�f*މ���/U��f͡}^����+W-�4�%��X�Xpo��]4�с�H��E/�5]a���9�[��Y#�Ϊ��ԅL_v�� qM��C�4Y䡱�����P_��@l��r7�1״�o5+E\�yV�c��g%2�6���V�H�}�7�S :��ԋ�?����{��U���2�;�Sƍ�a�[��Y�q�K�X� �eqƟ�$�@�|�	�@��}�`�+$1A#�5s��9��qw���	C���������E���E}�g;�\��TY����`��E��uL>e�mS���vP��xaL�</e�
5�S�G#��mq�ÿ�p���un�<PKp�ba��ڎ^�舆�������=t-$D�M���O������9��aF��G�������8҆��꿲N����ۯ��dQ����R�-ܔ����.>YZ��q���d�2���V�<-��áa���u��@0~YR�6'��h�  z@ziWW�kLXK�w�&,���^���{$�E��~L#p��,����� ���G7E+��
�����1�o�*��bنwt��d�`O���9���7�v�^�E*�`����ʱ�%�zvrk���1c����m �v���SR�6C9T*�{�bܣ�er~����z�YH�9�4�!�Z�	{7����3N����p�e?��>���u#�˖3m��p��	F�� uq����Yr-@Bz�H"7��eo�Rvl~5�K��Y����9ƾ�2��B��iJ�y(�q3=@�%f��h"��D����x=-B��t
��O2�}���	�d�*M�= Ú��%��s$���J�h{+�n��H�R�|��OM�z�L��541p�#�x�s�RdD-�O��;ϠGX(�h�:K�y�Fo�͔�Э�^����O3R'?_�Fױ_�G�f~;�,������W� ���y$Za=SU�!I(��H�p����a�w `�oO��Ҭi����|Y������0d�_(zO����"����?l��ˊ�h�t���� �����y��A����~-WW����cIK۝�q�v�F�fؒA�P�����]k���K��F;���-������R�2#��cS��܉!7��׀H�"ӆ��Ɛ݆�r#��2��Ae�:_ڲ[�����]�n�s�O��y��v��{]�Ԟ�0TkHHOn!�߲�8" �
�j�@���?��=J$� �W�ю�2��_N��hN�p_��{6�[�+(ȀC�M��ފ��������ˆ�d�rb(�L&f��a�9��
�`�>����e��ލsAKu[��
a�}鳧e�Az��2�p�� ?�����dжB��*j��ŜQd_�k�(���Eb��",����X��bʑJO£��Y��o��IIi��"j5�
��c�E��-��S��q1�Y��VK��C�����'^3�ns~Ta�~&���'iqT�W	��Y���ǖ&ѡ�2�s
1��@Lǁ�*(ñ����8����2{�ȄWN6�k �H���H�m9�D�rqf�ޮo7�=��VNT��{�N�P,��mv>Y�����ę����qeٗ�!�4�WыY�(�q��$8wǅgkN=�"I���Se�	�V�4?����E��j Tħ.������R�T�z�BI��l4��`�iq�8ɸ��F�j�J ˪b!�L�S�1_frF�$0����m��qݖ�����:
8���m3�b�qd^q��V�Gђ��3�_�,_~�\����Rr$��.WR[I�(y����ԡz��Ս�d�X1�Ս�¦0��"��*�7ۧ�Ї��2�%��6��P0x.�zqC��@D���ჰdS���������"g?w ���Z8��|ؘ�C���D�9�iCL��*}�>}`.��g�9�v�븁��/B�g	��]Q�PKv۠t�:��g!ٯ�GG�P�?	�z���4*��ciP��Hs1"Z]���$�KJ�uC��b�}cs��D'�(ƽ�j��z:�4d� ^��J�w���8�B]��#�GX���%3��G�e�mO��:����L����p)W9oP������͞cC�/E���rU�	v|���ܾb ��Gf8`��Q��Ⱥ���y�
ebC���.6��P�,�ԥT����?����ËM��T�̃V
�Г�I+e���0G�'",CR���A�o���1se��=���h�����*�IyR�}�H��)N�P�O;��__k%}�x�l��D���VӦ|6�;@�JH݀nPM�XG�p(h^i7�E1��R����	��(*M��~�D��&��/�S ��*"Er�3��q�m��i�� �IwC�m�c{ЈvJ�m�	��vƇtH�ĭ���4��T
��*uY����k������=��@i��Rs�2�n �S'��({{�klu��l
*ӏ;#,�}��W)j5����C#�<��_!��S�E#밃x�{T� %]�k�~W"
.�Y�2B}��An�K��*'�31�z=(L
&�KR��e+��Z|߸�oG��\���/	S�=�YƟ����B�b�|� ��}A����¾���,	�$�6e���sv��߀bIx&nt�]η*v�Wx!9���j�t���L!R��^<����<{#%/�ZЯk�{���O�g�qX�q9�k/Ѣp
�`�\����d�r"���q�_A+.�:�V�l?�R)"�1{ݦ0{:Hd$�����/��r�#��7���~:�s�Z�e���;k9�3@WEyͬ�RZX�L!��@��Y(�@���#�l��x���Mm^)s{��ƌ��n1�2�@�g�l��/����㼾h���-e6��0�L_QH\f������?�04��R�OL��I�䇭J>�)C�N�1B�۝S�[��s5��{�zY�b��|bk��M/�a�97n�gR��N+/g��Z�Ə��S"�ɿP�*s^7zʖ[Œ���+R�����E��A��U����j$�,z)�$Q�J���혙�5hBJ�e������H�x��+^�cCC$�?	���R�%�#��*�p�I��ǧA4Fg��@�}j�8s-�.M'�^e�)�%V�;��sKX�΢x�+�Ge���fh�)��DZ�?W��P�7��ϗ�AM�b�L�`"�vF a$���۵�.��hD����To2c��Su�!��E��{�i�6���1��WM�pvG��B2��J����{��?m�.�hc2?y,�LM�R�\z39���Igb����Ũ\�����ʐ_Ny��#�t�ŪzRA�%aC��K��� 	���S��x���2�>$_��k�	|8�%#C�Fa�]��S5��e��&���;T���;�X_��"_o7�H�m��^)�W�8�Ɯ'��|�v���Ң�j�3�� ,�[��ns�+FU�{d�$Ѓ�Bs�vվ�VF��d�Z����nZ������$�N]������?`���nRSGY�bq�~ن�uWn[�(Zmy��{���R}�׻a���)��/�5J�U� ����O���5|^��m��rm L~khJ��Gm�Z��	U���D��{Ď���O�[�0��רKtL܈cX��N�%��[[T��E(C_l��HY��#���򕏛�eG3��g���m�܀���Eb@>W���B�g�����1(�)����2d�"����4�����绉ԚĤ���T����ȝQ��q�V/��{BW3~ue(*g�+e�t���Γ�󨽴	?�E{�e��R�qE�hJ���p0��X0p$Jt�Gpj9�OV��,I�S�"�=�a���-a���5�)b�R��+,ˬ1K�*��O�^��c�l.<dy�ↇ�ᚡ�I�Oq�A�Ƨt&�.�qX�T�a�FiЮ�d��t�E�B�Ζ���\ҙ����`TDT��[�}�ª �Ew���6ms����9��K�*`�"ؙ޹_�1\ �c�TMIj&��w�;M.9�Ą�3p�������V*����
p��>n��&� }�?�Qp�ܞL����Ѣ,φD��C����&�ksG��T��l�I�ݛb7�>�E%���Y'���"�2�[�}�-l�Vùįy�3Ww%�9+1�A�p���T���<��A~�ģvc3\(�.���rx���L걃6�\�ާ�=&dl>u�,Z?sN�L��5�T� �k�Q8��������Jm�QӅ� �vyl�e!���G�fe�d��pЖ6N�P)r�%Hn��b�؛�J�@w�+�e��j�=|����n�Z-��'���������᜶k�k�0H>xn��X�m1��^�^&qΜ��x���`�A$>.�<3?�S��W���+���a뿎�ftH~�\
�Z$s����댷�����q+�s0�<�;A~7�k�Tz>�&�c�o����$�HS5,Z{��`RX������ $%��|KC��oЀn�{x��L���\����C��P��l����dz�ׁ��)�����%��$��O����	��͔h�ݽ�z���'h�'\�Β)W�Üح�&�(F���2��'�W+�`Nb�˭
t������l�HI�rb�����E�c���^��-@���ux���<�1�@c�w��sU�$��N_�|�GAC'ޚ��sh��C�����:�����pd����O%}�q�}^ 
;��D������������; \�s $�or�$X��u]��������+Z��v.��v,��G0J& ��!�1��yRq��14�Y�q��k��@�����C�Hb��Z�Kn��j��]���K ��λ�I��mZ���6޵`�H��?�c~�&{�VG{�cl-NPַ^��c
�;֑��̊�#g4�5�>+Xm�t�t�b ��}�]���4C�v�-�|���U�)pH�e)�Ȭ�"�L�i��p�zm�&�"�'���M�LT��&t�R14gἌ�������:H����1.�2��x&�z�۾V��̴�y���qT�1�=#T�ex��׼/)� �L\CzTJfހ��j��W�]\g�V�P�؉\T��e�F7Ă��3&�V�ݒ�z��������H�g�� �(���t8QH�ĚB�h��s�������֎���)hϝ�N��l-]jQ6k��fͱ�7�xȕ.   50
e���+��$��k8 t��T0~{�A��_+�-�sdu~��f^e
6���#3�Gvlg��Ƴ����B���|��p+���!e�b���y&[-���ӕҔ�`ol굤K�3E�qOu�ȳC��-���.盇!�V�zB'�Cg��6����ϖ�4&���M��Ş��'�8�»���A���
�/�����L��9>U��s�Ԣ������L��w�=��ʶBsq��g�!��R�7��힦o��8�1����ȳ<E�V#��߲�̆Xc��}*����2YG���F1 �����:$ �=���Dw�����l%~5�c<F��� a��(dW�*������no+���M�BON2���ս�D
�*��oI���t�Z��_���:�+��@�H��%k��A*�eJ��dxhq�=@�oƷ6��: Xծ�q�W��%��*���&w;b�v��w��
-%���r  Q��Hs�u�8^N�0CF�<ϊ"�lA��U,`���>Dm/��F�L	���ah����d�����߮#R�ha2˽�zv����ۡ�γ������7 [�9��4ݜ�~=�����wH�W��Q�+5j�9��c#��Ӏd4Kt~l�XN�A&����'�A��1�6AO6�7�:�y�� ]���&G�4i�u��Vj�Pw(�n�o2Gzp�-|M-��F\�&�,�����eZ�j�����~MygS�K��5�'�-bl9~��k��t�-���Qחbf�M+��6U$��b0�J<��^Վ��~�ͥߴW�YX �!��Kj+;�~��PQ�W	��:�>�����@����.��Ɓ��
Z̋r�_�	��/��0�7��G�?(�gPrѼ��H�����%[�[�f0�
��,��5��Q�
�B�h�����}�gJ�9��I}����AK��=�l==�Gp�Ϧ���h��ib�.M~z��BJ�~jG܃���K`�&�Ay��dPd�vf��>݄R�x����:��GɗI?a֗����W_�^h5#����8 X��׮���B/_��7�\�x���7Zb�|�9�
HH�ڧ>�
�/�P4�������U��E�a�S�Eg0ݼ�%����YN�i��
� ��y`�0�Z�`E_���#���C����&cm� ~<\p�ʇ���k�9��ox��N� ��Y��uU����jP��D�P��'���8�եBW��K��̭�P�'�^ڙq�����1���Y=e��e��d��9����%��tz��I �~�����̬�rr�:H���'|y_�g��/,W	�+z�,���2���\?�I�Q;��y�Ԋ�M ʱs�nLz
�8�����:����#���1�1�}M�]$DP��㴃����0�s�E�P  #dczL0�2O8��ai�/m�/E��a���Iu�ď��v�JW|P��![`lJ�4�#����M4��IEP�՛K���'�Z@��[	��1^ �6��-�����F;a�_����Ȅ@٫J���y!�?H��)C� v1z&�3���T�"�)]}�s8Ӫ��oS:�'�1�*�%.PgASj*o$߇��.�E9 ;�z6[��-� (Y�Ta<k���'�KTG�B~�M�pv �S�b�9K�EZ�
���pL����v���.�t�]:-9�	cĨM�R��D���F 	&X�"��gVg�$i�om����f�	W�����2\�g�cu��I�t�ә_F��%p�6D}�"���/�����j���y�u��q3�qt���b���w�	�xd�d��b��\�6U�W4-�����yFɱ�H�!U%sXX���N���ƃ�[XR_��Lt/mr�`��ܚ��.;�%��i����#�@���E`�&_�U�:][�``����"$�9g�$��+rd!���FtCg��+A��0�H�Hy�oJ��AD�	�
�����G�`���4E�#V�TtGW(~��)�+����M/2���<�r�z�SA�1�q���2�2�h�dА�ȱ��N���!�w�9�|�wB�Dj�T�-�pr��e��9�,�伖�]�ơk�T�=�y�>{c��J�}"k�_�PQ(���{�r�۵W|�I��8h2AC���v@�P(�!Z%c����	�^=��c��,�ܨ����������_�#�:ip��پ�G��@���(3���e� �Xlq�j�m��K�G`�5�`��ۗZ�'�N��F3-��/B��tcSu���������A�r��g-Qj-֎� �c#��c��Z�����F��}�]J��L���
��԰۽Qy6�s�ց]��u�;���\����al�b�����h�/o��EN�["�@�{SPD��zmNA��Vȫ(3����S�N�:1+R26A��x���_b��p�DZP�X
�&�p&��F
{v""���4.EP�K�VqYk��Eej�ˀ��=�Z�?�ǔ{��Gc�6��4���wC2�q�8��1���Ɣ���ytYg>��C:s{�A���K�l�y}�w��>�c=Kb��T�K��Ԏr�HZ��V(����E�,P�T�J�ހ<�wdS�d�B.�x$!#�>|�N,��̐�jp=�[g�w��=�G2�Ʋ�yOǴntЕELo8M<�j��	���]o�>o�-H�y@8�H�J.ʚ�)���Ӈ\����P��m����iG*Gk�x;?9[du�t�áꦰw�k�0�[W����#�ꂘ���^�VYИM�'@���k�,����:?X�~�I�V�T��b�,r��t9|���b�L�^�������b������$U����غqA�oH���ceD ��z�����U>`&�o� �KCK�.��ӗY�]��| E��������W`�}[`9�5a7mA-���;6魖�o��Lrϋ匞X�Q�`�������@�����[�/m��t�>[�h�p�Np��	A�����ZZjK%�4� ��	կ�?v"���������Gl��P~[�@�_ç�&��È����0M�4%�<��NU���\P���H��
�j�4Ya�Ԡ|"��B�G��eG�~�B�X�r�l"ϻ�yu�;	�r��A	��3ÞJ��˛N�*(D������v�-t��yF�^֧*�'�t�q�5�� $Xj�i��DPC
W���nU�V1�x{��R�)��䎭��q��-�!?�-�!���Q��_�,Q��@|�ơ::�mc�9���e�5؂��O'��26�&wK�2�����N�+�~Ǎml�uW��k3���[��0�p�4�	��r69h�w��Y��@4@a(Vu�ٌG���w�@@�����pn� �}�*��Lְ�P� �f����4��l�ݷ�J�EAv�<��.
CF�n�;߱m�Qf�n���f�9��N̛)��]$IZ �� �L�PE��C�3�N��\��ǝv��8n�<���ٙ������7gQ\�B4���7l��R-W>^����F����V��|~�m�1�!�<\�X(�X�,-��V�2Mؕ�"]��@�o����ẕK���e�'�R)�2>�g�W����,�bN�K����z�\GAt���t��w��Vܜq�������p����,�� ����eP�5}��{�oX��`H��v�st*(��G"b}~�����C���������D�<�t_"k�gQw��C����X��S��ڧ|�8��%Aq�@+b��v�Ò�5u#�D��մ��AH��e��\�g���)�֘���W�ui�?�h�
H�h��S�:��M|�f�A�dBE�	�#5.�\!�	�b\SsǬ4}Z�$1����0/'7i�Ҩ�|��2�Q�aw�q�Iņ��r���P۹b1�O��u��"�u�=���[E������ղ4\(/��9CPO|��������F4�H�}gMV����d��?W�w�r�5%�ml��+�h4��>��P$��
��H!?��'��V���}I�V�
�~���7��e�iوs��ՄGR'�k��"x����`�W�6�I�4*�3�!���=�\	�yi�Ϳ��5��r81��n�jX�.�t�j<� l6�X�[�R �j3�Ed�&�%�{���J�>-7Yp0ci~���V��zΞG�v9��-� 7N2���2�X1��_����7nX���	6��mA���0�e8IB)SǄ�^ݒTt4��a��t�e{����k�eM2%N������xbP)��T(J^���LTQ3vG��)>v ���:ru��4��acG"ƀc>SF�mFh�Sz�I�uj�c�j+��2V�]�)V��dN6�����8 ���,��e �C%8s��:� _�t�v�Y���FM�0)!䅋����/�s�FF!�����z��~W7�Y"������7��`OߎU�m�����*�B�o?j2�dc���o�\tD�3��ht�$���]���R�;�"	�~�k�����H8�!�uMvm�R��m����6�o.CRlx|��uڄS��ot� W6�i��9�Ua1g���Tru���0�W#J>-($$����|(q�&�"OG7�C�ˊ3܆��3娮�<qF���s�&����9��z�cЄr�"�˰�R�Ϋ������p�}BP%�,=V��3�a���<��Z���� ��>a�R�s�|�c�nX���k�ч+�D]+�ÿ+V-w��^��H��8�RѽR(; ��k��Y ��w�t��/G�_8NO���L0W�Q)��ImLs'���؟��(q��r�]VF��M7����4^ۉP���!���}��E�dB�n���\�����T�JY:_>Cʑ	��3����pKO|^�]	g{m����o��7���'k��٨�Vn��X�}P:Y�	+d|��TM1����0D8�o��_�!�"g�_��͉�n��Vj�v�1���^�8$Ǐ� {˰�"Gp�K�O�,Ǉ��ĳ����VD�߶2B�\���s@�Z�`{���7��|��L�"=� ��W�����/��p%^Gٝ��9�ᗆ��N����h��ɰ�V�"�ˎ������-��|GkN�3���*^���5b ��W�,�zbG�c+�E��=h�ԂJ��"��O�g��rF~�Y3;㍝�!��V�hb�85��]EAz�>�,o�p��[n�`��vhǎ]����
$^�m{�\q�EpNƷ8�X�D��8�v���G)3�1s��a ߏ�L�ϣV��eF5 �XB�T���]i���9p(ӿ�C����"�]�9�d$���l�1�_�g�L��]�S-cG��ć%�q's_;���	a�q{��F��(�9)�z�U���HV����t��x��ʽ3�&�<3���Q�GC$��3]����-���%�S��k3B�P�2FT
ڊRaK����I�ͨ3hzo��{h�*���/��.�rG^z�&��M;�G�ePϡ���M�we����9�Ip)3e,(�ϙf�E�)x�dμ	�..��~N�>���\��R�~6LD�-qQ�k�G�q�;s�ƽ�wT#�V��xHp��Jav@ � �zm�`�Oi���:I���t�(JyXp��X��}���=���uM �]s�s��b���M��7/�Qa��w�[۷S�Z{�$��ց��Xl��>E\[7x���{�9�Gȼ�\(�A�>nE^�����CQ*�x�`=�4�z��$�8{�ɘL�Y�kmj n���{���}�!�\($ct8�F��ߊ,|�.���'�Eg�<U�ȱS��M���]Jt�	Ry�������a盬����.8VH�����/��:��X6�Z�xB��s��=�G����#��|��Y�.:ÉW<�0(��Y�V�S�N^�����Z�}_���5d3v����4Y"���Q��:Đ�z!��	���|��\�{Đq"��a�z���/��N��k�>:&�0���&P~�K�b��SO�������4w�hp�#��^��g�c���~�WJ4t.}e��p���&�g�=��x�P��^y��p_�R�V��w�$��8:���9|#�0�>l�z?擎��&���-ڿC�_���y�u_�,P9��}e�{��yr��ѝ�1|��S��br�(�#�G�?�I	��^���|��G��!�!�X+��z��}[g ����|���_تܶ��5e���T�?D?,�RL��.$����@�6�&c$>��8��(���LW��I^��x{�Z�+�+�@���xC�h��a��qE(ov���X������ݡ�N��V|������VU��D������KͷNZ$�yu�cɯ(Z �*��|��;	���ݪ*S�d�����?��_g4܉��h][ş������Gh/k@���H���z�}�֠<i��>lIt��,(�(&ߓ��/G�jj�B����FF���� ���*c1>�0�[A=�Q&�������X!&��n{�}c��7o�q�~K�O���ⶵ�*i�qё~c�oٸ&��WEt�o��+Wa��s���BB�;��W��X5�@0j�V�*�ƽC"��'A��îu=p&��A2Ր�Ko�)�y.���\�#�GNS��-M���U�W{p�K���ZH���)0�Ÿ�\A1�(S��� 1��,x���ngS���!���5~-5���!�X����%�R[f��r������w݁�ۧ����Z)H(�IY��"+�rj�O}��r�u�)	��p��k������<>l�=�<ڄ���:iG.�v0��w�^�B����x�Ԏp�@��4T4}��T<�y����FkP��	�7�r� ��g5�j���x����t�澬�\���Qn�^*1zJ���3�US�~E�r�������$��wG;��d"���,�� ��:�6���a[.4!�����h7;h�|�˺�!����p��g�O�����	'�f3a���;�<JD���m�ۭsz΅r��J��{X��MQ@v�apQwTg���E��~[��d�ÈUN^h��7j�R�:�v�v�a!
qe�V^}���C��t�S�@r�~�x��Sm��hY�'��n��O���G�����ў��z��1n���"�zJwd�$ҥA�f��H?�~����&�Y�Φ*�R�o��h��c��3"K����0{���ɼ�e;uj
FKeޝ�6	�80��`�M#�t��T��D��zw����y˟z�Mk��4~\m��T��f5~�)�y��h���Wԡv�e�W���}��q*�m�fyd��-��~�nm��{����DOJ��-��۱�
<�}y�W���X��B������w���F�ʹ��j�����!�Ѹ
~u��{��lg�Ǚg�@�w��%L�Y���TQ>�ˬ�'1��#��m��G�(�X�P��"���Iߜ�ϱ���\0�j�k2�?��Ѓ@F��!aV2dN�]z�ο��	��h�G���޶h9t��D�����ʬs#��Cx�DXxET5ƋY�Q9#��Vno��)���ک��_�����!�ɜA���?���V!(^ҏ�<��_��ȵ*�O��x투d( ��3U��v�ր.�ɑP��+�)j;D�C�� )zZ��w��|�v¬�*8���}ɬ�KZCq�l��"-���m��L�n�n��4���;H�h������w��Yyj���j�VRD��E��#��V͌<1Ql{�>�1:��6PXyŨd,��H�*C��|H ��/�4ؓ	ê��%�����+[I� s�b��85�n�l�0�ӹ`���H�0�e,e����c�Yy��̽��=�	/HX�ԯa&!nT6ɺ.|�]�菡y�S1H<�%\�yV�h����z�vX鄭�P"t��������B�qPR�;8�L2����80]��Im[Q2n���\N�f��p����t��b�c���� 3�QdB�q�ZP��34zL_S'�|��U᭔$����@^Q�����&�� ?���f$��|&�N���R�M�6����w������fl��1Yk��@����r�@��tmr�_�"ɰ�8�z�I�OnQ��G�#�?E��E�ݥ��A6z�皗��t�o��|�������f
���M�W#�| ��}��y�~+<V��4+��|�5�P\��伸Pq�`)@��U>��6���a.�+#�x��_���|
 {�헃C@�%:�ʹ��t<h�� =Е�BB@E�����Q��Y�;h�P7q)�U/��@�g]����F��ͅilS�we�V�t쟊z�e�+Q;��C���a���l��<�CV��+��#��C^���Y��T@�K+�ӧ�m��=�ZG�A؜q67Pw��t�F(�3s?��/�웙.T�j�e���ku�RsmE�/W�D宒�ԃ�Am�3-���퉺���؃..�Ԩ�O��+�����H�z�"m��C�2`i�\�+8�X�0�\7��,��
 u/.���3%�f^���>�Ɵ�$4"�FZ[��XY�2��������?��lu�پK��V�A˞LpK}'��xs������;8�HP�!��,�4�K ���/JΦa:�P�8zYv�;��v�Q�Rh��x��&�,�5��D����QZ�]qB�ͻcѬntab���t3+��f�'x�D4����+�q��H*%�2?"/���jm �<=0ėy ��8� LM�I-|�p&��L��%�@��OD�����$�5^�%;Ň�O_����n�E~ �/.�F�@QT�Ky�����K��e���-�a���o���?R�NԚH
MF*<���瞘���4�h�}�'Q%T!��~�^G��-�b_UR&J#�V�%QD�GN��a-bҬ�\1�nc%�^j�o4UMՇX����6@}�GAh�L�����/|�M�<�*G�Ȥ���XTߑ�۝�y���K�u�}��">�e�r���_��lA����h3�!�C���C��h���tP]jWI�,�=ݐ�du��������$~_���ji��\��W8� ��*N�~8	����.�W�$��)/ʛ[HA�I���<�13~n�����
�}i��F� {\���$.v�H��!��ua�b)�/����O�_��+�<�Z�gW�����bp愺��qjB�v��S��~~�
ۜ�����N��Y�+oO��\���S�n!��J��IHi$85f�OVi�V��pD�lɤ�]�9N�Q�� ���x(�!����p{�L�
��)˭-�}�l����ߏ�����Ģhm��;�/��f�灠Ԭ��]-���9�ez���J�=�����S|�aj��{ʸ���.�PȆ.���r�{�d��`��f��ۗ�يq�߷�/	�O*č��u�1���v�NIO�f�|j�!2��8��_�ҫ�r���s���o���=���F������H�w����F�<Ԡt�Ɉ��,�����۪<�[��.Ɩ;"�׻�s`:B�W�^�"�4�$#h{(�"�D{���۝�x� �T��~$�K�pALv����߆,o�HΦ��c���b�	!"d�E�8��V[�&�y��z�����;#�f�7�\d�-� ��'{�<mU�'�>�o|���6��a�U|�m�#봕�_ԡ]�2N}
�����P�-�p��_��J��y�i5�}�����<�9h��$���?�:�8�����fX�h��bJ܎�h�qS�[���;Uѡ���aߝY�;�ƹ���qɖ*[7s��m�'p<0'c:'�b;��9/�S_o�Y����@�k6��-������gP�6z� ��I�
��g�s�v	�Ҙ�[p�_�s�ٓ�����:|�����S��d�I�	���>vvt��S~���#��u�}�iK�1$��!����~c�4\t��?�f}��뺔�ً�������U���e?�+�������i�l�k��^[��C�U���X�#���+��~��2� fG::e�/ �%���	D<tM�ft�s��n��U�*s��=H��9˫9v�{j�VN�9�(:<��>�"T��v�'��-<��:�N��K�FKN1����,���#�@ƕ��3zeXBI��Z��sӴ���T����r���27��$���ϑ�Mce�KSbVk~VaYH�T)�pm�5g�7#�*�xo@� 3��":�91�EH@���o����>�s�Uh3��餮���hC�T.1�=�CN�&!��te;��4�a�7>I2�� ����վ��3�7�|J�6���msѤC�o�#��F�<��Pz$DG�{\<��O$�Sb�E]��%,�[���i=���;����q���n�?4�b�D˭d�%�F�o`!��N�YxR\����(�'~�^���n��myq`�F&�'����sw�d.{	a*�3��e���8=:0�#^�fG� 
gw���G�P��_��a���?��D�Z��>Nmi;�!��Ƈ:?��;��8X�.ᐒ��\\ �b�� M�:~��G9$"�+����=�#Dd�F�|楕�Y�LxB�S�ψEڼ��ڥ#��#7k1)�{;�`q1�Կ�z%%Ĳ�(h1����[�+?a_���kZ��X��[]�Vݏ�,����b筄���eh�hE�($y2�>sG������C߼U�I�+�@ŚL�f�C�>��L�Y��l��
�H����m�K�H☇��f��p�1Kq��	���H�`����ki�}�@��4�V�H���Y�g�܀�7]3�����g�I�A̘+]
N��&���C
d��c%�Q�9�^��CrʈT/��l�Y?.K���	�V;L���)��B1}�H۠t
8ftwv���a���Օ-�T��"�VL�����$�La�R���,Q���͛\��=��Q&����;Ʊby FDX @xn�	�2j�^���z�eVQ���f%!��<�tC/�~��	���w�Ƶ�����5��V2��g�v���p�+9��0�G�X/�Nψ���||&e^(��kD[5G8� U���R�T��Ȼ$<����X��F��I�:i����;��)�YU����mK*���c��DMog��hwĢ�}���pr@+��2݉�a#����XwW�+ͳ��F�Ȇ!]�j������w��95>�0�Z|� Ӡǣ��O��D�q-<D��%O��!ZQ`�p�Ǯ�ϳ�4���� ÿ�_/@DV��\�C��#G_�+xN�.d�=���� ��e�b�����{�5jƑڢ�N,l㇁��ģxI�a	H�#��9|��X	eS	2䢜ca����@y��+\�Q�"a�KaT��X�����Ƨ`��}�����^j2Uri7B|r�����߆�*��M�������n	K-C���B��"�������zV|-6k�ea!5�h�gO��ҡ�0��8��EƮ��h��µ�ߞo}&ȉY����q��+蛲r�����᠖JSL3���t�&�qej��U��5UAf�A1 J�á�&��e?ϙ�d:� R�uQ/�~�Z}������.��qS�8�uQ��M�����`Ϛ(�/��J��rT�{��[v�ҕ�K^���~Ն<}�/��/Mq���[��Z��n������� ����࿦��oJ����R��`��6�G�i�c�рf�[T��u?���|��!��GA� ���bC��������6�#6>$��E�[:�_	��n��Ty>�b�9W1�!q���ܞ�lfW��>(b�e*g�1R�L�^W8_��k�T@�?���Я�Z�+�U_�T�����XB�٨��tB��(��-�^�Vlw���g���h�eO�N�ߢؓO������C�Y���(� �+�Lk����Ӧw�p�7���ytI%��|(�c{4���u�1+*��v���P,�^ل��@�3a�6g�4��m�>,� ���(I;�xx���>ND�V#)t���Q���^g�+��<H8�oU�\m�	cA��uA��?jb�u��7�fm�S���$v������U�e+�X�jy��F�er'ް"��M2>@�V�1�s�}+��޶e�P�6y���D�s�����5����\p���ʄ�;S�Ӷys{~�M�ܶzP��v�x�T{X���-��Se@nZ_u���|��r�Q]�HoL_������z�=���m5�=����PEc�-�%w����ܳp�B�L3��ۨ��N���.�����E]=v�F�s4�\x�'��)���5�7��w1�v�3Yjb��5 X%��j��4cY�)W�< \�� Е��^T��͢��ӏ��i�IҾ�%2c�jO�4�g���h�������eH�Ƴ6Mт�.�d'�$�S�Ts��}���3(��t�0A�B��|�i���e������r�?�i�6:7��@���q�=�H֖��\p���q`TA��#X��2rЧ|��&�� ����,�@j���Yq[S�2k�.NV�E�ʊ�̹Hf����j�5���H{��'�2⚞x�#vZp"���n��C�"D����lCF"$�l�2����dD0�=,E7��Tb-�w�3�*��h<�UL�z0@¾<�u�|R��"���˗؝��d�m�U.Vh�Z��i$�#�Z>�S��3o)�ދ!�z���?�X�H�%�tE�����Ս�I��*8���6!�s��7�b��L����1�P�n}�}���IpD	�P��S�.����ό�W��Jx6~�Q:� �fN�O5��579�ن+H|����-c�9�&����8��c1P��󇗙!�x���55�� � �0�,P��\�t{����n֮��P�b�CĔ�/��k�>bpFk��l�f�r���ѓ�ygR^��U����;������@���6FX��s��'5wuz����&�wo<a���u���p(g�h_W�B��q��O���7�wt^>U܃߸e[�niW9�W��w.� a;�u�wk�a}����]�ؾ�2e�^�O���/�:o�Y�u��:�}�ی�P�S�S
�\ߵU� �}]h�䰕b�8���pPl�k�kIOZ;�К�R�͸��G�7n�l[x�c�)�ݥ\�;����錠޴�x�)�-�:8�o����r�M4�J��GC�G�jhf9yGe�@��P��}QU#�.���R{�O�Y8�1%O�g��+�+ A
ެ�w]��3���3!��f��+�.��-)J�!~��H�1���~��n�l�Hg'�(Kշ.>��вN��������V���qKȐR�
�vҽ&㘕r� �ۍ��{�çh��>�(�5[[ȼ�-#ڣ�
�O�	���	��E��="鵧g�J*f������*�N�%���H��8X;7����ݑ���]�ß�$�jw�b��wRf���!V�<pW����g�����ZSk�:�n'}��%eteRb&�(ϗH�3\��c��q&�k��U|"O��W�i�+%Q���2�H����,O著e;/�:�\P��|��uı\3�y�q�h��邺��?#��#ri�m��vL�9��F�ԩ���J0)p��	yl��)�q֗��'��c�9�a-�-�y0��� g`Q�gw�<���Q��y`xN���p�$������9�L`���{�#���+Y����BL�k�ӂs���ea�./�Jp��ݷ�	:	�nט}3��3��G@#}�U��Ʉ�Sh2"5�V�p��q��0�owj��Z�?S�?�4��
ސ��Y��_�;�4�	�ƪ97xE�0LZ�����.�7�8�g��oM	Z+j�}�B�kͰ�ǺZ��+����}(d���A	�+�{S
����_T~�+��O��(�1�z�1�a�6oD��_ފ?<nොq%w���hqH3�e^�c�'(7��,�R����I�}x��ӻ(��A�] s��⢾�c�v�� P[I{6hy1G&��uFZ��;<kϸ�����`yn�ϝ��Zy��St@�����L
ژ��߄�?�l��S~����>5���~9�^����m�L\T�a2E��>�j� L��'9�y(��b��g��-��O���f�3�@/WR�pA�%��P�4���k�*ř��u��t���;7�\��%x]45����A<x~����;2-�s�Wv�/�O�69�-�&E8,nX�|���4�/�w�(���]��Т\qe.Y,+4�PNB�ļΙ
�u�
��i`�QS�<�����aߎ�49�Ojhp��{����t�ߩc������[?0��Ցyw�N�]:�@,� ݍv}^���Q�zm^�J\~���B��ҳy&�1AĀk��ݧ���ZoD�#���v���������:5�e��0�1Ɖ2H�R'$���^����>I���P��.�,�h��?�5�!��S]����5W��|�As��[<|9��Ha�\3�"4�n�5�C���EoZ��pm_9�D_���z5-i��:2��aLԄ��7p�؛�n�	h�G��M6����|:R�Tǌu�����7�5��S*q�.���ިj��W�Z�@�=��bH��@�c$=ͯ,���A��2�M�aD1�0���_.5"�-GGkǣ�_ř�����J�X>�>�D8͚� �9}�Ȧ;�2� �4�Wn����.�姼��$�V$��0������M�A�{̉&p��/l�R��N��#�	Κ��5�NL^���I��!)��W���'��#gз�M,d�5�h2������Ϧ:��������o�W��AI_�u�+�������wE]��Ȼg��u���Y"ZX���d����� u��F�qR�oL[sX�q�I�ѫ�面%j��O��]���#5(��-�2�O0� ���H�bC�΁	�g�t�g�v�E\���_��?���s��^}}�6*|��$��O�8;��O�3�\��Ch��R�Kڰ��;��i�s^�g���䪢r�*�Aj��q;s%�g�A%��e��Q*�p��T7�1K+q�3F3��%t�W͞��.,7_�Zlw~�v���	8e%O�i؞������9��8��r.:�����q����"�&;H��c�/�G��\�ݚɾԫul�t�FSi��*��:�{�B�0;럕�8���H>e%
*���q\`��Oq�N$��*̞�JO���r�����3?�)�n���h��V�'k�de����߿��|�5A��	C����RH�J�.�:��cZ]�vo
^��N� �c4�8���l�Dƻ�ńA�`)�Y�@��t2(5��J��)�Է���j��Z�0��dk��&�r���Fg�0��γ��*G�Esw���Pq"��$A�Vr<�6�Y�x�{m?�r�����l"��$��VJ�,6A*
!����0.9b�������Rzs����?,�@�k7��H-�2EH������P�&�m��'֟��ǽݦW(*�����-wŞ� �k�S$���L:���@2�~�#@���֢�eE,=R���5�/��1!��ګD�d�~r���{'��pG53�q�2>���i����x��&bWӻZ�>[q�<�`[�Z���"f�C�j�e���ț��g���(&ٹW �|���Ǽ!���UU^�xPQ�rt��Nx��T��l��K�."qb��z3_��@�A��D�VU��4���Ә,�_\t"uq���LB�"l�k@�Z�5�%���D��z�����L��G嫶��]�J�t��.X��F�n����l�$���J� C%�AS�?�=,;�SI�1��J��`��ҡ�RY��B$QRp����[����W\S���I�nL�"M7����?�#[=Fp�Ne�~�Z?�w
���X��G@:ˈƩl47�c���[� ������RB�!��o�x̌�J�ظ'�Bk2-4��f��s��F/-���Q�
�_2߭��]Ձ���2�a��/|5��(�@	�p�׹fk�e��
<8�2�����%F��vcwr�'�߄�߃	X����H��Q9�O�^��0Vˉ��<#5��::��eGj|�ʩ���Z��骁��#t���2[�UW7M�^"�K$0�1���p;�u�wnV��D��u�����}� �)��l5�b�э���6��E��Q>�D&�ib���>o���S�>�H
	��j�*��9��yw�ݰ�&I�Sř	��ݿlJ`�\���,j=�5W��:#k% 'X�v��8{)��Q�����*`U�j��l�r���)���T�U�r���cF��֘��.{;�~g�ME����7�=<��G�|�����1D:��i�zaf{�<L!sJ��?CӺ��#<�p@U� C��+�CPs�Ab��u��}% ���Ao���f��mSU��=0o![S����yl}�:�ht� Jd�Z1�)/�����bWv�+q01�:��ܩQ/Υ������,E��A﷌՚n��,�����l��>`"~����[�U-;$�X@�Yf�u�`Q�6������nQ�����yA�K\Ȉ�k]�_�FA5W�� RE�V �3xLI��W�8���@���˽N�^�Ƞi��2�bM�Q�2?�0G _tK���_�e@���̺`d�!��v�mݛ� �F�Ic�& <P���-4.�wN����)2�C��$
��-���r�Y@m���[	���k�V��?)��d����Y0|���jGmDI1SD΍�D0"np����+�?�Gbln$�惒�q|M�?��b��aV���ۤ��J�K��5Ro��\rK*`�����/����v�ȸV�-�&´>���4aD�f?v�	��$��	�}����c�*�
E1��>�a,9t��}�ס�2Di�E��VI~�2}q��Y���`�[+�|��2�ߍg�$
Y��s�����N��k�Ň��[���x��f&1x�;�_�F�X)��[`�C[9ef�4�F0�6L�i?���w�M�F>R�I�-T��uO��%Tƻ���y����J
�w4�y&��C0Ix���~8W�U�s��1�ܰ���b�`���w��XPu�c�Ŧ_C����̼�e��.\6�wVS8"Wy|�s��&`���	��+��#N��0:�O������,9�����<�����L�
��z�z.�䩎�PA�lV@���F+����_�R�q�@�5X�S踂]�����`sDe��=O�*~�n�OSu��o�2{�?i���@.v�Ǝ�6���2�qRc�J����2L.}d+�J��'oa	[����޳��UVa@�8j�&�c��HL�q
���D�����g.㖿݀���f1W-Zb��XPxIm��L�ե6_��'��qQDN�-�����r)��+�>~��SD�-�|�"rXAe����ʸ������}{dz���F&k/��,��ws��8��WZ���~��׌H�[������\�'!�	�	�oY	��U�{A�-��
�6@�O�`M�q!�c���Q��O��n�W�� �?����لj�7.���+�*Y|���0��~v�I��W<�05B�j��J,z��f
Gt��7�~1�3g�vq~��P?����VzKs�� /�	'�w�֒��KW�){�b:nQųHJF<���		�39ӓ�������������fq��|&����êyׄ�a�»�����vBG�P&��-J}��5��`FA1�'&@Y�̚�@}u-x��h��H�Z�i������,�������^�	9�%��e�� <�.6ᯄ���L\���$��koC�0�b��� �0d��f;�3��H�6�`����a��k�Aۋ�@��F)x|f��HЇo]�J�����f����Q�d�����3qK�� 3�z>����ε�)F
������y�k$��=�K9�C�!�`�����9��;�v��܆~o�͠w�x��dõ8kй���һ?�I�C�t��d���|�ڿ�y��ۜzy�$�����٩�gģ_|[�%�� â��I�`�f�@e c��|��iƞe�0��فJq�6Yn�ޝ#����፴$o�m��Z�`39%�O�$�^; �.[~�(-�ޝ\�g_�k�<�Tsb�� mO_w5������
��ڈ�5A�![�Z�y��M�!�.�81�MT�!Y.�܅�s�I�w����p,3�����v("-��6�P��k�H���8� r��4�$_��H�?�A��v'2�������B��E]��z��`�/D��ϛ�َ3KfY�M��4@T�=��?����g_R` ̀0��G�<�G��Zd���TC�|���M;�����ʷ��p�v��[���?��;�*�s�
�خ��tg��Eo5�/aЃt�>���,vX��锁�Ln��-�����#u�b��^����|y�|��z;��A�7R�����x0Vv-),������3��^�%��C��4B�@c��[�kh:����8��\䈽�+���Z�T
o�׷2�l?(~�x!��&�Q`�M2��"Y%F�o	�CG'x\��T��<�*s�?C�V��x���A3n4ה�*U�^�3(U�����
�%R4!�����{M��%��K	���7/�C�r�q�h��S��0ۙ&yr�mX�R�lA�|cK7I>S�\0��;���Rt�nO�c�R�aT�3�w��x���y��ß p�5gO;m6���?a���NꏂU4J�5�)WV��V��^�ři=��n��<V���U�#�P�qS.~�ju�lo`�c���<;Y@l7p��0�%�{!Wwx��b�J�#(q�O�nO���*�v�n��H�Eј��by��N�Kx��R\�����/�r!��2]v^��P�3�!�2i�	�s>9�S�B�h������1�M�?d��B��.��@�TL6t�=���k�3n�R�*����P�V\���sy}h�}�Y��UP����}�o����Dcp}[��Xt��0���5E��p�oO��:�	��YE�����ظݠ�`7k�=�(��P���bLs��^F��-�����j���p�{1�g����k�X�����NN��;�D�Q��Ґ~]�HFb���$}�T�kA���?;�r4̧> �J�"�W���V�ɉ��Q�<E۹.��N�	��iٹM���\�S��t��G��i�)\�Sɇ,�M5+)J�A-��U�`�*FF�w��I�8�Y/�<�ܾb��N���*�R���
��������r��h� *�zYF�}L����P�
�"� j5�T��49w*
��_C�0����>L�/�����
'ڒ&��+���c��	���&ʲ<��d�`f<[u���P�L�Lt�u�)es,>��"�5�Yy��Fß�@�~	Iݥ>s1���
nt�89�'�"��q�(��fM�Z���
*�*qő��|������D|�����ս��z ��d3��q���m�9$��ؼb6�3Rs93�
K/J+��jr������R�J������xI	��a�-��&e0�P�G��U��ߔ	"X\Q�����<b�m���w����FC��;]��1G��9o��EDXm�������l��z��XcBm>�;t����FGP��S�8.0����e��hR�%��?�F�s5'O�SO��u:/�WܷS�%�J�5C��R�ȇ��T0EYhV�_)W �\*y�+��W��a�+���}:��l�y���aPH@7ͻ(��,����	�UuFC�!��c�W|�v��ũr�
�f~S=V2�b���6up��Y>��,��i�#q��7>��`���&iõ�m����8E�� �������j�،��V(e,*�3���Rx�`��1�yN�W��cZ����h��\��N�=�j�F���[��;�KJM%�Y^Mc�2C�OWw�Ϫy0������В��r����J|.�.���Aok��;z��0���f�sE���U!�+Yn�4-�X��vǤ����Mg!��U9!Ax�WI�4눅�ˬ�l|��6sJ	�,)�_��;h	'��6W���2�;i�����
[< Ϥ�hN#-�Џ&��+���2�ΠY���`I�E�ޢ7+#^��v����E��5�PӜ&3VW�� ��&�������XL���AӠ��w[{c $&��L��8���\2E�[�?�z.K�g_�D���97 ,Zh�`l���G&a��T�t���nL�����$Y'�`[�祩�
�32I��f8�!��{�er�"]�&̍��*<�I>/���@��+r�����X��W������,%Tu ���G=h�@	@& =����aQ_j�^�§0i��ZPba�� ݟ�[�D���4����/��{:��8"!8�v@�����u�����޽K�s���)��ސ�q��Dj���u�oW�^r*�5��ǋ�!OU��7!Մ�F�w�dXzTT'?���#Q�������,�%�k����9(���_ک���]�͐��QC�J=�/�c2z>tY#�����s���0-��I����VέhA�t����>�+G2X����W��容�������jMې�r�ױ�S���?�8�z��_9d��F޳�&��3#�)N�+��8��u�lsO��5Z�e�b�vz~&��j���J�G�w6 ֻZt��h��<��o����B3vp�M��s%aΏ��)����-$�VmOO�k-��QW��a����0N�Y��S7LV�h�ʞSR����*|F�.࡚)�D&�

��%j���~�
D�ZRv�N���Y��L3�����ő���� ��j9e��u�kwQ,�-)A��5{�\>����8��F�Tl�%N%³E�W��ӿ�����i��'�P���n��[(�3����\�پ�@-���]��33R"M�H9�U/��2�ċ���F�
9&��d�`p&5�����v�d�ю_۝,xn�<<�Z�����%��0t�|��7?�ܿ�gR>~��54�Q�[���5 �+��9xZi�L�����zâ ��U���)��\�*>����Z�&H�v�q
�����)�^bP{���U���d���]�T�����a�d�q%L�Jjw0�_A	�g��"�-����*�Vh롩���@��4��� �Iz:�cL8�S,�i/� ���7���v<X|P;�i���dI�c-�h�/>�xJ�{F��Ǭj�@~�Ѭ�M�ok�52=c�/���t����w��	Si��_�`�6�#�5�e���t�AS=�3M!���m|� ~�7����/�:R�X���]��$oX*��������rG���{ĕ7Z%�m�`1qU�4꠻��pr�I���w��Wn�^�R-�(�z��v_ �R@��,��f��+���dف"� ��w����=��kЦ͙������P3�Z�DRZ�\]�mǼ��:v&�e��[|������鲀�kI��#�u ��B(\fg����F�jWF�[ɟ)�҄`�V������|�媵B0U�C�+���fkss��fB����9����3����2��~�;q�r~�V�8���%�E��?Gvx�n�u@��g�]T�6d+L��"��+6/�m�u��-`�f$ 0�pS��aJb��%�9��LѤOs�E�ܸ�$��a	��c�%��x)�~r\m��<�a�t^����uv�]���j��.\E^v�N�����8�| 5�#g���B<ʤ,ˉ������m�ܚ�dn�i����`�;�'t	",�q*�!ɫ6 �&b�&��SW2(^���s��z�>��8��D��m�8�N��9���aC�)?���=?xg5���Z��^[���#��Ki�4]�aV�47�d��9�_7�����P�7ԍ=DQ�F�@-|�3\�%?$:���ӽj���DwilA����}� E��Ks�=r�� |̌Us���y���|����og��wΆMPʱ}�t�ow�B"<r���g�I�|�h7$����zӲ���49o�W�'�	��Lf;?�01?02�޿ֆσ�D*!��o*Pz�A�*�:h®�j��J;mg��0��^"��Y���b����*+�I��
�:�3P�T�,O� ����������G,rD`����-	T��K�=늝B�� i�P�Zk����(�[+�f�@�[I\
Y��v[3�c�}��l'��"ȓ����W��hL��̠02\�ۉ�X#�"�������lzh[	��U���[���A�	o��k�J�
H���rJn��� �R������x���^���.!���=��1�6W���v���\RYgT탛+��r-=�
2�P�KѸ	f9�s�j}A�q�W�
�	u��bg�˴7/���1pϊ�R��yF!�T"����9����+B1w�x�������J|NQ�����U��GǑv�.��5 �3^�#q����Δ��Q���#��B��&���<�S2��n'���y�n�,x�v������̪���\b�z��Y�8���7�lOY���t�*x3���+��?J��w2+�dj\R ��ZT9ؕ���-߱Nar|ں����eK{y)�����pvv-��u�d��s�S]�.��->9�H8\�.�L3��S��Up�X��w^d�#�=�/h�i�n\�x�J��CWJ��!�0���e�S��b*� e>�<C�2h�����k���`4jkW���j�7$m�\zP�RA��`<����tU ���8`!�9�O�M���+��6�B�)�M�_���˛h�ny�ȳO���"#�#�\�p�+��]��a�w��C��R-��mh��gС�6����(���I�0r'���➼)Nm��7x�|��݊�kȌ�tL��O����d3ih��Pmt�x_�Gi���m�_��%�ׁ�֧�x*P$�RT����x�Mj]GS*Ӄ�^R�!��{y�������e���ߗ�Z 0��e�Nf�`o�a��7� ՉkWȌlŴA�4�m
�s!O4���yFJ�1����H��믌��IJ�T22Cp�H{��８���VU.���bڛ�,д`��b��[PW-?߱s�)��m,�ȕ��>C*BM�#d�!d�u�p��?`ތ�28��yU�Ӕ]T�
�W �� Ú�\���H(��!�6����0�5E�:a�˶S��N^��>��n�M�A����{n��.�Nm��d�-jIq{[S�=]�4H_�E��ƮĪB���b�5S]�1��
��VeU������yJ�Y�	k�R��?�n�Mmb�����֥`|f��?^���4D�Ŀ��.�K��)]�ohͫ�\%[��O]�m�zT��]�(K׼1]b����=ZT.w�"��,>�$��R�c q	�r�F��\�BY�X[�\O5*�7RȨMy(46�\��?/8uGo��h'0Yr�q-=!�߳ EDN��r�g%��)�M�`�[���H[!�OHP,��[�i�u���x�ze�fJnSU���8�d�����!�xE��+O�;C4L�5t����zOh�	����|Z��NZ��N�N"Tr<�,Lӽ��w�#�e��<��V�K��z��ֺ�V��]h\�e�d?�p��k��<��(��|7��G����T��n�򙸧�I�T�q�$=��ގv�~y�s����\�I��t.��f���JW��rjf���<�@
g�}����ױ�Z��	x���f�pf��S�'�c�y]�^��8ʪO%����ê �T�fCBt�`2����|}�d����m���� � `y��4���������Q�M�J��� 	+$�"�}��B��׈�n�V�JRނ����$�,c���Kv�?
���c��̊���n*�rANU$���Y�V�}��+�.��G���f=�>�jX~�	�@�Q���J���D������]x�ZNo���υ�������|�h+����[X���oH	Jw��h���mLT1Z%N�i�]��/�3��#��֡m�.$���u-���Ck�7!���Z|��Ae3�
9��{����j�hz�b����j����h[�����o4��>5����� �K�(�9:3\PA[J~�#C�q	a1�L����W��4�Xv�5�����dT}��
{�u�(/Œ������?
�����Z�dE��ќ/�<ۆ�犆��}�	zzm:?.��s3}��pB�1�^�P���A��y4~ԗ�%�_;�/�n6搱���wz9/��B��"���3�X�Ex��),�)�2�bL~7EVM���>1'� s�e=���G�!�2�k���u�	�7$}E����]�4Ƥ�y�ᕇ��@���C@XW�[��[j��&�,��%G���N�����d7x�%^DI��1�A�� ��ͧQl�%m�l,gɭ���\I���/N�H�@
�x -qB�O6��
�q�w}�|f����h%I����iU��'��(�����m�=
�6�`#���~��� �@;=��y�n��Cm/�[���dc��s��T�xÀU��K;�ok�+tk�ÛY4f�̱�?��μIRP.�-��c7$��IH��	1ݮ�q37�O5d5��h\�`�XR-O��wK-�P|-��F���*�k���PDC�;R(ϴ�%M8���Eb8h�`eԕҁ��o�  �&Aմqi!��誗�J��o����� ���{��dr��a�6]�.��{�wO�0��G&����v~���i=�8��I�{����Ƙ޽͈�-��;�g_�9�XQ>�g,�[H�	!�=���J5��b����g�8�#���Io9ax�����s6���_���i�K�I-*)?��d0��of�	Z�@��w������ˉ\5m�2.�57c��fNN5"&�n�O��r��Z{�)w�ir�{�TdG��5�߷���s�&We��>�R�E�X�6O�eQvV�`U�~~Ŧ�h�0�5�Hw���t�a>ﱨ4��|�z�Dm9�55�)���{G�(����^[o㷷X��	�� �q-R���.n�a�ؘH�m%|���T�d�:%��,��`a�g�2��|��mD"F��,s����tr`��J���2��j?���˄����sJ\v�����0�2&N�h��R됹�P������\z^R&�X&	���d-ȩ����D)LF���=�[$�EE]&��@/���EFٹ̍�l�d�.���A��k":R��Hg�2�J���8T|�q��~��	H!�0�Qx1��Jl�i�tAx�������N���H��<<g���Ԕ��3��c�BE��֋1���m�|���'][�����N�C���@e��
~4��'G��1�n��󵛦8����p��P]J<�茵R���a�9���� �Z1����6�W7���a:=B�r�W���=��
/,Q�����.K)�c�"�0�MRʟ�E�Njh&==1=���w-�����x�>DJ���=�rԔs��'�a�*t#;<E<�� �ʒu�"ޥʖ�n�p������P1˩82D!�5�E\1����ڽ�e
�c�#}L�YV�2��x�?��rPP�%�\1������*�Sw�K��1��l9�@���0ρ��j����ۺQ[;������9�j�ܦ^~a��$ό�7o|�w�e��YY6��w��;�Q��j��JL�Z.�o�Blu��(_��Tb%I@��%�7T'�r]nҘ�E���lg[����9ǹ�'�
�3�Y�>����>p��9�&CЋL�OlĔD����e訋�E.V:�C�"�=��wz1+�$�K���`�@�i�����rV�D�M���J���t� WI���(l�ugI:�E6|��'�<�䬋a��I��/���L�]�SX�#i��*m�� E��|ޥ�(�+�1����ҷJ$�o\,u����r��$�l��<G+c'�:$À��ي7�.�x=�͉��r�I{�H���EJ/����܄����z�@����#`�dRu��XN�<	���2�~M��}��.��"�&��S����B���%�-�忘X_�^�DR+%�.�jh��K����~��Șv�j�͌ާ bob�Á?����j���s�]�4��)�/� T~�U��٨�����O�4�VV���ι�X�l����.>������P>�S҆Bt���7[F��]�sI��7T-?5�j�[��e��1��Q{B�,�T&S?�����r��Lݓ�[x�B»��2)�����B0�ݚ�a�ɖzX0v*((0�($�Ħ�P����|IK��7�0L��1W�,�zX;@�C���+�S|��iJ���V�5��F�$d}��h�z��'�@ƯFbtW,\�͂��^2kE�҇k��y��m��J	�eR� ����:���"=p/��6��*�W�`��U��㬀�3I�ł�$�RpUX�a6���"R+D���9�o��s}�>��p�� ��B�Et�H�Ț�Rl.7���`�UC嚨L�Y�Y�X����������i��gohJ��h�N�܌��e10�Dђ/�K�)�ᷥ^9�u7��Bɩ�r�*�s�vyɹ�:��K��~��o+Em����._�M^���`�Ď�y�惟�9S�j	Qv�Y�&*�y�Q�n���Bʒ��l�ٞ���Ş�^V˺\�+<���Rw*�&�8�#�����yŤ˔w�i$�9��������q�_�!c��=�Ჹqrz�kt<��ev4G36��>���i���4�3����X4�%�G��>d�s�1ksia*��M܌/��x8@��Z������X�I�q	�����s��'],U��ɡ�@?��%`)<��1v�+���[`RK����y)�MҀ����������>���2d����!�=ӈ���$a$��2rQE����q�19Vk`�0�����P��1����\B�
I*p_(]��{4 OMǽ�?D�|�O9�۝�wK._��2�Ҋ�ɟB���l��d$�H��Icp�K}���ñ�/yf�YC�'B�v�t>b�ɶ��1׻����������Ͼ*K��̶�[P�L��B�}d%�;������O���)G�iX<)�)�/!o cd�" �5�ػr���{�FI	;�' D����M	'gK�M�"��(td��<h�ݜ�}E'�h�g0#�2/�k9]p�jl8L���~$~I�ǥ,�aX���`�v�ܱ$D2���@]D�+��<�X����HԀ�A�F�Iv2�ΤϚ?.h��<d�3r%��Ⅴ�]bVࢾZ6LR�o�$pa���i3f"����������c>�.F6`��T
ף�:�:}K�8
�e�A8�a��	�!q�Nj��RxK�������Gy���	��(�������;���WrJmӬt��������hOa`���|�P������b�sAg��n�7�����7�_)����|��9�kp'Wy���%��woj6hK|8�X\8�!f�եB��z	S�ߝ���Z������)?���B ��J+�d�2��qz������&��H�74�^:����ݻ~s'T"t=��Ɍ X�Y���9�U��9~�l��p�$x
���ɞ+zlK�N�qځ�.ׄ�vۀSi��C1ϑ�e9��5tH�bCc�r3E����WAs��9>�X�/��`���j{h4g�,;��g���z���J�m��ȅ(�� ��I��|`�K�D��3
�@"|��U^�D��zP谁�Z�=����^55~+�r2��S�zݴ��NntJ1<�C���}D���C����౴ȇw���OP��go�~��p�w�T�+nY٠7SC���{�8�ŀ�W�]��6��=_��p�$���[rK�$�>S����:D��b�q�qP���q����Y����kv%��l�����.��%R�W�:|E�4`ɖMmy�[J�*����]/�dN��]a2�!�>�C|���Hziڀ�}����lj�F�/�ԃ�@igĴ�{���5eJ���F���#�iqD� ��Wܤ��0��q'��m�Q[<��h����Q��T)z�@x"]��xB�	���K��~n0 	^T��lʼ��~�I<彌+��	���o�'���/�T����)�?��1��Ƌ�U��ۊ\޼\����.l����C���
���C��e>���e���i$.1���[�����~�dLbw�Y:ܳcn�3^��>Q|�%L�jN�n�#h��>T}d`d%����@��]C;��0r����t�w��ѩ�lQ
�"q��pD�Z؞־7���m�K�� uW�����me�'��5�Tk����④��P� ^n��$�ꊔ�{��ynLN{��S��?r���X����ޯ�8�%=XG�#���.��akb��u�%9D�w�"$ID��3�L�B�xUL��yum7¦�Ʈ��_��0n��f^�{��ƍr${#��3Q慰:�X�C�}t��x�#��o<a&�/�ј|���P�U�fK1k�S��Xrf����'�xޕC�I�Ht/�M��	Ñ�ZKW׊~.�Ԇ�{�o�@BȄ�WsɑG�#�7��ȯ�!����S{��1��l�f*������doқ�3���K��@�O
�ڿ�q�
t,�Gg��{��`��7��!�8�/ڰM�ʴZ3=Q�g7�y��8r���&������;D��L>�H��"ܹ�~�H�������s.����5S�X��HC�!����iԀ�3����"Ң΄r����잕�<�!w偶�G7��vd�a���`�@��*T`lP0qmD�������}��E<���Q`�)�;��PKa��&9{��lF�d�R6�9x��o����f!.��I���F:8N~@J�"���wVdX�_.�����l�vL��ͦ����'뉲j�)��ޙ�xk�4qs��Y�G�>dW�n��tcP[��:�cxﰲq��%�k�&�S:�X��a�N/�@ո1��[ފ�7�]t�`K��1ț\�S'L�lB���KD�<}���i��CE��>߁m�����ϋ7Z1m�I��{�_�ݯgM�'��
d�0��X���PBnU�2��q6�S����צ�b�/Yr�OG7s�B��:��_e�����` q�[G�jI��I9�[!��Ò�IFK�A��$�4�E��F-�`�Zeǯ����"�]�eFƕ>5�ɩ1�:Bv���66���!4N_)��FH~�o�E�	z+Tp�Mվ�(M	��X�K;w��(���jS�#��O����y爽'��
�.��y��t�Z_Nį��$o�d��>�����#�u���#`�	�֓EJ_6 j���0����t�=�*�J���y�d���_`�Z�����}3o����ͯ��(O6�A#��r�V틱�1!i���T�K�<���C�=tԕs+�$pP�A�XtFtu��>��(p��(�y���9V�uKM%j�ؖԯ�gd�����qv@�*�m�h�����\�7��}0�9	C>{�H�A�և��A�c��<:ї�-���*)o��D1��RC��b=�3B]�r^�U��Z��u��K|�l_	����^�G��7:���Et�G��	K������1�5��f�%Xlau���M����_V�J}�����8b�0�5p?�;Z.
�u�;,���XVL[x�f���ohf�ܜ�'�N���y-��TIi]V�=:�05�]�sLBʋ������A�D��PjL7�ړ�9��q^�Z ���Z��o� Ϭ#a�k$���F���Y�'�x)Ր�nޭ�ٳjkcc�J(q�/*	9I�����k]`��ۖV�{���-2���JU��	�JeR�eQqs��Ή�U>$����m�Ң2�QJy|�nH�ƍ盍��0��� �$H�����w,�"Y���}��/r���#P%��#�ChYj�]���nU��"yB�b,kl<i�|aZ�|���l%��J�P�CQ�_�ajS5$�%�5_H��ܖ!�u�*�#�����Yg�>���wGQ�ZI}�d���o�祰�J?<�$7_A6�^V��8�6�Ȭ ��v�	{Dp��WƼ}�ޢ��&�M�V���b�f�s�4L=y����� j�9�V��MWP�{��`��ka?�!���q���̮��i��������=�f����Afb�u�5�3rb��4�drp�.����Dl��򚤸׸��N/�V�[{F����1µmT�H��S��@嬜
�TG��a{sЊ�c��~/I�� ��-?�h8��"�ER�4�=[ük��,;ݸm?�d�ׄ���)�vc��W��R�,�A�e	L��R���K8W����i��;[�piV���%?R��Tt{k7(�'
Fx@!�[��\���
�S���ьr!��jM�݄(9�����a����f:����~��Ax�Z�%B�%�Vޠ-��Q�>ȴ[YS��\Ǩ~�a���*Fv8�<I�S�E�brs��Q�T�<O��h�m�2�=Q��(Q��>g[ڀ��6nR4�U9�y�b��uĘ	��+<�UrD\���E�IEP��HU*�}|�_�A ] Y��գ��������ʦ�R�[ ٸF��5�����~z���a�� ��#yآb��cl��(�*��s�
�����y۔���W9���rvY2�c)F�N�o�M��S@zC)l���R�YV|�C�x]dk/,3g�鏩��V8C����j�e�b<��j,��>��ꇞ
x-�߆VH��6sA�_�-U�>	]7��iq�;8��:]]�����M��rnU������͕w~�IX��g�t ^�.=�3j���B*���l�z�~��X?&�GZM�`��͈D� ��q[0�a&��r�6��a2@C.Ę)1�͗\/67e��L��<���ԅ�rΐ���A�0�DQ^ƛ��~���lIp*r���
��?#�������H[���/���"=}]@�xq5��cl���g��Y�a<Z�?9��H3�� �{���:�і� �7Mn��Ί�p�&O�:<����)�H���DH]��*�x��(,�&J�%��J�?sٛ!O���A�P�R�x��u3���)��7m�*�Mֹ�sqKd����T�ߵ�2��k1?Z!�cI��)v�h�\�uSQt�����M�p!.ZKbz�k�=�u��Q�e�^O�2~9q��&���_|�"�a�o:���x��z#���PDꚸиw/�Ş��Hѷ*�H�nl�=��4(��ަ�|yZ�:������,`��"������E!� ���զ�:{A?���gw�U"��6�g	1�wG�䓿*���0"�V`��v����cK�@3�y��7��U��u�$���}�o�Y�z���=F81�"��f7{u	��Ȕ��ᰝƞ�a���%~H;�4
}i��,������WF� �umU�0:���q�M�U�è	��D��gjE[�%��-	{�a)L}:�au�p�hug�	n^�"�=
�G�jE���Ə*c������(��eΘCm���Ƭ
(f�S��a�dU���ls����'Q�_��%�dF��w�����B<1��? (�><�]X�@�^b[�J�+17�����Ttu�Ń�=WB�BD�8�n&�j̈́�p`�\���.??�%�x��p���+9�@c�I��nL�{����b�G�2�7��sV:;�>��r�㶫�P o�{Wq=��c�mƖ8!�wlmJ9��{���i��ðWsNvK/~i�q�	h~8o�\��x����u\5�������׸&לM���e��#��:�y�]SǏD���.�c偉��j�����<uF0�|���h��aj �Me�X�'Nǳ�~}�+�ڳr=�����x��E��`��)�fxRq��"��JY��8������į�q8�SN�����|W���*��	����J�'t��8%y����<I߻MmF[�dQY-@��'�ݧ�m[��N1!Q�@�d@��b�/�z���{/o��Ma�F:o>ٖ���X���)�:Q`%'L�D��Ft.Uvu���N�������Mǽ`����` ��/U�<��̺%~�O�ϟ�l��~�F��Uy��B�U!dB�ц���x	/�V.�%���'E�H���)��y�*@n�|!�ղ���DAP��kd���x���k��T�Mث�����U�ǐw`�O�>2.�&�ɽ��Xg�8^��=ǊB�w ߶�b{��g�	�cqJ�hN1�r��{�/r��국<��.n+ϳ�`#_��_q�T5�X�x�s����;C_L{y^�.�����O=���������8���g�����@7�r��d���)S<x^�!��J+�{� �!�E�5IG�` BX�s�HȘ�K������!��X��`�s�Ӆ���'6����Χbf�.^ݞ�E��>��AՖ���z�ي7��dо�0;�Mp��v�B���X(H�}�sY�#�i�I0�}k�-��-AXTR�����Ed6L����:L�	�NjYM5'�^ObK&��0�a⮎�G�m�Ml�:�ﴛ]P�ca�d����@'��UhpDT��Ň ��E(�ұ_��u/�,�����bC��>��
|����]�S�1rNJ�u��O�}��c��w2��դ���j4<���}?�`���6}!ߐ-�XNs�5�5^�E���/��n�n���k��|��4�O�:��Q�-������D[��0�G]8�"�)�t�V�Ӌe���@�Z��h7�e���˔H}\G]8�,�G��[;RuG>1������NU�p�cNfo��`墉��/�u~���2���l�Y�!���Ř_H��ô�xi�kjzDۊ��B��"�L�Lͤ���XJU�o3���E����An!9UQ�晞OP;��S����t%Շ�n�?�M�\#ٷ1#��Y�ܭ[(��D�����-X�Gz?;�O�v���,�����MMq�²���m/I�&���,�����qt�|a=Tp�����C��P I�;�UҐ���-�]�Bm�6D�-~���� S"'�
#������ y�z�a���: �z#-��?�_SU�t�F����mی�����Z�����IYJ�&W ��V�����W:��+�����m���i*��+���Iu^�ŃK&�\Դbg�b-Fݹ�W
����bD�&N�>��.O��7/	/�0��1�_|O�l��诙9
��+_�9��F�u�!6�k�l�ӯ�|!�=ݟ�!i�ST2�ܟbs-����*�/��QŜ������1�eЦJ���,��}�� ����l�y�GD����P�%Od�#1?�+5XX���ɦ?���L����"${/���F��>�bL������!���JϠ�''��^r�r�[8�:�9|�ђn�����E<6�jzmҘ_�k�͒F�9c��ӑ'0Z�:�'L�<��ݼ�*�>�&>(o%���ۘ�����h7��%��Z�hL`#�t�1n��}��/](��Zs�h>Q�O�8��-���]�K�kt�r���zH�:&$y�6R���g�Cuf�)��wu��ą�Ӷ���'c������\� \JI�*���F5Z��
q3�Ԩ%8u��
t�yi�QHR�cip�x%�TC�k⁣oJ$�[��}�[r���� �6͘_F�N@j����Nחg|6'
@����Q�t���"�o.I(x����a3eqG?�}v�9��_�M���/q/	��wh$8&�}�oR�� Ի3N_)���#v\Wc��������"�'R8
�9��X�����\�U�8�W��xu{�c�wST�8���P�@��b�g�]������4z�ܘAbFY���g���f�J	��v��>v.amK�o^5��tC����E��PS���+���nm�1d�J��0������9��znE�+�>�&BT(��8�-)PM[�����C6B��W�u��%���[�����&E�E{HP��gM_!���>ՙe�f>�kl���H��+m{�e/% vg�xs������=H�	&'(�J�m�U�{�(q���^BZ�M's�t��g��Ƴ�-
����@����0�9����f^�\��
����<$���!�[$���C��T<5�
Yn&R�"?E�(����a2j�a��hT�],�a�js��(Ar�~��ᖩ]P�d�_�����?,�
��9SNb1s�`���s�D"̖����g �2�D���N��y�f-ʽ�5��ܞ��XfA��!c��o�X��gͥ¯����w�D�ׁ��FXW���t�X�q@�x�E��Ĳ�HĔS�V�z2��L�QE=�}�[�� �`�?ǎݽJu�k���Nr�>߁V��Q�Ql���t�vo5{3s��3\:�^�=ԪO�!{v;nH���g��j�Df*]x�����5��t/���Q �X�6���C�]�n`*[��.�7���ݭ���N�ao.nTi���b_���?QՀ��A�vԗIs��Ïp��ʲ��~�o^a�8z>��ָJQ�D��RJ�ϼ�&l�;}�ݐ/I��k���+�[K>�1�g~ u�x���{�s*����n�N",�,_��Z>N�h����U�ދ�m���,Bgl܀ᢌ�T��۝�ן[� a������qőF�ͦM�x���|Z�����b�7#Ҥ�d�+U���<�����Ww]z-��zB��ls�jB�b9&����FV�o�y� ԰86��uU���e�G�ڧ㧗>�n,�q�jNb?tr�~�[Mk8U`��zar��b�����FpD�BE߷2��-��6Hm�S���P�YD�FiWcR1�v�=8�V/@s���7����s���:5x�*��g����ߒ�nPx�+���(k8A/�����P����ي��1�l���,/� =��(�*0*}g�����M+�<w&��D�Zכm��m����Պ68���|d��'��Il��,���M��4<S��w%�1��{�i�VV0�֓�w��|�)�+���Gm��*�G�N�5!u����Ip�W�ܛZ� �� :!ٺ'��:�â�� B��Z�{E�P�lP%�����C�ku������ϋ	e$���aT�!�8��-�Bj�)�௘`������!�Xr�
�f��Yx�n��0����2�E��� bm.���JbtZ������j�)J��ŤM���7���9x��o�D�d{��~<���-ܻ�������T�0���[8��ZXe	K��}�&��3���EE'#O�+��GQX�^��JPI:�Aɹ�(2���Z���|_���:^�]�¸쾠?�rT7@����N�W �4A�l}o�����/���7�(������9�a����a1L��:�fIb��8y�*\�s�)w?�#�YK��6�.�9�֯?Fքj��3�Y�n���ꖍn���ަ��-�W\E�v�<u�L�����a�8�eaޠ�P�q/g��bΏ�g*с]̲��p�ϟ��o��f3�a%�羀��;t�b����mH�]�ܖ������6�{-�P��nt��oT�ƕ�/��*pd/�A��~�kfZ�]4���I|����ֲz�+����y����q�_��&w<�*ȡ� +(�S9n-h���X����|L�(�5���_V~��ű�	���!�0���������$��L�����
��vjX�A%b*c��t���ж�y%���`���7�-]S����,Rѯ�i�~J�:7l��W��g�>���ĵ��G|��"l]�35=<�fq���M�\��w3�!S�Ñc6[�d]��,9'�M��Z���^D��Q�N��Y������у��]h�͏S���oACS�t.��;���1�(�Ȍ��� �[;EښkT4b��!�1f����љ�k�:>���a���ȟ5�fOM;;PU/,�տ2�&�3�������=��_(�ad��"��D���ٶ5�136]�5���.Tݛ{p�k�p �0|��%�m\���m������։7��ƥ����a �
�MWwu��H��{S���S�[B����E�V��X�Ȯ�:P����^�V%�-V�ў�d�����B]�(C)��r�q�O3W�}&Ca0R� ����\1�u%A{t��e���\|���hμ��+����a��Z�В��$�m��G�!D�z��5&�xu��}Q�滟A)voC2���N�{��C��P?����#���_?����?�Vx�&����C1�	m�$�	�/�d_�G��s���6oW7�<�qH��]���_Ϗ�����E�K���HE���5�m��$�*��|@+(�Zeb34���s֥�������,Q�ِ7��V6Va�����/%����KJ0�Z�$�a����_���s�}`��t�I͢�a[��Y�;W(�0��h���!j��6��0dѧ���z��4�����%���@�c��DAO7�+V�I�o�2R�� *&Dv���n>�2�n+o�������Wi�?_���?������NT�m�.�m�O�M��$b3bWF6��zY�l�8x[}`�D�D����P�q1���O�&J��Y	j�b��Ě�b(�#��7+����Y6ڃ�Dr|�e��Gx�C��@�I������/��m���/�_fQeh�]=�?`�kk��3�zH��;0��]�&�
�{�G��RD��,RL�L�-�����lS�=H��Q��c@�G�×��AY����~��iY����-�|)?�wP^�s��I��FXR�[�^��_����$3����m�[�{��}��q`�q�#�mD*�$��S|C��]���M����މ���@88���O����M�];kW���'�]����S��]�&�u�9�:�a��xV"V��sǜ�p��>e�_��A�&�Hᡔ{/t�7���=79Z�+s�$��^�-݁:����,Ԡ�*���v>��Li�tkl��kho�� S�p�kj1L�9D�u\K!�΂r-:��a(�I��D�Ơ�u_���R��[p�_�"�(�k��ڻ&X�:�ш�S���#EZ7��E#Y��(r�Z|��!����dY�C�npN�p��At�%�ذH�5�Ŋz��f�g7��#�U�\�3Z�
�Rd�/D	t� 0��B�^!�i�k�Ԉq�(�7�s^�1׻�������n�/V��Õy��o�`� ���AE�2bMtZ��(}��'{�ԡ��P��s>��nM�ݱ��5+�{����G�6v�y�r��������@k�w�y^7����^�N�h񡲿�ie�Rm�v V�g���pא�bi���d`y3[`�A,��Ë����iZT��.�S���A�Q�!�iX�6�:�1�L���ª�P�((S��S�aZ�ߴ�KL�oT�$�#J����F�?�|���㺈.'�r���~UI��v�Z�+�3Z��z�fM��_g��xȉ���*Ք䯏� Z��Pse�R��2�,�/�ʈ�����#������5���0���q:���{��4⑓�_�6�[B�=t���>i���s9(�	��Ƀ�)���E��887��Rmj�N�|
�,fR����Ge2��R�*����ϼ5��mUh�u��7յA�	��N�����xבj�u6� ̀@��}��T�~U9fV����������Co>��<�z�r���9rc]�r���E�Y�39]�gH�����CJ9T}�wG{d��`�amv'�z�_���<e#B��X��5�x�8�K�=�*�(8tv&~S#��*D4�H�n��c�Kܳh�E���:��?��h	����%�^�����Y���(�X��D%6��/VkB��`�hj�������s*�ѓB!"�~3#<>�_�������BN ��g2[Z�<Q]�ߎ
�ܟ��,������̓(�LH�)��}(�/qu/��snĿH'ED
�
q�����j�r/���8��k\^m�A��N��m{�/:˾:@)��_b�lC*x2����6i�a=�2�8�w���7�1�󢗇�(_y�YC�oT�Z값&�IY����İ�О�Ӎާ��Lh��G'�H9T�_�d�$>7�c�y��?Uw��s�>�#Z��c �)b� ��$q�t g%�2"��b�ou��ͮ�L��T'i�	�:\��!�!��9/�i�T��JJtB�]�va(��M7�L
3�R��5.9��Lr�R��lM=��?�jO�j��v����}���n�}YY�5�"�
㘬(��,�J[��އm'���<�`� �>�+��{a����T��]j��ՠ�[�r�}JGV���Y �6��X�Cyߍ���ٍ�zM�����K3�����7�8�s�G ��U�:�r��s�w�~ww�ь�
�[�M��Hv�Nu9�@����i���L�������Cn-���sm���Z��2���{������Z�t�"��㛜z��6`���m�,�ce��2��]���7P7��Y	���<}bn�п�1;uU[=8-Ӗ�18t���F]�� �����袎���v��Ò%q��IW���wy�&�sSR�������7SX��v�[zB�Jx���𭹄j���3y��!��{wtqNL(!of�P�)���?ĥ���CQ��m��X������icP����V��
�Oh�������,�`'�^����tyy�DS��j��b������3#	"az�U��Y��Ϙ'!�A]�	���1ʡ���_�-5��#5D��Υ��Fi��K��W�8���A�x�hB5X��g3v����ht���ү�I;� �	L2��?����pU^UY��oS*7@�0�3L~��@�C��
.�Jz��tN}LF�lf>�m������iwt{+ɻ>5��ۨ���/x�� 9@��Pbg��5���u�0�.�������05��\��p�q��q�Ԁ���J�	�t��+������D�*?�s��E�²v�J�o~k�5���NQ�q�k�������=	�Q�C����u���@~}i�'�t�LD��*/+8�M��#/+�.m�5���}ѯE�IS�{=w=óH�;���0�����	��B��W3�^ �T���k꧝�]I��h���o�e^x����@����0e�sQ>+?Y���^��0W} ���5��#�ׅv�u�F����4ǎ�7�/\��#�-�k�&��Q����φO� �29`Ł��3���b�U��zP�|��,�Q���r��Cb��Ғ���	�ٗ�&r~R1�G������4/nw����9�4jj�Ӯ�9J݁��(�*̈́>�����3��{C�� ����H�:�`��r���cɔ3�s5���7qW�;?ۼ.���UQ�<Vgp<Z��xF�i]OL�  �r����m���2*xޝ������
�T;�j�-�6m��>�*4���4RQz�#JН�\m��;pŷ��BG�k�I�]���Bgȍ4�K�ZሳNc��� 7��t4�|�	�V!O�:!�if/��T��jr�mF��^���{-T�,�i�Y.�类��)B��it��Lark�.�ϝ'��,njp	��^Ba$��~��y�o^���,�%�+������?/d e�x��YYe�j嶪&�+�4��(�p3�L-e멖��<� 'b�D������	�R��H-2=I���~��E������P�%]���EuLT��H9�M�g,�𠅿W�K�]��aF��)�݁�_3����bS�O��D�EX�F�Ƚ�J�JfG�9�&��>��3�F8�j���q��+-	A|����Dj���H�5n�a2�Į�v�l�Q���X��lW�(��S�:�Q���b����ɞh�9��G����5	�(��zU�2'o��.-w�,�x&ǥ�.ϩ��Zl�5l���y%�1�t���i�Zؐ)N��a�i6q��pY�#�5�0�):b����(R���������I���IQ�ܶ�\C7���n��:N0�p�׻>@,1��n���n�=[�H�;�`Q�g��|�+��D�/�m�5����=p���z�S��9��Ѩ���N�̬ˎX�C^��u���Rĩ�Ѿ���	��V;��������*��a���ӎh�%�N*/`�	!�S�i��4�Чm�8�fg	�,�p���UQ����0��r��K�LJ�.NW汶Ghu7��g>�f8L��	�Ps���06�Q<v�ޘ|��6,�����������[z�L�y�c��TYwR�Oc���1�o�E��臭:P���.�*]O�ae��^�� -�H5㳥I�R:)�1NME�<ŻLf2�`j�����J��ٝ溛ltlv�a6�7F���h	�J8���1���Q:O'�H�h�n,�W���`)tI-V6BNJp5��,��'�D	bs���=�>y���aubz�P��A��� ��H�z�e_�t^+R$���O�ts�9cB�	�(,������A���01~��ɿ��t��y{P9���5JǌZ��݇]3��i�������z�8jY�K]�gA��N�c��Bʭ^5�\���u�*�Ҩ�63R����S��f���*�'MU_?�T�j��!���dG���b��\f"�[���gѻ	�/Y&�1~_&z��dX6z�kf��{�Cz��pt@��˻����Q~ٚ�����h���W$=��?OވZs��l��.?{T��r���Ib��k%�䡏nX�1�}f3:�#���pO���z�_���f�`gMs��ٷ��{�fz��@^���о3&���g��Q�1���TT~"o�_B��s�萿�qW�۽M�N(�'ڙ2pj
��W��fϡm%�@$�W���Բ\�|ID>�j|�G�f��:�=��n�*}�}/�Iu�Ik5�2�z_�Ae�rm�;��SB����~Zq�W6'��S���<?�I�m���-N�n�� �{G����D9^�Φ��
QЛ�~�]��gq�g���FVx�낥������g�3La�;3k�6 Bsm�jWo�5m��ЈK���D�Y+81�%`b����t��f�2֟UKW��*�V��04�f��^�qt�Kp�C��5ꬖ}���Î"��0;%���`��%�m�Y��ln(P�b�)S�/�C2���'��r}(sZ�`���/��S?k��T_���d�����s�8�J��%�!.ه�(KR.��}����o��E�D�75���T)�l��6�D�u��m�+��x~zs�%�;K���Lq"�p�=���MՄ�+!Q�,$��[��l5c.)y��9�f��|x�B��l��o�v�;��4�����<�l��@�m���?n��i�[6��M��n�L�r����l���f­�G�����-�$��mnP&xy"���Y~l7�
�^����ib7	��vĳ^zIw�n֑D��w��^�x�jA4|ʧ�mT"��{�%��� �^����-���j헝ԫ�{`�Ĩ��Ϗj���;� ���k@Jq��$,�f77�ڷh��Yw����w/���0��B;�K
^2P�Q	�bX"	M��ڿ���E�'"&�����Q�KW7�ڗ%j!���p�ӡ-@�	�"�Թ�13�̒*wAo_��b�I~�C6���z��Zy7u<��K&k�(�#�,�4uV�+�\l��4���P����p�i��Q����4ȡ�h��zo�b��@O�b�Ҏ*�S��K�-���@R�{sFL8��ͥM����c|�@��"������o"�����C;�PA��1�Q8������R���2g�y�������r������`&�,��ql�,�6u:~���Nv������y/m߭ wI�;7~�
e�0j W��r���J lS8X0�n>�{�����3�_���@�����b�y2Rcpt�F� ��_���KZŬ���^M����ZZ�Da�˥�[�ge��<Z�L����ay�`�	����:�s��%Y�X�?C�(�7���<+n�.c2�B�6�WT���������l�y���[M/Z傞�G��uY*�Q�K�К�Ч���u�Ʌ�4ݎ��g�y$����4-���S ��u�܍��i��q���
i�l�D��4�i�sr�W�gC(�c3���O�5���|/E�R/pc�������Q�;%:���ID����>-�Gx���(�P���d���L�g���#�Ej������M�U����r�P�!!64��:G���w6��[Ym������������4i��$WĒ�-g)֣��Ԏ�p�ۡ�x��2kb��r�dL���>��Ek����w�o��Jm9���)�0�4��ݴ��cf}��%��;����\
�rx��n�$6]��&��s��?��!��-����?�gX��g��c(�}���ڮ Έ�Z1!|Ǧ0J�
P�C�V�k��Mu�t �c��9z5�ӑ�}M�Πl3f�*)�j���.o��`������� V��{2�
I�����J���*!�I��Ĩ[�dJs��̫q�Q=c���f�H�mT�:��b�WH�Q�g��'hJ���O4E/�	��tsz���\,�A���F��l�\���籀]Z�9J�W�����VC��fG�U�L�v�wq�D�N�l���Z��궪���i��v*$���D���6B��@dMd��� `�$��Mr24������D����8����ÊWQ$���?q���(���u�D	Wp�;�P��Li��q������P
T�����/v/E����Ϫ�rl� �h�	��YJ�	��T�K�8��ɹ���1J���!�pB\~�"���DX
-ed���Hk0�:I`1>8�zm�ݖ(�T�Z#�����^q��æǎ ��i�f�&����e�����r	����6+H,��Rka�J���'ĸ�ԃX��9nva R�t�TÉ�b}���6��hg5`�Q���^�ŧ���� N�V��c9��ڱ
M��z6���q+�(	A��Ӹ	��"��a 5�KV���E ��hh�>���*F�:��ḃ�����X��~����K�KW$'Jidy���m�G��쥮��u�8sTb�=�1���N�s�\C7�m��C7&������B�@������m�����[�t�g�a��Da 4��[��=�+nxȤ�;g�"a�@�- Z��De�5G���Սy������4�+����gb���%N7z?JE�]��"����ol���z4{ ˜^�$�'ģo~��P�=��.벟�r��y����9 eQ�
�ԸC$,�p�N�,c�
���:���Scu�R�C0\�]'��k3��`�8�	%� ��M�ꌁ����D뤽�r��ϼ�2�{��`��kh�.�*�1�I���4ơ�:�_�L��]e@��N!I~ͻΎ�~,�6Á�R���1>@�"b����ٷ�&�����W�}A$�q�H�߉�� �����Ի��'7b�{��kY������1?��.�+yc�z����f��*9e���`�z��~FЇ�a�`k5����¢�4��jEx^i�^��y���l��N����8��-��Մ6�,!�Y��V��5$r�>n��9�����Lұ���"��u?��!"���M��B���>� �>1"@q���)�c���
�����O1f_��@�xt��V#*�p�@�x/���ebb�$���[��f�Rj��ݰ}��R���U"#�.0 ��J��6=����{�c�	㕪^
m#���9=�d;d�}.����<�"B���Zv���`�,�:����i�yL`@lw���;T�R0��̜䈿�h^�B�A<C�&)�q؋��c�����|�qI���4�e"��v�V�B����fSΩ��*�pQ�	�*���*��zץ´O���$.�7�9��aE`z�-Ttc�6��*�j>F�k���_3��{B�^�����W��)N9|�sl,4��9���QYvΝ�U�({n,% ������}0J2�g䵜h7���({�������>Z�`V������/��I�Q� X�$jf�O�,�B!��O7ߒ��!Z~��{.�
�����F�	CbY3�L� ��	�G	摤l�yF���BF@���5�:��D4K3i������	��s���af�Fƾj���
s�g�&$��Rt���ttf[(�I���r��
lJ�m�'3G_S!9J"&<��O#�Jʈ�g���lƝ?�z-�����loH5q�^j	PeY�� i��ZcȌ�d\��*WQ��к
?�jM�йH�� ���o�Mؚ�W���8���@	�Ҋg�(��S�['�||�\,�_�p�(�pg�xb8���;=�`ٙdp9Ujh;���Z'�d�r�����E��/�x�r��K4<�z�����8XZ*��uI��?s��C�k�����lsClvt�H8�;5����l�7�{����Uo�fe�tm�go��4���F�M�w�>lm������7��u���R�c� 3 �N�K��ck�bl�-�v��?5#�#��cN�e�t���DX���o��8k�'#w�M�O�t��F��f��t�
����O��}^�P�����m�Gj<[��ZI��
]᪰��L喙%tMi������}0��kwu����VNu��[g*	���
b�X��R��麨ɂ�mO�-LR��|�ss�S*m"�D��X���"��+[���!�5��&���L���w���4�39`^�wMw�O�}�T� �x���aM�#�f%�I�Y�j.��!h�*�ۭP�Jn�a���#���a2+��X��y����ǎuE�_w�>}�
Kz�웧�-1��a�X�rPW���tI�Z��+D���/�v����1��q��2{�dI]3�h�2ǧ�i��Zà��E؜��xJ�Z���Zy,$k5)LW$4\HH� ��k��5u�t|M��]�'�74�n\�%�a(s~�M��ms����ӭ>���i�@��T��n���2Н��L@�5��	��d� :�`m*����f'7�-��
�O>��5P�E��|�ĦL%���ȥE��S�.v�_h��X�pe���<no�$���i� �[m� ��ٻ�$�u]�&�3T[��|5��ePg���f~}��к� 
��鹿�ey܎fgb�vC+����	1b�I�*���d���G�Jk�6��=��}_�J���`�n��W�	ʱ�*q�Mj���	�S��Х��L���m�M�c�D��o�VR�p������ݦ�m?������}�3�`��6�'s����Xy?~�V �Ծ�N�*0�uԼI��|fe��_�h�����.�P���ХmrL�f=�I��(�z[����ZҎ5A�X*��`⨛�C�uhP���V����$���V��J��G���V�$��'���!~ �uHs���ۼzT�"�0��w3J�ӧ����Ԥ�|�1����$�b��}�[hr�O4��j��1��$��xAe`�ಟFE�pd�V-���0R�7�r�hdaR�p-+����&pJL�y�6����H���*s��!��& :�P�i+H���ߑ��x������ ��߾�Ϲ(��PX���HqE�NIݾi��6k��X��|��h�j�Z�@�Qq�u,@d��K��N�[����Z��[IBt�HuT������� �nh����HR����6FԹ��uy��$<�-�D,���x�6$�&���=�8GЌ	������ӓ{)�u/�'	��]���_�<�t�N�����1X�Se�C$�h�u����8#��ݏ )��8Y�0|�05�7��۳G���6�"��DӒE����R��ӯ���>�p�}�L�j8�}|�Z�Ci�����H�|	44S&��
�L���z��59�Y�a)��"���oHaN���b��� ��a$V���y��=z���L�=���s4Ԁ�b3���jB�i4
>�,ߤ�������m�@C ����'��G��/˲��˞籔�R=��)uB��(	'�y���/=��XM�����:Zg��uM�s���(|��z�6DQ��g�ۂ3��Y�lӻ�����������@XL��V��9>l���V㎣��ms D� �~�sUeҫ��У�*$V��`n}�5��=Fw>b�Y�>���V�A�����Zo��G��-�y��LB��.�nS�Eb(љLhR�hE`��O~D�҈ՆP��֕n��egw�5�����9"�\f� F�ΫM4r�?Z�u�V`-�g&X��w����!+�;�x�"��=k k@t���n�f�d��̾̕b1
��A� I�(&}�h����܍�ޫ�=����t���|N	�R:ؐ�t��cmN��
8�X���?k��Pԕ#�n����ƪ��\z�Ŀ�)�Wd��i�����N��F�*<�9�=��'�	v.�bL6%��<m<�q�mL���3��"�)I�\�6�CĚ�qe�qR|(N�ʒ�������}t5�G��J�P�l�?��[-.j�_��Hp���J��`������p�	�j�Ǉ�y����P!����]�4����pμ�� ���ޛ� �'f�����,�#�rx#qiG�þ� �Y~�MqD�GSʴ��ú�K#�F!�B���>}��)B�5mx� U+����M}�;�:90#��m��>2h��� �Ber�i,���![~�eGm����1+��X=�_2�&�v��-��*��g����:.2e�I����m��%ȥf.��e�x�I�
��ޙ�&+Sq��h�Yu��;Bp'n�ܧ�4�(�RB�3	��Ѱ.^��NfgL�o�%�@�ZY0'��fXւmm�Jt����W�P׏=��+��q�������E0Q@ ty���L��iJ��p]�x��yO���&F��W���'�.�4����ԕ�Q��ڦ�b) �> �0�������1����եT��%�\�9d��& ^����U�E�p'\���?)�^t�'��o�?1�ͬ����pH��Y;p�v��|�"r�1w�}V|q� Y&D��aU=]b�o4�?��4.t�[�V����A܂�U��g��eIo�C5�i�=�:��cɽ� ��߃jdc��b��53S+ZR�";�x��N��W�З��
��+�I�U�#!p��9�݁M�Y7��}w*Z���2|>{!oiZ�(��8�a��%DIc���yC��I?l��zI�a��(A:���V�.����F[��� _M�+�0����t�:C>v�H��K>m�����_ȎZ�#��e��1>��$M~1:O��-4����]A�����ՎM�Yyt��ǰQ@#��-���=�ΓGes=�dF
���.��
����|�p�"<њ�v)�w�ɌpM+N�'��V��@���	�34V ���Ҋe!����r`�@�#�R�j�1�:�K��#A�CФ �>b��å*��>�:��`���샙y��r|T�(K 	0Z��LE����]���,�t�/���a��졎5x��Q"(o�|�ϭ�ۧ�C�i�ʗ|�5�(�ƶ�)h*e� ��-����>�8 ��m:�=�6���R����"}�#|T�@K�|�F��-�R4�5�B���Z����ۭ�	��\�A�q�$����pm�/�!�j��$��o6�!�"�5�����������,B�,��˻��J#E��=b�,*\]��9��ȵ�ޜ��)�*c�r�j!=1d	��/���o� �ߊ�c���B5z���V+	)���O7Rq�_N|���=���u�c�q�M�si��&��#B�0��29S�v�$قXZpn��o�byV�U8�O\ܨ0�R���9W������p{�!K4`b�psC�_x���/N+�����r����o`*^��y��jKU�U~W/�)���0�*L���Ɩ��y�kO���7^i_L�\�]�dM�z|�˟h��N/�W҉yF2�D���Ք�Z�+���^�.N����KYۨx�B�⥛��>JD����śZ�df=�vF�8d~F��`QϬ��6��慄��ˢ�.0��d�6���ٝ��dVa�T�c��-9���l�^��6���3:���bf�1�̴�b�K&�};�P5L�$;N_~��^S/z���|�K�ƕdh9U��o�s��9 Z�N���=_<Y�L�K֑	.��߆�@"������g�iЉ��ռ�	�X�^����8�0iG���<N�
\��=���!��l
;uA���f§s����W������ ����:āI?�
e62l��6P�Oy���6�emi�Ȃ�ȡ�oKbCǦ�ml�J�_�������8���t����e�b�h7'���Ǳs&Ͻ[)����Y��].�t�Ϛ-=��N�XH{,�77�n�~�~��=Q�|T�߮�[�����Ǻ�6�Ej�,�_�ܕ���hkhe�;:�Г.�a�	����^���j]��W2�R���U�J'���ko�g@�,����s�0��$y�f
8�e�����"�1��8s�Lv���F�P�y6~jJ�l3<J��e�`
j���[�$�ژV�������g�o�l)I�oŉ�?�Y���Ǒx;~����`r��o'>�sR"(���ǫ��)�=I;�sZQ�V�cQ��
~�B�P���FVG�����+^P��]vX,���Ix ��؈� �a^Q�q"���c�M��ǭ�7M��<U0� -�tRBW�`le�J9$�:r�4�#Ώq�b��W�s$����I�H�m	Ѱ�vc\p:&wp��ѡ��Rzn!ˎ\)&B2�h�T���:䫣�J��ihy���g�F D`�S02��Ȋ1�����C��;$J��Z���w��O��p�o�m�$-V�����Ψ԰�qF���m@�N��2��U�m~����[l{�IQ!P���.^��sytvS ����R�b���=�Z�]��rO���E���Q���ubmU�^�~�R��g�g2����ζ���s��Wຆ�M�?�&`��p���Wn/��G�r��i�������z�H�:!`1����QK�C%��K_������b�{�qZ�i�].�r�������b�h�a30��Nd��,����@�&-���MV�V$��v`|E��������黷Фp���"�G�i���Ue���S��+��r�jA��^�c5%9����EӧPPl}�x$p��u���Gc��$��DCLf��l<w�5@]
�>`=��r��x���r�����[8�����7ԪnA�������'�"saz��!�g�`��fb����<&+����
ɵzߡ�����ai
'�����!%<����c�}���6{����hƠ�P�'�\[��$&�&|���o��,�uoU��1��VG|��5���"�-�5"bs���8����B_��L��Y���?�K�+��ji�j!&���	�6^�i���`\� ��d�'��Z}[!��W�umj�����5��!T����u�"�:�E*#�;(ĺ�S��'K��-Ca/�'�6/Ŀ��L2Y���.��G�T���O`b� 7�X�� PӃU�q�Bz	�~̊�q�c�Q�[���]$"�S�Q�{�.�������Ȩۆbd�:MX�{ԯNi�ȟHl��p��m\���v$����U^��5�����8Q��"���8R�o�B|=>|I�����*��_RQv�
颺i �]Q@by�B��6�\�0#�S��c�`�U�	��uܭ��;D�Ieʾ��{��R`U�V-?O���B��0|���o�����vL�ǹO��2��5;/��'J�b�\|n@��,�U7z)0�m�#Bh7�!��/(1��l��j�P|�8S`������ڲZ������!��+ N����~�ޱaV�����Cng�f��lDߗԅ�+�ƜVi4�Y2-;��Tr���g��Z ��8���SP��/��N�y�݃bjP��8�Ο1-�,� {P��K)��F�W��8��2m�@z|��@>��l��h����+��@��}4��W�H���R25`�RP=�y��(�u-�*�!��Z��~��B8��I���~w������!��p��6�Rm#��ʈ�z��#Om�H<�VTj��{G����:�}T>���~Ȩ����p�m$��'��2ďUJ(��zL?�vM$g����Š�e�Q.}�?PH:���`!��oT@��t����P�S��\3 �.f��FQ)��M�	��.-<v�X���qCN��Ë}7�E�Cn��o.�����,+����kP�G��'q���@Z�o ��[,� ��ٗ�̲�f�O�e�U4v����qy3.��Ę	5�lT=��&�w�FW�}U-ͪ"�(-�ue{x�\WT��b�8��G ��PԻ�X��x�?B��E�H��~u��65R�)r�À�U�L�GC}bW}�b��i�V�l_�)���
�������N8i'�-���Ԑ���Kj�Os�^n((B,fbE�hB6�(�� ��p��b�S�u	y��P��pOi����J��]3h,����&��p{�����/�L�Y�	�'?�J��r�11�{L7�º우&�������9["�>�i�R�u՟�`�G%��u�D��~�������I�dl\��zӃ��Vc,�~��Io�]����ktB�Rc��^�3�"��y��Z��bK�Z�ł�ZX���b纖�"ǩv�x�>�Q�Og�yw	T'�^WGv����VfZ�B��z�'���;�E(�;��_�7��X�{ɧ����T.�wV/H$`�"�4����3+s��진��A��B���]	qi�s�c^F!�U��T���`�=r��u;��4w�~�7}��g���O�l𪩋5����_�%7���:�#�x��ɒ�m�{�;���(����k,#���@J��� ��j]�Z�����碢��Ee��G#%���-~5��"��z##J�3�K�u��!��Q��(ݣ�Ks7
�;vZ]��l.6��6��Gl������佺H���L���[��J���W���0�/F���G�︹|�	Ŋ��N�����Y7�ۧ���(;đsq�����7I�7�^���f���pJ�bjm�|k��pDiJ����f\��\޺K��]?��e7����Һd��9��
�>�P�&�N	�_���#4�/ٓ��fl�O���a���v�<�ĠcZ���5-0�̺CYŭf�5��e�ґ2���Yz��Ad���7�yl��,�d��/�!^���k��tae��y`�*��	�e�������Rg��
'ѱ���lUU/ܳ M_�뇹.5)�Ԃ[�؏�q�S�y;��a�
Lh$��C�I�����^�6pJv棻1H�I�>��OM1:�Q���rQ@���y|ԕ�x�; �30��<ƞ��H��x���E?��H�%����T�&g��)`z֓,����H��
��a�ߟ��'͝J)ﬃ���U\B��A�
���=�,Qc���2dy��*�]���7b֓S���܂)�y�d��x��&^7�k�LNX	GA���0�='�[�tN'0�H/� �/�&>��d�q�2�0��fh ��ڗ��#��ψ��t�p�i�y���׉���BX��t$��k��IS�D�=�2�[k�����-��2Dq�Ҹ��Y��F /��P]�(%?��P�Bm5���+�Dj������ ��TOǯ�טPœ[48hd��;��v���1��(���3-���e�d�at�����.sٔ:���5�DF9�����y�\���mk(���G�	'-Ŋ����"�g��'m]b@_/��@��hH*qeV�y�=Sx���c���~K�mGka|�sly�Ҥ3ߙY�T�ˤ�i�~3���m�C��e��:��Omx��	pӜpv��6��ͥ7��7�qU�;�rď����J�y�b�R���?��^�i)��U16���H��/��[glF"�<���+�]P���-�u,��^��Y᛭�������V�Qp�J���*I�̛�����[IdN�FĻ�X�m��,Y(GPGn)*k�Hr���21z�̀���K�	�:+wBDw��;�p3����byψ��HI/�RI�j O .����ӂ��V!k(�{\��P�Ü��ku:c҂�V�*L��$��</h7ߗ��۽$�M�7���F�|�	�:8�?y��<�Q�uc���%��IP!�C65�Qk&U�LlM���{a��O멛�N{�{-��S�\�f����cL.���"�U��7��T_��O���:e����,�}۾��orݔP�v�5���F��<Gpv8��T�&��N�
�u��zu��4�#Nfz���j�G�h;�0<�r��Z+n[����ĂKP+^�$>�Ƀ��2��9�nJ���3HCWdl��,o��3�ȤTӋ���wc|���s?`��<�V(��S,�"���窜����=�t�|L����[_-�ׂr��b��y},hK-�Xk|fk� ϥF �]?�m�c�
�~��E6�N�A���M�#�(,����| �4�N �Y|
Z���)��2M���6&Yٞ�&F=o@�{�d3|i�t�BM�w�_]��]�gv� �K��X�uWTÍ.�,H(Z����"T�,�v��+Y�`��H�e��/��ׅ2�M���.���Ѐ$k���A�]���q7�Q�#Χ�݊���&~�F�@!�<�[{�+�u��#��0�^��hf�{�ͱ���F��|�;M��h����%n���+=���n	^N���c��B��3z$#'��=2������P�oQ���#�.H-[����j�$��F���� S.�� ��h���Ka�D��HV��6���tj�C�oJ�]B�v>�g9lQ��&p#] ����s;EG�lʀ[�M0x�p���#�)rE��`�&���)�t6��n
�UW�	O_����cK��T�=Ǚ6��u�ѥ�D1�iB��Lq��h1�`��Z��>Q�I�	r�q\����3���"^3r
�:���I�Je�8O�(�7��c��C�� (�
������m�3$_��E����
s(J\�!��7�QUE�y{$U	��,2��B��w3E�q,
�l�⛐賩��U�M�9k��1�%,��6���W[P9���]FMJ�E��'5mLgB1]{p����u�1B����K��nj=�<r�Ew����;�~9|���m�k&arOT��>�����؁a��1�βIJ���CkL�8�q��T(5��!ls�E���V�N��� �$E�~��9�\<����Ul���GL+�ˡ�8�.��u�`��J�ev����mh����T ܢhH�1L��R�ed�{��[�D�ScHE�YF��׃"׈�W�C��.�"�a~m.EY�Dw�Z��Y�|�WΆ�#ߩ��.���XLjP�d`�E6�|���Jxnm-z�����aɽ�-1!������L����O��c��!��C�Ȳ)S��V*�\��X�>	I���v���4�>�����ls��-���	r0����7��t��)��0�E�Ӻ��"���v�Է�!:�3]��^�n/�0u�2[�^���⥂�ڭ�s:��;!������X���ا9LJ�$�v݌�N�F8|��(��݁ 0X6���g{�@QN�M3{����d�O�n�~��3�>�\u!��!�;'mO�3�G�x_�I���IL��/�]��0J��(�Ln��x�N]C���沗j@5�����z8�$�a�M���p��c�=xp-���5�ӷ>C+a�U�!NMH3`��f���|�ܕ��a����?���wG��O��qY¼�ދ~%���Kis	;�k�Ռ�m�sCi��d�e�<YOLWxB4�Z'��������6x�43��U��U�|p�́'e;E�w���V�n;�よ@��1]�g!���OvL5;�m�ѣ�c�-����6�ȟ~�_O-Q�qX�.N��Jpn�/�xTX��g%z�%��cQ��z�`�מ��1G���F��u�}��/Q[��^ly�f�>���zSH�>��,�p:��#ف�VJt�����@#�~x����M��z� �
r��&�a��
��0�b�#M!d:�,J4l�� +��_7u��}Q'e�,[��7���I�0�2�q�nZt�	x$8�,-��Ţ�{a��RŬ���}F�9����F��i&�\�)lG-��ѽq@�"?� �����'B]45-��n^}X]�(V"��l'����[�S��i�.�^��R��w�x��!0c����~�s�e̮uH�/�l���>����H�� ���)��E��{2=<��6|�6�]�B(��?3�^���?���BB�`/�G�D���<�!"`G/=-F0v�L��}rK�4��U�Me�&2�Y��߷�T�^�`I��_���/g_��|�6��<ԇx�d�Щ�W�N�8����O+�_������t�HW屮�h^�U�ɫ�����7u�5�\���$�a�*�AB7U8a��w� 8��aw$���ǉ�7@�邛��0 � �LV�t|U�ɻ3Bc�<C�ۑ���%��bGa]����%Tɂ���݂W�,�����&��)��C>I�@Z�k����,Z�}0$��m��%rr�S��f����qKf_B4���3�v��\hN�uR�t�������G�
 �:2}(2�G_4�3?}[#��K�T�����<�t��+�gh���c�J�u�!b�H�۳���Ib�U�o�v"j�u���Jl�`׾�U�e��Q���E��C$�ϤB�-Իxca!�<��T�S{Z����H�KK����ƙ�mݔK4�O�x�$�E�z�#ZL�3ƈ]$��MY� �LY��z�%���t�Q���DJ��FЊ1��|,SB\�V���:�[� ��	�Z�R�O(V'�0Z6Y��ʄ������%S��h8}���'��є��ϮQ�o���-*�O�| �����y-��?[���♤c�f��������T���L#����8օ9�����F^8u��z����q}[	S]<x{��PiV��rqs��Da8/TS�X>x���u�@_S�9�#�E�r��i4-��}�*�H�<����6A~�D;��A&����ۻ����������'Ib��ɐp^p����W��.�k-b���ki/��pc��v�D�S�'1b�_���$4|Sa��٢$ʨ�ԋ���PwI��+	�u�;���Z��6p6�)��9'�T�a����Lc�}��?��	e�1cC���\��m��R������F�թ$���C
k8��Cd��"w\3h�E�?���kݔW�{��`�R�\#�%�r)ŝL�Fd�� �[j��x�61�.�^���r����M*���l�۩`'�	�3��JO�P��.��x�u��b}k�~��5��̸�Q������� �٬vQi����R�0т��\"y���/-�
��x��@Q:�g�n��nU:vj������ƶ4�OUۚ7ȤQt�D��'�Cpk��|��Rpɹy���o!����~�ݍ;ܙ��:i�$A�j�Ɂ�-**�PFFet�}�oR����X���zQ�����l�Jֲ����6Quyk~f��7Cv��A0��kF� ��Em���q"�#���H�h�	�9W^(1��7�|�^�7��o���AR�� & ��UN�Ek":�ci�&�u�Be�R!�n��}o�;sr�Z�8���TT�C�nɈ��C�@ �Y��{��d�cj���Cִq��� ��32I����&e���	�k�v��S�ĥ�4��WO��ьp'.pz��yވX�T����t�����:�^cG���R��%�	��Ep�8�����V㥀'z�5{��[|g����A�{�.���$Ӧ��;4��-d�׶���ՒG�u��_J��*ጅ,�����yQ]�0P}�u44�d�B�����c�L���_��IC���S�T���G|���`v����5u�f��ŏ
\��嫙����}����ĽH�/+�l��hqak@���UJ���.sM��L��;Z@gv��"�5�N�xbE�����GX��( �K�ẫM�)HL����<�H���0n+�4�x��f%ݭz�l��;V[R��0'���O�Ŭk�&D��n����ۋ��h5e'�*#φ9_���N�ibM��(�`G������o��z��d�Hx�Y�S*������m�De=�Rh3������	'u)�Z�W�!^V6��!�X�$�Z�
D�+5I%Ҷ���Шb�?�J�4SQ*������
�EjyB��># �7��������VA�!C	�Je`y�b�j�<��4|J@�a�Nb"r�d\�l�*��Q1v�M��?fַc�)���a`ʾ��uڕ	�A�΀���Ͷ�׳���0\{ί�סD��t0F[�r[�M��z~��%P����p!��l���9�?�k�� 41:�bw ��W;��rJ����w�%�k��4� F���AM�no<9�|����J�����f��AoW���pgFz�)8����6e4��cT������Vb�z��)��o�e�ء�h������gf��t�B�]���gܗ�hs� �5DG���������73��M���)PEl#:f�S�W5ο�� �!�S@��Tcļ��,��F%���/�}�VP���v8�F�K��WQo�O8���e��M�m�b���J$��Gf,�(�.���Q緙�%g���]H�1���lUc����8��)�G������S��f��;���R�7���Ƞ���=�F	t��Gw6�B*�:
�a'�����z;�纕��-��b�I�U�]�e�_�e��!���iF�����y��cv ��懡#w�'0aH.��ֶ��d5�2�(D�ᐞ!~e��0+��%�g����mX�e�����4���	�M&����q/L��mN��#F�����G4NL ��a��³5��~��U���[��h�Gd7jmA�m�?େ����g�v�tpj�Xdcub��*1O|�BBGGVWy����{���0�uR0�Za����>���'��X��{	!�,��g����uXjJ
�0�m�W�RI`�}��L���s��\��<� �;�;��1�T'�g�`���K�!g�����:������X^���
z!����E'�J�.3����,׹��l���T;'\Q�Y�W$T���+�G @X�Y
����'V�ETb)c�kC�"��xΰ�م:�X�BD�Щ,���!��R�߅�qA�C"����;�5q�>�),lD�Z�\r�������k-V�����Cp�&�s݆Y�_M�7�N�l��$���|	�X5��W'"���&��+���\F��F��.^"�ǯ̇+��<�z2LA�mI�*'b��`2��V�G
Ҽ���?�>$@D~41D��c0iT8�83����g̨gQ�̚���"͐谤k�D�(��(�U�����ў�/O;;�ܺ�T�x�wa��������"���̻�C� �CV$ ?��)Ԭ��|U�woA�-m�I0�!��l����u!e>��Q���x�{�A�����}�� ��}H����4��s���V�l�/L��Ꟁ��t�GVip�V>�S(��<}r�������PbIw;�(W�P��~��J��9�V�F3[x�)Ͷ���*;hRC�RX��h?��WJ3�(CwWQ�{`�T��7�cmWS	�ۜy�j�-EH�w�ߚ�T(+���_���"i�U+D�E'RBtwI���*����*�L�QJSK*;8�VqY\*R�"��X,c7��v8���] qA9q!V-���|Y����g���' �Yt࿄��1"�AV�P�[�<Mw��sV��~{7��P
W�(��oڄz���yyX�������M�w�bql���^AS\Y��3P�aWp#Q�J�c�����wj�e{Йћr�f#�x�o��"����4w�:��BV�_Ta��2?�v�f+`�V� %r�C|(�g�ٔ�3��`���h�1��G�:��(ɐz��uAP��k�ȝg���}�c��N�jh��<4ڬ�GƛV�1�ZYnJ�uޅ��dny�X6��H&�f���݆;��cG�B�؋"�Zk/��Y��8�C���*���Z<?#��D�%JZ�O�d^ϫ�(^�rŘ��(v�oz�6���3�~�Pk]�5y�q ������[�S�L7���B���g�{"θ����3 �R\�~P�lv����/�Pr��v�x*65��:Y5b�<�܊����[�����/Ż��WU7Q�.���2%�WXR�0�ŪG�czQʲU	�{���@|� ;/��z�tV�yF��7�<�F�0�)�jh�xn��!ńм�����ZvT��Ά#[���x�����ʂ"���P���⣃��ߌc��;�Z17��m9j��H�@����&ܵ^OK�iT8|=��si�;��ȦD�v� �lb�Hi�g=���Q�R�9d���'�_�����[C�����$���0VB�d/(LSV�&C�˖��}*;m�]���Ϊ��+\��5y�ۘE{�]џ0�mBjw�z���-5�j�^�	J +���4u|7(QdCL����!�׏C�"� �9H��@�5����]a�1j��U�Bh}��b��%7�6��� ��<V}���f�	I�t���J$c�U:�w�(;5��(���^s�����[N1�m�kmA���$��t3��g!�bc�]��5f:�CB��ՙd���LŢc�1@��?+�(��N��R��1�H[�am��Y=�Y	��<)A�v�����%R�{��O%n�m4'H(�e�kBa�Jg;����fh�@���&:���Q��\o����ϖ9{:<�,`mi(p9�^7�1����caty�*�	��M����8��뤠�����a�@�m!%�U4}{���"^���J��@�5�N��pS
7������LD���C��0�@0fx�2f���2ڠ�B�QE�] �=4>d������*���
8+AհZ���h
l��ۯkh�&�?q�����h�H�Ce&�9h�����Wt����L����.���O�!^��V��l������޶ą�"��@{���!\��<�ݸ�
-% ���7�`���"�$s
��[cȺ�q@��eVH�ǆ�7!��۸#����v�u��t|�R�ybg�؍�WԞǪRYv��?	��)�����q67yG'����d���i����`�$��;h��0~�=�x,x��jQ5$������s(\�-U��/�d��hVh�T�-���ꨉ���%��6z��Co�%YQ�_[������B؍�6?VQG��n���ڧ�'�|��*��a$ǈJ���R�k��1�5ƯǇ�+Ҧ4\��'���+e��x��� ��>U�����8=����g xz�G�;��	�6�'�*�pD�E�Z����"^��X���ފ����<����&Rd��#9��M����n�U��t�f#XV��<Oc��%�R(k���=MOӜ�M� �@�j�cَ�x��@E�Fs�a"�<?r�r���-?�F12r�(��*
��ku�^'�p��FQ?T���?Z�n�5�W�-ԷmC�7���]�8ntC�@=����La�rV��7� �& ����|�6T&��T3|����?��y�e![�u��P�t�8�i�o0�P[��!z���;�y������dNni�B��nK��H1)uxGb��r�Fnx��[�(3�tI���'�F�֐cH����vm�t�mA8��G�,]��W��p0�[�3,#�8bp�~/���u@�A�ɏǜɕA���9RV.R��pU��ՠ�鞝���dlo������`7��9�M��CQ�4�i����	vJ���R���i�$�v�v9S���$��s%,�/;=:�h� 5%7��?J�SR�{C#c�v���"%Y��^��g�R'�eQ��W3��=��A����=2x]�C�N҂dP���;�|K�ƾ�=�SǓ"���켨,I�	�>6��յi5.�5�ș��)aY�=r���<����yH;3��xRϟ��ߺNmKi��KpX^l埆���|�����Vuo[ P�l��~h���ͰY�3��"z�;ӈ�% �]@uV��#��pR��)KO�X#(�`?R5� ��-:��{z6��A�H7'��Q�9�� �����P��r�;QBg��7	�%��.��dG:�*;�%�����ہ3��l2%�������F���zpZ?&�ɨ��������|f�\��T��`T��bQ��+����B�I�yx����5ӳ��,�3K1�$�?�)�m"2L�?����y����9�<-��ث~��ڪ�]�uL���>�]^$̥����/D'��2�w�������i�Nq�y��'��ݰ��f��� �8�UN��f�9.ѫ�q�ը`��c��0���,�R7�,�IkW�v1Ks����k�1�)Ci�{�/f�ؚ,!f��;d.�	�N��xS���z�3e���d	�����
/iHW�v�^���E��Y���I�Zf�f��A�c�����ʸS���W	�$����ưC�� 7~�gX-�7�z�OWO±c,ª�v⛢�h�S�"�j�	�����<Ղ/	������`έ���&+�d_��ϼA/��7�!���M�'�q���s���#�V�n֜ ��
��b�z��g�8�w��:X}ƚ7�;���r�8Pܭ�m�̤T��Q}��_2���Гݟh��j[o�`�.��M_1�e�	�V6�4ܤ�&8���W�Y_zi1����B�M����r��V�f�`P��( �օB�6]�����⃔B���Y��`-��)��r�����D`�RE����SA��8�S�	��^;bόvӶ��W�8���nl9u��\To�[�:�Йo>���������,�J��4l���)F%����,c�(�=A�Z���,-�T�� [�<#~=�3&���b���٣J�d��5�a�ӨG�B]U~	x(D�#-�q9�������G=�7���m#�I6��p�\�M �;�9�W)P�#�_t���Ӗ�J�(n^��X;#�V"����h���	i65Akq���%�I�� �й��O���бv2�):&S0rGؒ�^.Ű�cyz���mhآ�m�y
�U.��2�&�ȄS��k��r߲ �A�%;��Ade��x��PC��P \�}�D_L^�as�A��.�|�IY�(֯��֚L]*11N<X�G���Q*T^y|�{�𝂽�::���	��4`��a5	�k��+�Î`'ݛ=���&ڜ�)k"ik~2�'j�ה����ߩ��T�(��A?Yd4M��?��$(�yIy�M�r��:I?����Lb��S¬}3� �|��؉Z�z����W�S��(3<�4+�}E��i�ް�8�ad�j���p����̳�/�EfC.�j���Wl$j�/X#�e�W_Ǌ����i������*Z�pf5��;$(G�4��`�tx!|N�������ϛ+����e�k�L�bNa)Z�O>��2z���^ Ĺ���f,lҨJ�4��m�"���+�����p�UlCY�@ĳ,��IWy�R���?#�а?n�w'�]��5/�����
�����?�,�e��7��o��6R���kl3��z��r��!ޓ
8b��N�� �Út�	a9��OK��5�H�D�vB�GM��� �a5�w$���Q�n��������H��Ag��iL�-
~��0y�Hv�"!)�p���j誣8 tXgy����u�^�U?��j�#���d�o<��ª���6���T،��)��9��P��MF{�� sK7#�<nlj9sL2����oϝ���WgBwBK�a�X�)~8N��;#Y��o"���j��I������6��v�Ik��kg��ڹ���B�Q��AcXV(��n�]R"�Uڸw>:7���3z�[zoܤ���"}�t�87����+����iɓ?�*'����!~E.���L#�ET�Ur����	�풑��Uh�gZ�Y���"1�ohB�nђ� �pB�Ǐ|9��G71�,;�ԡLz1���NL�(�'���F"5ؔ�ϝ�"�A�P�H}݇�1U?�gQg��蛼�a��Q B��+����7j�n�|؝�t���&��8��!+AWC����P!�$8
O6���4���[}yD=���i�w�^7���Pswg��R��h�*�������ꇽ��U�����j�hSR?�n�=K4r�M؋��vx�I;B�E;R:�~�ӫ~Lf�BU��3+c����Q�h}]�X0ԛ;��=ڂ���p
vh)�hn���� x�#�1kG��Qt�u�Q1��i���[t�2&H����������d�x���B���z�(�w�2[V��]a���V�5�+�l����4�@��1�࢜'�ó� ��C�Xn�z/��10"�F��lA/��k[��{�<��TG�?f��@�+b����>���[���>Ca�,���^���>���B�#Pl�{��M��F)���3k�w/�3F�ϓ��^��X@�%��b��ک���{d����y�3
�2�|8W�J|D���#:�ѧ�z;�z�K�Ɍ�G�2���+B�O%�����Y���y>�ٍGL�h��+"d8=b�h�PW�s�7V·;�E5���0���l�rH�t���^S��s���JXfP�MG�¦�ԝ�^+�n")��3y��B�}�̮]�0H��4�,[*�f��EiӞG)���C������� ~�yG�^�<�1��[=:��iw�d.���a�t���{�>�c<$Ă2ؘ\t�f�߶a�m@`xLT�J08M��7�mxr��u�"�4Y�cq2��yq=B��#9b�h��x��	��(�Ͼ�dqη=F+h���P]�v�m��H�sΉ���y�U����)d��S��a��vp���,乖�0Zࢌ�n;+٫����P�'��0�����)G�	�T�q7d����b4`�b ��{��������QQp$�nc�5N/JꝎx��0"�H��V`0�*r\���q��K����GV�F=�	e��K��Yݣ'��a�G +8�	[>妚�Ve-e����o�A�k������>��a^��'��w��ˌ@���g���כ�桍4�g�(�4)$�UI��kd�I�^�(��q6`��kD(��Μ��"��ZZ*	)ձ$+.��&��:�螠Q.�;09\��<�c,m�eKcL�;��,	�省�* a�����>�d�+��F��8@vm��͔��ݦ�+�w���7���Hx�����{d��
��'0����+�g�<I���G�ԙh`&�,�mxϴ����V�=��j2�V؀�����Sa@?/^wD�7?�2�y�����!��br?�������qQ.JH���.��O��O��48���� ��Z-캯��M:����;�h2��J�9�=�.�l��4���ga�뺠R�˼c�N9�!��e�>D���R�=����8���ܦT��Ǟ��U��ѣ�|�f����F���鎳���>�Uӡޓq�J8�R6T��O�o�b܆��[�g�j�u��;���	]�Cw��?юY�G��,k�\#L�����h{ʩ���%`��6�c���21�I`�n�����u9j;WN6���}�h��7.��Zy�j6��Y�{��k�,��k���z��?l���;[Ē
{W�j��a��<LB�]�R������В��L���#��/w�{�1�@7&`�S�]�`_7W)�n�\� �-L���,h��VP^7߅�&�Q@I�aY��C&���|��0�I�P���3//e*��K#G�����.t2�=�*D��� �HxлT��K��[41�";��4RW�eZ��Nr�܌� ������1_P��-KR\����!�3�g�l&m��O�]��\���lꚂ�4���F`��r_)�b�լ,�P�O22�t���f�w��������Qn@�~��0<>bh?�+�4$�\!A�
n3/�����ۡ��%,���a8���R������#����.�~��㔦�� �n�M���!U��{xOi�\ӐGkfe�$M7�m 2�l�9���%�/3\Sd��}H}6�Ua�u��͞�JK|�x��v�S0����0�B�O^�V��`ށWa��B��H�i�42���!ܺ�f5�R��=���cXS�S�ׁ�/� ���o ���&�݁~q�ۛ�=-�Na[j��Y����h�v���SF�l���E���|g�*��''�����#����P��]��i;�!ܪ)���r5az�=Z8z��F�y8ou�)I����wf$j�����j���wF�w�f��o�f�� �F����� �c�� ,�#�R��|S�r�"!�j'/0�il[�8vg��ߢ�\�-���9p*�:�D�+��Э��Pk��S�q�T���dg�/JԎ@9����۱]G�����fv�lp��u]�?��7r�c���w��2[�6�t�U9A��X4���JDk����F$'ND3�#M�麷1܋l�ύ\b�|��d ���ܯ�P�?�� $ʅѿRa5�֭y��I`N���2���0��Iu�q£F�saLu���ֵghg�U��)�5QQ���-L���\<�^<n�z{�(�%��-���n��H˪T�S�ouǍaf��_��?�� ��v}�q;��Қ��^�y��Cnr���T�q֮��on׉��+v���,�
~Ϫ ��ī�"{��b�3?��	)ŲDحm��I�x��k.�i��]F�?C,E����Ӹ�R�>K+ @M��H�|�-t�����y"'�_W/���Tr��c�%��5�o� �j����(�n	�r�睹ي�P��N�Nޤ�>�Y��u�q�C:�K�2�_ܬ��5<�0�AI��w������IoZv[*?Aӳ�Ԟ�[�B����;���Y[��/��eIE�Zu�3��촁w�՘�e��}�ԎF�$�v��Lk�#��U@���P2���S�؏e!����ʐ�?��t�Z����=6�4 ��K�V��B-��D�e�s��u <�g_N wRk���y,�t�X�D{��o��\�(��®U����r�
v�3��W�k���{�y���6��w�] m�>ҫ�G�
�[f�������U�p�5�ڥ
fb�l���Tw��a��Unp�
S%�GDE�r+��%�^��5�j��/�	L�{��)��(ܜ�E|�s�	yȭ~�V�^v)�7��e�S�V��
�C��txaA=@Í�������^N�q��ȿ��ky���&Kr,�KT$,��:~�<�I�L�:t���4O}|X�H�˶y��4���K.�Ґ��㣯d�oXqt��n�T�L.4��Is��T�����>�`�w�h7��hA��p���S�&|�7=�e\2�MW�.hM��V\���5+�Qn�׺}\������Ř�3���)�HCS�k��7k�j3�Ɋ?𩌄��O�Pyj�S�fW��?Q�}=B��q���^�����Ӄ��>�,�8c��x'��u��i��׃LY�o`����N�]t�ڹC��w.8	؊'9.�95t����P�k5+�'M�},����#�3�Ŵ�0@,�R�_���#�q\�M Y�a�+=���� @"�ARЃ$�HNa��C� tt����R��T3�z�u�����+�\�9��s�����E<?E���5Щ��ߞ�b/�Zِ�Z���0�ɑ.ݖ�8�2�̿1=!�< Sӄ%Q�w����p�ҡ_Cp���Gּ6S��N��K��}�v��I�*�y.J����N�b��0g��N��e̺����T5�U������~����ө�X����~��G�'�q�8�t�H�뮍�Q"�c����5!z�X|�R���&�'K��R�o�������V�]� 7�׭�S(��~�掱���W�[�2�ģ�}줅[o�	n�3���� �0�xn�5�]��;W���OR(c�y.�1��m�Q}�Rzr6e�66�j����
�f�r��d�M���K����ǚ���ͫ�<���R�z�S�f�]�A`RH'lj����V�,#Ӑ�!c|bBsx{e��.�(6e�Z�6��+n>�H��U&��g�c�+j����-��R�n�L�Š�o��������̑�Yb0-�Oѝl�Z"�*:*#�H��U��aeq�$����s�>�t��mٷ�8�B�G�,��GC�g���Jl�F��m�Ʌmaq��hG�.�W��<Ao0�H$`�}5FR���U28Ηs�%�^w/T���Su�!��;��/NnW����6�9r��,�z|҄�*�'ð�F9��42��[��[i֤E�J'��0~(����VNpԏ���=V�e�=r�t�S*e����.̵�r�&:��pV��è-D(��)��>dkgS�V�n�,���x�aхDu(�Ztv��E�[;d��>n�9K�3X)6�m���y�r��-|;=>A_!�E����%�q2���c�!h��~�c\:F��sa��(�[��R�|�Po��jΔ�4s:�Y����>�k����^ q�[|	Rά����.mԂ�$�C8_i��G����� IEƨ�����e	b0���Ff��x�I�g�0�L>�����#S�3^E��M�4���
p)骡��;� g���X��{V�ܽ�4�?l[��˓K�kt3�d�G��Gg�#cb΅�'��v:L�iM�^Ԡ̡Kx�K��l:�y<��[<|i�Ekx���x�f�>�}�����Fug���=c��٥~���Am�D�䭧R�/���Vݹ�x`!7/ʞ��kB
�Ll����U�Hf��M7���������0u;�"O�����gu����/�FZ��;C@������g��y^��Ɏ��#x~Q�� �K��T$fn��I����7.�PN���}�C����<\��>.�y�ɕc�n�pJO5B�LY���j�(��5�y��\E�c��^'�I�J�C%���'�^eJ�>2K�$�o:����"�xICy����R����ӓ�=N8t��I�@�9�*��v��@v3N�	O���i/�V�����ku|ٜV�	����u!s���W�6�FZ5�D�7���g2s#I�:$tP/�F4fn��ˏ��p T��J�=��;�fӍ[��N�	�{!R\�Q���� ��۞.βw�	��Ky~��'��)���B�SD�ʒ��A��)�Ak꘢j���e{ȃ
�"�"�3�C�!n�c.��/N��0xJ
������!��M���M�*o�cN����t�	�����k�^)V!ܪ����M���2d��k��
������'9��Ƃ3��Zjd��?`��4����8�q�KA�����-h>�lr�V�g|�K]?3�+W���`I�q��]0
�=ݱ��� ��M~^SY��h�e�xn�U��X��Lb�w��"^`�<vR}b6Vȭ�L����x�P�N�p��,_��^�T�h?�>�K�_���a�jضi9]kv_@`�l�*n�Վ��ڱ��v�RX������"'6��;���V�>(�=�� a�����h���lq���@ʕ����\I�μ�,��@���5x�k�M��庈���A;��cb뽲3�YU�X���c8c��a��B}u��+pM4!����sE���!b���o�w���0��!D9�k�'��@�``��1o{�`���� �Wڟ���&��L��w��g�|M�����Y�*ˀ�d��Z�>��CD�F ��� �=�1�*w�6����Xd��tR<u��(Q��L	Va�!�����4nz�8LB��&�[Q�KJ{�2��jg����[��Ҧ7�d%��p�����8:����9[y����1�Mtf�6��V4}��× <0(h�����x5$<t�ߥ���MǱ3��Ck� ��O�:ݙ[�2�2�Q�!�~�g�*@��Y�3`��cSLi@wō_�ĵ:"� �9���4s�Ϋt�n�RX�<11��a�q�$�r+�_����ę3��q�����חy;N����\�u���LrAu�����uV�Dgx���y��I���@�֦����yʨR���T��{z!g�Ο�}����!f��	�,���.�V�]�O= pxB� �X�/(�΋�cΧ�x��d�����?��r+>��ڮ8� �������r��Ñ�T!�1�e>����	r:�w�%o���/�
	Pg�
$5y��]2���"�=}��F��U�P�6ѽe�_�Ҵ�l�p�w���:*�;wn��俦G(ҹ�F8��6�
��͌|�V�8�]���X��i�%'�0��
����{�7A�Ĕ�~m
�l�ˉm�@������32K(y|�o����f����ji�q%�&4�#�=|j�*��k��p��ˣ$��̘�"S��;.�� �b�S"'��3�̀�\������SF�Ű����Z���{��R��#X"����S �?�M�DV��e�-��������>9��Ff���y`�����Ml�>����┇�.&��|��f�������4����+:�2�z�D������ڨǨdt7K@�L>IȷA!��rAр���/����h0�@�|X���5(׃�7ć���fp%���b	m���_������Cg�A|��9�܅��r?���*i3vڟ�A�!�<�Y���lf�1A-���/P��eb��f]4� ��G^�D\ĬˬcÂ/���4�)�c��I�Y�=l���}kXb�l� ?�����7�E-�&�l&uGρA-�UI���)�lf�X�6�w����ZΧN}ֆi���t�?߰�8-6e����./Td�
�0x�{�kߺ_|����6@�т��jӅ������mC��,\=�h�ȈB*-����nŎt���\�ԅ���Y�5��ٟd*<��;a�;��]OX�k��H
����QD��:nӵ��h߷�W�gK�G���ֽ�vw�I.ّY]t��p���װr��z�����B)d 3BJϪB09�ra ?��ϔ+�&�"Rx?�܈��H��r��-iMf��!��6�����J�J�C��|�b�������^.O�
$�,<$��s�2��)��|&�co�&�Hj�z)D%�N=��O�z�'{��=m�?1f�r޵�� ��'�y����Ҧ���CMMq*�X2M4�v�#�08��^�	��ݔ鐂�����·����-�l�z���V�h)�fY,Z�Ǔg㱶���ƈ́�{�{�Q]D���tK��������Ҙ�^�����I����:=�j�Khu���.�7�2�$�%?��kY�]��>L�jj���o d�/8ؒ@�,:�4:��W�yx��w$���2K�q�d��fm���������k��в`��4��B�/ˊ�1���lOg�a�a�t"̍#i��sP���U�߂��﫸-0�o���(0�ڒU�[N���9$]���U���9� ��K\�-�S�z�d��۶���@i�;���a	�%����׷�����LLR7�X�y������$�G���y<����D����J����j�2��E�J\wR���9��q���(Q��ϯ�Q�2Bw@�KY���J��Ʀ��h-ѥ���+��0�5��u�̻���U�zEt��ʜ�ZgZT���E�Akm������j�u_��!6r��Q�/���L�5YR-�0(�85�Q�d�^��w��c��f]6@6NЅ޿Xseς{m��W89vcY����6����;�^7t�4C���B��8Z�wC�ɓ�XdNDcO�f����s�Jit�$� ���"X��z�eÝK�a��%!����_�uyw����UM�� J)]��j/��l'�������Ǜ�zq�S��tF[��ѦZ��8�S�\L_,u�����H��r-\#q�?�=R@���zC��_��l�I�B�[	���qq��NV�����lm�4��"�q=��K0qU��@��cg$;2,�5���7O3�������@�+f���/��|�X��ͦ�O!� T ~����5�������j��u��c�Ǆ��ɔ浤r �,d�&e$�$O���q�����:W�;~��%��ն�^e*gL'QT�	�g�c9am���ĊM�:��[6w�:���V%�Fr) ���R���}`�c��ç����&J��~��-W�^������k$A�ZO��5&��H��wkY�^��;Ap�Q�ΐ��_o�!����0W��ϧY��J
�Uf$U�R\�)��=�K��Gx_@�P�s�ӆ��*:=�4A�:��I���������[.D+��@�Y�����BJA�(eO���w�<u��e�Ԟ��Rz�i+kl:�Ϯ����Q��t{ై�V�3>G��ki�3�g'vA�| 2��<�1
��~ş0jor11� �h�c�Z�~����!H�()��p�Êgvg�I��n��l��?��F��� )JD®��V�X�[�(!X�Y8>N��u�]���}��yOJA��L)�(��׸��@�g�}��9b8F�&�*f%�w��Eg���޲<�S;Qm@���9a���S��@K��6[�����sg喽B�\�x��zbJ2�WX�1;��3����;ܥ���X���~�B���@жv�z�(�Y[���x���G|�Y2fX8���f�l�_o���4�ea:l��g��y��)�	cwЩ{x>���	D�+=�j�v�1V�RuAplm���HL𲉓Y���?Bߚ�%�pۣ����Y4�_���	�{O'�k�k�U����\�r�K�X?[M��Ю*i?U�h ��`]ܑ���Rp�om}�(�1�l��\cI����fP_#��C3�b#��!7�#i���z�|��t���C:\��c��b(��G����[��g��=���B`���O[·V�[�4F���5Ή���ï�3�cj|_S#K\��T}�W�����m����L��Dcs��ĵ���ȹ����{�\;��
8
���l9���B5'��+�]3+.K�ۓ������<���q�L;����fm�x�}5�k|"�V?չ�x,�h�}]��:��	1���9Ő��̺H,8,�}*j?5��D8�C��V&�'���P����|D3�@f�â�D�����u��5��@�v<�>bV�|lh���նDS7D���<ms�I��I�EsIֈ�)k���u|�y�|a)= ��V�[�3:I'��]�h�^�A�cw%\4���3�����4`�e^��_�6���TA��/��(U�W�ɡ��&r�4qG��h�) ��1��|�z��$��_U�:Q�ڴ�iSH@P��Dz{g0���a���5�w&>T$5{�B��ɫ�.�$���!�ܔ����2L��%fm�k	;	��%_{���3ƃ������Qn6��Ε�"g�@���K]���E��
Iנ۝7C\}�+Dl������4BB?����).gt<tCFVB�g�=0VI�G��#Y Gi�ZbM��@�",�+�)G�)S�p�;��?���tT���e~�,�z�u���r5�/�oEb�Dy�Z�C�}Ƥ~X
����ͥ�&k���>�:4��(R���(��{"��xDԟ5l���n(Z�-+�'���x�^ZI#��t��2�X�_.X;tR�{J�� h��AW�A�Qf<�F�|�l��SŔ�R���)zj�J�����e��7���qz[,�W�9�Eo2��'`��̄��?#��&��;U^?T;�΃*�
n�k�Z�L(�"���kL�ЄP���ة3>���"
��ܳ�k}E $	�Co!�h�|�0�djlӟi�O��h���_��}YW��Y��+��|F���/��)�
��тZ%���f1�ؤ��Ƽ�7>3��ռ�q&{T�Ghqo�N\��
�j��C� �!�Zz��h�Þ���k�G�Ϣ?�'GЄ����p�ޘ9���j�U�dmY�f�Nj§������l���l�q����k_���Q���L��Qu'����Hd�anPv�f�$��H2����S�������5|��T��8��hPokx���P�aD+�n��q)�{��BkF���v|�6;Q���H��"�^�t��MQŴ�#�\g�~�ٞ7�c��������է�/3���?a����c֬���:T��{�1���R8yd�V��"tL��'�,��"�fvV/��VA������-IS(o0���XCb�'���Ka_�4�����+��/�7C���Mɭ.%�s��)e#J�q�ņ����z��84�!�M�`�F^��y�uh<$�H��Ʌض�b�uR�ejE�+��ԇ����c�t���!	"$D:$8��dѦ�^l1
*�� ���NW��?��TF������$t��E,�R&58��L��!pUt�y�^ р�h�-����������(4���У�u���_���f�\=&��ObLi*R <���l]��]��?p�E^u��I��k�t���\@�􊔷_Z��}��oڊ�{+fR�L7��%G���	�k���Ȗ4u�������d�-�x��x�k���쥤��#\7^�`�� c<h���5o<�l+�{���2Џ��U1ppE&������5�.����`��x�лLnz�u��$����H+].�-FV���W����WY�a�w(���DSdۛQ���x+��֣e|ip��z��:Z&I��ri�4=Ԧ���7#��/�+T�,�'��0:t�B[������E��P�I\��'�yJ��rKugk}�w��WY�Q�N�bdW쨿蔈b"�?~W_��/WG��.M����c�ZKI�o�Wy1�n_6JP��#��Ih9m�zt�/�0T��j����cO�)5B3�!�)M>��8��d���	����c>�� ,��L�)��$�P�L9q���l;G�3���~ڛګ	u�+6N��#�|�5�Fr�K�k�5���4�N5JR��v����l��W��� Q��<���+x1�uQfϯ��I���8\QSrtu���w���¶�ٽi��_H�6�Hќ�=fSm[a������9UM��d+��+�`J,� [��m�<�4e�R�bD��1���&_���k�#.m���+R��+2x"M䐄�ƐP����5�i��jO��r�2óAm0E
'&vB q�q-�7w��B��K����j�2�<c&� ��2���ǀ��D	��[oN�d����g���$�w?|T�Kk�[�ݭ'r�����)_��T�)4�)$�OL������4n-�%�yĨ�ش��@�
`^7/�g�-��V�ڀI���Y��u*���pU����)gD1�Έ�W%j~:@P���Ɵ�u�x�;�[�#�^.��L��mkMV�?̭��'^��U?R��]���S<�?d񦜠���V2dU_тД�HF�I�j �K!u�S�LƋ��#�^1>�|�].#��6oܲ4\8wٍ=���\����ҹ��xJL4X��ʚ�[�LU9v��m2
^F"�g]K�D�o�*Oc/$S����(�v�4�
?D�`dzZ�%�g*.n]Vy�wy�[��@�Q��f(�t�H���QaHC�WnLvv�S
�c��
��M���9�X d�j:�J��'��W����W�U���27�*��:�/�m����=�䰪�u��"��#NKc�Np7>����A%�"J ��v��=�I\���%�ڹ�����,5��g
_�0�D���O-��r���1c���l�'��r]��ճ|yt�MQ�]�w�֎�'����b�x�8Ny��Di���M�b՘��}���o
5��u�vTxgf+���LklԿx_��B?M���6p��`�D�Q�ю��E*��<oz4�/6>L��'�ٌ,*E��/?���[p�g$TP�۪�i���&��U�Rc��`%��X�(���.1�J9����?��9[�ОC��"'F� �(�2��Q��\7ܱ	���3��@06]o"�e��[�?#.[&�wVy;`����^Wx0���*yn��xb�/|H���6;חO��S�ࢳ�8�w�0��%v�׎�ggu�gN�Ux)muM�Q@b��'�����R���5T��{���T'&x4�;{���N������tE����M�1���x���"Z�����V���{��j�♝���MQR�@�/�s�Dh��sW��-Z��ٱ�V'l
ʰ�B{�!��?�uN�8o���ܢY�E��K�?�����um@���1���{W�&�M��9?C� %H��O�XR��Q���uq4f	��-gu#$��pr	]��Y i� org
�m%Y�wS�y��qt���#����<���Y�*��M1�$���[y|�,��^I���]N?d���8^�=������o�nE��ȝ���$��C~�FGgo���1ȅ|�O�j�O���&��-#U�֥<@"B.J� ǝ�}ed�k����6�:\Xu�#���J��i��SK��(����x���R�&=�p`kV�db�ι�\�
���a:zvrc�}���r�.L��Ngw�D� �I�eNԄE{�d��Eͯ9O*O�	�֋2��-gP�woCe�uȂD�7��4��6}���ǹ��x]�jU�t2�ҵE�LV����/��T�!��W,hc�F7l'/�@��F��*I4Y��@u�"YO�6�,:�I?�Q�uh^�)�Cq����Bӧ�����Q��]�	�[l��b�ΟT0"�.�bx����%*���4�$��������xll��gn�9��|� ���50���f�Ӯ�f�����1���T����R�f��"�8�~�[- ��sqv*���2' �ݑ~b/X�7�wbxպ( ېM#2f�鵐�1��h_*jt6`��\]��_ �|�[�߱dAHQ�o��'�E��ܫ�<�z��X��%�a�LV���]���0�Ib|�J��Y	�	v�7����-j���MrgNM����&mЈ��`�qݠ\?Ep�*:d;*�n�8��;��y3�	!������~��ۡ�=6��J�#��D�.�?��RT�[��pY�ߧ{HL?>nGg��ɳS0���f\1�2@�doo3h�ة�+�ME
*�ۋT���2�ɧ	z�+����L����ODT�Z�3���6mEIQ��۠�LI�7Cˆ�@��QI/�Һ!�:�'����|�Ѿo������O-�jm�[a����q�8g=VT�%��䘟G}w�+�t������A�4�v6���K&�@����2;d�2=��vlL��s_N�ٝwg�5�4@>t�6l<Ė���g��H�#dgB�N�ԑQ�g`˳�h.w��O.:��9W��f�ڊ������e4�"��:��^�Z�x�����)p��˕�,T�X��s�V�B�����$K�_Z��ȼ]2)PYA�=DpY�U��XDXU����w,7�" p�5w�fI�]ީL�ߒS��tf �x@�K0>��� I��mx=Э ��sB3SŌP�����O�v�8��[I'eC2�z���G����pذ��6RS����֠�@^�9ݑl� @�9���5�BG�/�rTU����>@B���*�ݍh��}}�[c<lc�-��`�v`���'0���wMt���bm}/�tn|�W&�62W2�k�t��"{��5�ᘋYN��Z ,w� B} ��f�n4-FW$\�����P�hC`�D��d�D��9����vpdYG>k�,��%.��j��5ٮ(j��Ķ��h0�D��S��6��8�%�n�C�4*O���a����jj��<�1x >nՁ�Q?V���ei��RO޷��#���_���2g)����T?�pb�d]5�5 �,hѲ��~�ɟW�W�|�T!��0�s��T��h|�9H'��������!$�TfE�����v��_�p}5j���C��J"Iz�[�i茏4�	�0�}�DnR_Y���a�KnK��ŅoK~�[׌J�����8�W��e2?C	-��n��������]�������2�4b����Y����I��X%�>0S/ߞ�|����}2J�e�����7-N e.�Kc� T��j�d!��m�!��w�Բl���W��Z�+>)@{B�������ѶXb��׉?���]I)r��ס��_Qf+����yq�O�2�;P���w�[�J���͔R�y��'Y{��`�y�?��BT�)4���d;MZ_�]��L��0�C��iRW�l>�YW���݊=\�Q$~"4������1]��jsb���
+W@�T.�5���/U0�'O�O�T��Gʀ��v�^�r m��N�b��yقy�
W�������B���H�d���z�&O��6tK(��lS��6L���
C]������y%�p��x���S�<+�F��-5��!�\�އ�v���3r�f�ͦ�/S>�+f�}��a����󙔖��E~�7���ӸNN��~�d�pM�BWdT%��V�J�h�1�b����PUn,� t���+W[6����Ɓ���l���V��\J����y���K��;,��W�!S�3 �?���cP~�ښ��z�`2�5Չ����4ЬY���v�k;3�k(𽝊6L&�0�8��Q�	 ^sʋ�zYW�d͔@�� ]e��&9���l�~p�r1�3wO\�3�h�ۧ�)�rq�ƗnA���P���KΜw���5�%VE��'����i�҂���R�N�|g�lv�]�Tu�2L�+$t�^�:��c8����O0z�	�6� ��o�l0gp���c�����y��3��Y���K��J<1 hZ��'�JI��gK)�y�����T�f�I��N,�l�0��G��#���c�<�u�U��J+��^<�`/.̬hl)���eyv3�Z�����z���"1�ġ��5Q�@��2�\.s�J�w��e܅�i����4G̓��N@�SKxxlb���r��E�@��_�^��w.f�\S��od�I�)_��e�z�(��[���Z�4�	�
 :��L-&f�{�O�SVy"_��8`?�h�[(�FL�hغ��0�������)m֦�|�r^�43��E,a<�A�w�o�R�L.5��:M�2�g
ۀ����R�}�mp�?��bc^bOұ�DrN�7���Ʃj�>d���ݹ:1t�|�Q�Ñ��"�$��e c�A�S�6[/Ӧ ;����(�cG�|��	��ˏ�ž�andk6���B����L��������e4 ��%q%�q�釰��Ha�x�-�z�>𥱞�a�zN%h)����dr�7����<��/�]�� TǼ��k3��v@�v�J��W�Fj�&�����Q>�U�>*�BQw��Zk<ԭ`���	S�o�@On|w<����7@�#�t�]k�sm��W���̺��N��rd��U����f{/�fKR�)������U�N}�2[��us�L�K�{�W�ߨ9�_���c��e�� {9���L�IC碣��]5L�����pf�g�Gd�}nW�Q�E�w�c�jvgX����E��Q+�I���7A�!QL{�Z�-��91C�`�>��:W��y�m��\���B�@�<�EJ�|��;��w��`���ͫ�ʺ�VI3<�p�nkS�sC�-�da:\�������e�]�� ���K�h��m��{�)ˏ��dt���x��UYQkQL��_���k�!�����z��p�uQ���`��]�o���9sJ��ǰ�����	s��f�9�`Z�b��n|��/�u����P�̾q�=sДn;L��Ŵ[M����Ͳ�!��ae'J�}^�Y����J��-��C�c����7�����Q�(~Qu�ho��4�����F8�j��Myj�<e��:�:�#',}��M�ƈF�/�k �����4��L2s­Ð�4`�$7�����~P~*��Y=�ٱ��'u*.�~��yس�%O����R�ojm�d���A:�jd�tX�f�*G���>�*|�C���j��,����7��<��K�z ��t�C�(�(*WK���(��S��\΍#i�����܊����a�uД�-3AD�X�*k��f��Z-��
�M���#x�Q�JPLq7X�J(#���}�y�pU�J"	3t��9<a$�@e	���;�,o��#_���>��>WG0���l�Ȇ����*K�kL���/h���&����U�&��v>,x��3�O�%;���M��+9U����|��J��G[���?[\O�yx:u{��������A����aGBg����wS��
�=�C�fӇ��e=���Cɷ8�����E���?K�~6�T����y��0�~ �x�7��������z�3�.���9p�Eh�ǣ�\b)i_)5�@�	��n�@���=
�$y/�?�ς�F#�!�|B3͌cAC�͓�3���Ă���)�ơ?�l��(�,�xZ��)2d�����x���H78-�0p	��6آS�A#�r�5K��y����
�ؙz`J) w@���;o�x8ǝ�lڟ �N��p�-��r�E�iÉ���	l�{���.�n����dN�oC�[�m� 1)����~�����I{����ϧA�\B�K�<ӚT�ka3hEU�b�<�)C��֦��j14_�Y�Fz�Ơ���<�TE���9�@ �1�K=���ʔ#iSy����.S�Hx���	U}��Z�KX�0��5Ry˭,�@s,�Ù4��,�1�V��x9�5a��Rc[4x�/'-�ބ[7���
�*({6��;�%����Ob�����П {��L"k�J<(��_�I��S6�^���������L/0ɡ?�r3�#U+>Y����˿��^����
�T��7Ǒ}?]6
w�����jr7��$y��R��[;>���J�����}�C{� bR��|���%�VLq��?+V�3lK��|S�0n9�Ie4.���[�$�Zb-�j=Jl�2�W�ja��1���x*��}�$�Ƕ�q�H�P�qg37��5��Y�j�*�N?E�K��/�.�h�=>�F�!�`�t蕎���z��u�Sf'��ބ����|:Dο)��ڌG� =e�		�I���)k�죇���X�|9q}����1�!�1��	�zR�l0��W�͟(s.�	���N�l�R�4�Y�Џ��y"N�s+-�[����p�Ĕ�9��C��Ypx:"�g7���l#�Ne�����!Y�XB3��2�an�a'��E]G������:��ɯ�Y\M�2�n����|�S扸0�)�v���H�MӊI�E�79��G^+��0_���ͭm-'��-a�Ni��vG�O�=6�äm�W��H֯��Da����Y�E�M�����C?�js�1� 5P�K);G�	�Þ+�1`�d=&�&pͨ�X��a��΅��XݾX��K��`���N�$ް��X��������[vf�[��"�P�h����]Pi�E� ��{^B���\�IW_ͺ�o6�c=�S�rlS��1+�)��a��A%�)B���m��ys����q�Uo)1u�+��9�ʉЛ`��:���v�-[�l;.Lj��M���������f,���E���M� ��O��� ��4_e9�Ysr���
?P�s8�+ɡ�]E�to�	N݄Ok�� �����P�j(�3�λsC��ܑ����~�'	�a?#K�e�yvF��������Bl�6�Ո:�/1Z�U��K�.U�f���q2�L��d��]ݞ��J�3�xt�Ji܉�h��IK��@�5�Vub��|&0T� +���t��)a�u�]�|H�=jt2���ˬ�"�n}|.$����,�RY��j7�=���IeDI���l&�!"�sGө��]m��ULa�; ��M�d4ŞX����P-�cJE��bJ�Ih�˙.����ـ�ن,���qk��H�ǀ,R/
Q�X6"Vq�x}�ˀB���� w�4�����ۭ�9���>��e�S��^���S�D��%��福_�$���(DVl�K�y��bl^�(}y���2gOFB4{-��;F�X1�L�\wo�$8�����["²ղMKnW[x4�>6���z?����棭�ު���oT��2�@���F�E�(��{�g}tN�e�{�E��Q�\M����͠ˈ�5������D<��+�.��'�������	�زS��ģ��)�q�<(Ե�
�ð�����D=��zo:�D���{��*S��[�ٴ��t>uI�/5I?��e���gљZ_��оv2-�{w���珸
�Ky�w��~6���߷�j�=���H��"����q��R\	�G[��!����^3XA0��F����M^w�>AZR��](ư�I{w>\�e<d���4�w����[���!��S�К��?� �K�&�xK�o@s�+�	�Z�,.Q�����^P!���:mV��n����0���~����#��o���������#.��e�ۊ��ى����A�51|��[�φ�W0MR�D�
�&˘W����w$�J���*@N6�=�'��D����!�؂#�E��9P�ׅ��<̶�/f%=:G��|�R��fZ2�l>�IuuZt����h�ϥ��9*��0p� _A�i�Z�N��jc<�W���ҙ��y}�Z1Ǿ6���Sk+`���'���'���NHl0�T�%��_�����9�N�4x�"!s���,ɞ,�ʺ���~߂���mF:�,mp�@�,4�������R��������p�:H�pՏ�o:�Q�A<◥Z���x0���;�E~��Kݥ`W�g�J���H�Z���׷�%]Ǭ`��޹�����xm����x;a1??%ٚK�X���wW9�T�/6�KW���C/�Z�2��������eK��R)�;}���g�=���A?Vž���
�E�^@��Qc����[}K\.��a�m�_�blx]�a*\�v|�pE���i_��F�59��M�ͅ�����|��2C��t=b��_EvD���6a+����!`��?E��Y���u����e��Y�A'�ݧ���\yF�X���?"��Og	� l�J�Y�}L�+<�-r����=ҰfUZF�ɻ$�nL7���]��zo1�7֭�BU�\��<��� �2�t�OC�3%�g��Z棐��bF��"�ڝ(�)�հ�xq�.0r��Ҧ���ɣ_�?��F���f34��ȏS 5[EӐX����-1N�}��Wg�["�i���@Ȫ��zj\#�������rf#'��W��r�J�iV˹X�j��|U�[t�o�8Dv�$U݇�r@�&&݉���4���O=EV� C��<�t�6�,�x����p���I�T��hN�s#j��]�� u�H���n�X��1��TOd����&�Y�56����HV���.�I'����;�feuy^�O[��ᕉsTfI~�;��Dl�dWbj���t9��hx��V�������41��ȯ0o���Rhf:�kηNk���!N���g.�W;ݚUr1�Zɩ�
1�ή_@�����+��vv�[�]�:�.������]zd�O�2�(���qB��
���tӊ�b�R?`��7W�k���<��:���\��U�^���I�>���@h��r�:��	��s!�@���'^s����G&�2'���PL�e��u�\CZ'Zw���gѯ��l��m�7	7��tl'����@{Uzc����<zI��%�r��t`C�!���g+�o�Z��c[��޺���%�$��e)���٬��f��pY��+]��p���{f�W����&��P(.܍Ɣ;tF�K�1���r?��(O?J��+�0��	���j;)�Q;�{�!%�3�r�%��}U������ȃw��l� ����,
 �U�@��a��J=�*��_�����'�U����vE��Տa;���F���W�nU;�+�%5v,>mR���Bk��&�t*��)�����Ef��ї�ETs��Hs����n�S��Q~��ړ�VD{��h������ ���ܚȸvq�_�4�=�����n1�;�Tc�k̽w�۾@�&��Q�q�2�f!I���hɁ7�g���<���z\���6��)�~��k+���8ҧ�ep�Mӽs�d����X�S6�����vH�p��Ξ`�<�"�h��ZK��cj���Ǽ&CD΂�KU�	*�[S�&#��
ʉ��p�P<�R�>��޿J�:
B�)�0)o"1��	��B�6�'�~�RV��Ob#�9�(y2�G�D1��e-�iHD3 ��!@�I=�/A��� �2�c��A$��'�C���Q?m2�>��ۘ��&��L���]�����/��נ���i�0�֞.؆��wOҝW42�_m%!��(���*^� مw���5�\b�����K��y,SOn��|��eX���z>��휭:�ͽ�U��� �.?W����䗜��u�-x淯b|@���R�z(����%Č|�R�L֒u������Y�a�i:m��
��&�:0�a>8T���\�w_�w���a��� ��i�[�t8
-g�I�֭��T�j�� �(r�������o�-&��H����ےS�,I	t�w���o�<ʥr�l���se��Y����
wC�:�^n�Q����e+�A���ol�񞦋V��cZ��OUb��LD��Yp��(�WD�uH@wiu��=CU���6$;���Z��qi0}��ì���� 4����b�n�r$c=���!_7THo/�@"�x�\$�'̺���Lj�!��跬�g�-[�a����Ҋ��8�U����k�S��T)�,�{�sP{��o�+q���i�s�k�|�-Ú�_��,��7����3���p��b�J+92��=�k$'�fm���I��˳��:7�e.Epڑ�m�X/
�C�&r�~\��Ҏ�t >F毈OO�֔@��aK��U/r��M�;�eթD��R���F�q(p�(�l�YL��8�a�z���jK��_�u�oT�*qzU���|��џ%)I��.�� j�n])
9@����d�,��H]��x��u��5X�L� /�d ���.zcT¿��%�����X��B�O��Z��r��{���Gd���V����{���F)���"�z��N!��H�I�%]�!��JE�RD�R.��)K�#�#*X�,�������р��{���*n5H���L�B��@�и��	��=.�#��	���-7":�� )v��[#�{�L�	|Kݲ�hE:����Ax�N��>;�承A�	�Ӱ�4ơ%]g��'��bM�o"<X�ǅxp'n�:
 X��O��g|wi%�`k�S�r7���jw��`N�[1Wҍ^C`_
)��~�?T�5�þNA��A�����	�\�� �o��a�2���0EקU�iH���-6���1"���rc�8���C����7�4�����Ú������h�Xa�vA�;����4�[��hvg�cx���&�}ŗ0q֯�3��u��"��g�t����-
����o�D�>�d������M�i�W�&�y�=���=�P��7�}8����)��t�F�6A�x���M��Ẑ%R�n�IJ����#ہ�)�mt	�D�G�@y$��620�ZH?vpy��0�N�P���E�%4�`���ͮ�5Y��#���9x^�4'���R��O�"(ԁ�p�z��ѻ��+��x*��*�Η�`ŋ��f��Vj�*&�g5�WM�ȕ�����o	Ҟ��XhoL�O[�����i�}m��J�xyX��h����z���ٔ�v���� o��XӬ�<l� �ϳێ{z�N�|]{w-@�|�b�d����������u,��� �\�@�u+��I��G��#��5�;��Nq?Ě���B2������� �2a]�-wj�kQc��^xx.e�QIq��h���tĎ>а��~V�7ѹtp�%^�U2���g��g2`ϋ���a��>=Wf5���&5F&�S���f�0��b�z�GhM�h0�g��B��S����ow,���ܷQ��(�F��_�BТx;�t�OLƏT�KU"�s�Ad�F
�a�C��ڢL)���,��}����B�!��<Fͫ�dnҝm$��(�6㱭�-N�����sܴ�w7��x�skoX,Z4ѡ����CXy0sX'EA�_P!=ҽO.��K�A?H��K�����?�
�"���EW8�aMM�c�����[�/�����)���� ������64T��d��Xi���0&4��S����f�O�N�~�p��I\�X�ɠKP���|bc�(��P�Eł�����ǊL��߹fh+m+�=��k[i Ʈ�[��@�L:� ���79n-���c�\��k@'��=��S��%qk����	GS>�0���S������]
xyb�6�ܑhԕ�R{�*�#O��/�� Y�RY5[O+�1S�	�l��G��,,�[��V��	pM�����fa���­�"X���aY�]�Bkw���熼?��;�U]q��> �K+8@P�w�E�i	+bF;��J�I�^R#�;K�h��k�$=�WB�n�Uh��r{��*|ڥ�|=n��c�)��9?�?P��a(�M��!<�Q8|�am��ԃ	F�CV�H��Ɯ��p$y�R�v�	��_p�[ 8�Ș?�A'�=/m�SӼf����e0ifC�kUy�}�C���-a��K��{����+FB
H+[{��v�*0r�1�ɘ&����
�fv���^ê����19�b��{�'�ҋ�lm�!��?�;��~N"
0Lͩ�_�:���)h��:��UrcX�5�)�l�w��
#9�6 ������ނ�)㱱h@���+�R^���:̕i
W�OU��2-{���2@@r8��Lp�]D��&IH>V�:�X��U"��d��:)�;�so]���p�s��tjy������_#V"i��;X*T�n�9Ƈ�>�|�e_�a��5��J��F0������&u�k��
���ɡ�(5��,ĩ����wT,
"�L.b�[R�ϼ������u�&��ǽ�a�vSR	���Ⱥ_�N��\q%�5���8�Iu��$�u�;����t|��l�\�]�Ǹ��9�y�S0��rs��pJ9�C���.���5 ��v1�B|$�4��/?4ƽ$�[
L]�b�~Qiw���z�/�fׯu�� �{oKj\b��
hϨ�\X��*J<���M�`��������F�Ĺϖj4�͂5�ˈ��.�[�y^�v�q�/�W��4L~s�	3���P>_�4�_%���zAa�Jj�c-�5�SQ�I�3+��"T��`�גb~��K�|�,�^2�<���]zo(P�c���e��	�Y#��~�f��}�ܪ;�ﳇPʇ�wur�0���.�\ R�n�~=1��Ɏ�ϟ����� L}��/���*���%x�@b)��R��1��Q�9v�񥅻��Z͚o�?ҞZ�f3f̌=�-�]R��S`�5MU�y��]-zhu'H����+�����֭pO��3�����>{�k�M�	��!�m�|�:�C��k7������uU��D���Q��q�,���U����è��<�H�T|��]�ŚCe�<�B��8X�!B��O��fv��g��eZk�R$_���g}���k�.�t;�/�.�sAT.�L�+�R)�ک��%�ό�V`��hE�>Z
5/�h��X��w�����~�x��p𭇯5��|�M���Nxb��ip��#���C�9r�\K^-v�4C�h��ZH:�NX��b�<���d�� )�Z����+h�,��(�����#Z�J�&�I���v��w�ZU`%�CB�[�*�9"(A��s�nI��h*?�`p�hR� ���%�#?n�l�bn���@*�γ~'��y�9ov�5f��1���Y���H!*-�Q�u���"ȇ��F�"�o2�U'���o��*��,�.�� �{����'G��h���F��F�ݷ$W׭�b��Q�cǑ}��<����I ���U(��~�U�T�"5&��GMz��4\}GN�����5��VN����9�!.���3/S��=x�v��n��L]#��s ��F	T���bt�w�r��&+��y���n]�>:+��,X�c�$��wj�̢��~��*"?��E�d�����`���q3j�$�6� {��h�&�N������I�H�z�tN�6�KŬoO��=����A2��:�C�Qx�җT+�@�fwAK��>4�]l�[��V�K+VV�S�g��j��]e��� e�]��5�:P|�V�01�-����-��}`;����5~9}!�� �o9�J؜�Э5���>łoJ��N�����#��S��r^V.��12��Ex{nKU���ڣU��N��aa21�`���o��1o����j���9qP�ܕ%�Fq��[d��[���Ie��X0�t�Z��_���
�.�M�v��Zǣ�c�؉������fF�£�OR�D�]�	M����]��@�f�h����͹:� �k-����	��%*E���`]���Doq�1�#�9�e��=�2"&��؋u�{t�ަ�������j!Jy��M?cd���>+!0��Hٟ&}���b�ƃK�z��i�1פ�]��L+�:�\�3 MίAHo�/�D��\��V�Jv+=�e7����VW����]��7y�n�Ő�&t�L�Y� ۅ@�7P:a;zX�M��8�K�{���t�'`"�w>+�Ń���=�wB����h���3��4�Qt@T���4�5�D��Ar^֚�W>l�6�A�`�O1} �ǻ�+�O
B�w���P�Gؽ\~5�[^`�ݤSs<���x�����fΓ���ӢyE�P���\�ҏ(�GTB�M���zg	���T�3�2�`@�[Y6p�S�����#Ú8�w���=�P�nwsO��?�hC[����qz�^{�̾W���=b;���L\5K>�x��`m#;�G>������\�Ծ&���s�'6c�5!@�k'2�˽��8��pU��_����~d�Y��KW�����K�*��m|�GSI��)	ON�)zZ��γ3
N�KS���V�<z��#r|E`T�l8]�r�6��U �Syx�1*3_iCc�`�w:�܄A��1�r���q����êp��∡'Lt���,|n?��G�kN�ܕbm�0���DU�p�Usn[Ń	���z�7�������aP�i�܏��V�E�s_��Dׯ��\�r\�'cY �,ۧW�O�C���&*���F'�x������)��mƄ��k�I�{�I�p�������Y���@���%�i�ϲ>G�1΍^�6�}���V�S}�[�~��B]8���@?�;�N��~U��0+�PU����^���65��K�;���,� !�ye�k
<�ix�DTO��D�R���wGR��g֘ZǚE�#���9uᢨ�ڠ�ǫ�=��Bk�ǁlP{�A�@}��,�����1F.ji���������<�&r]���}��0�ey���x8���6�9W�{�2�%o�}#R�~Ω��"������b����>&�M��[���*f��b��4�4�1YL��o�i'�Xx�-���� �Tv>����?*�}�ǳ���\v��ç'��Oq0)Yn��Z���
��?]ٗ��!�mspmw�IxX�ܶ%��W7��B��j�*�h@*x�K����W��W}f����a�7E�|QR�ax�6�=i� ��DlLjW���KlM�!x@�!��*�)��"ҽ���d�Z���6<3��,�}tG�6*�f��% ��^���4҇�L*Hl"�|^a���`��Ky@�:[�j��TO*��B��`��^��E�)E�/�f8|Ep �*��d�7v*H,��[������S�\)��hUbT���ѵn�7*͠<����n��A��.�������!�.�F���;l�{��w�+���=<��;�����.���-������O��e��]��EX���YP���8E�P
�0I�Wd��r�4�.�����[�s�GR��l���P9�����S&q
4��ߨ�iz�M,}�L�k46�����8�%a飩`ҏȊ
��$���0�>T��@ ��c�eR��6�$>����ދ_����Z1�T�cu��i�$���ݮ��7x������C�c���R��5VL|�5�g]x�Y]+�&y����.�b����!�~<��ѧ�����@��3yO�!��RD}���Eum1��U��P�=� �8����i�!�9���'s�dY��n`���#����R�c��A�ۅor��U�<�\BHr�_d%���)c 2Ei�8,.Y'ps�c�;�x�W��9��ƃu�<]w���,0Ns�e*�s/]�p�.ޑr�tg�m<jF���л�c(q������N�1Z����� ��2 s�v�4�-��~vqZ��띻߂C��I�P�;<�>@�[��Hgn������z�{����֌
��a��?}���-��L��R�(��$uq��)Z䀌�b���H���C��9t��J�ݣ�Рj������w��z�Ǐ�R�l��n�S)b)�f���7@y�D�ů�����4Iׁ7U2�כ��IuF����N�N�%"�d
�*��9 Y�ТO� $��>g��#<3��5,�O��L�௒^1��7����2�}�}���{_����.=6�-<k/�WDdn׍�+;'�(���wp4�>$�"�r���Fz -z���\�EU�_��34;��?��˦�9JB��5λ��B����|�5w-@�I�$F!�S{��(��]h���h�#H��F֙��t'{�n�����i��.�Mq��_��JK�#w�]�tjέ�(u�-��3�;j��������W��N��a޼�����\�&�#��f�$%s�}�bF�. Pޗ�OWe���u���q�g>5�tQ�`���]���{��%1��M�r.T2_Rt!��x'��xOAd���]h�<^��ͽ���q1}��W��"�K�fT��kl�-���b$�X���UNT낌Z#�1�Ҝ�ؿ�MFiY��4�&y�_g�GɌ_���PQ1�=W��F��N����MX�A�=>������:	���ǵ��_~y�l��iP���^��t�x�#�5����ysP �<F����B�����r��t0Um���@�5����8��CЁ��~�͑����|_9t��X����P�G�b"��v~��[�p3�u�݁�a�%O^�pr`�,Y2�����V��SF�I���=�D"���gs��	��v@���\�,�jx�s�%��n�5���p+�g�r�)�Z����n��M�I]�Չ��-�̩(��3��i��}�β1ey�P�� �]րm4E*���<���D�~ U	@��_(*�+1�Sn]Jw�@�q���)s��|I5�|8p��J�JGA����ډ,	]>��H�����(�TЩՏ9�I.e+A��M�ע�0���C�ī���ǜ�T�����C8r�_�����fN�9Y�O��֜Y�E�!댸L}q��\�(Q@Q&�p���Cl�	�R�s�g��#Z�l�S��������-;&�b!�����7"r5)�>���� �>-\yn��Q)׏�,g~����/��(��+^XP�c�HZo��9m{J��]*,���?U}Ų�����Kl�:�m��#��L�֊��Bv����7Q���l��Z!�A�τ�Ex�~�y�`�Y��:���,{2JA~�}��q2��ۜsѷ�5W
���Z'�D��2Qt{'�,�SQ	�f���C6g!9�ɖҔVWP?�:���l�3���"���a�-5���t�:f��D>N�Yd(��}>�J]c����&w�=�Y�%��n�E'B���|-a����<���K<�K?�t���Bj]��i$��_G]9��h�g|�yI�^�z�|Xcy:=b��MaE6q��_�����z��Z��˰^��kǸiXp�1�!UBYT�^�[S|�z��]	usk��&y���,�t����Z�n��vʦ�4BC�j���C&N�D�,�ßiK= ����/�	N�"k	�uh4��W�],��Ճ��i�~�8��X<�|6��(�PW��J�m(=�j�O��<��%��Ƿ�M~h�X[�P�׵���%��F���/�Z�.����́`Cx:�(�sR�� ��_�FS��:�"���#��p�n7�lx��6��F�m&���Iu&��i��ݘ&�s���K�T���qx�	�՟�7w�|yk�C?j�'��i/]�MG%��v����c\?��	�=8��4��[6L: �n��Ɯgue�[�6���wzT"�B��瓥P�QE�)����I���Q�����9zWt��V�t��?=�q�� G��:��m&��$
;�	,��%���B�%�*�� �`�Uw�z���'c(z���G�!�J���`D-��ψqi7K	rR�7�)M�%t�(C�u���5���q�aк8���n�")�*y����qC�r:4x_�q�?����I.Z��LV�E�6BJ����"���[�c��q��ޠ���u��n�$����餕p�2}.�;�Wս�**��xoĆ��+�1
�,A)��! L_H��9���RqD�X�\}_���,veO� ��P�����#��\�^����;����y"���u=�(ʃ�8������J�3��O���2�^4>���Y�"��l}������;�O��h�#k��x�Dbb&S��rg5Ku�<��
B���"�İ�����q/�����Ɠ���+?�E���m�������T��|�~�F��� l!$�c��0P���� ?|�2țB��3R {���gd�]�Z	tg�Vn.�r���Nk
�֬�wB�]ʯ�k->�m��r�R��L�}��ݱa����QZ��wWA5`����7l�i�7���゙�<�&@�JJ*c�(��FX�ީ|���Ϯ�*����	~moͳ����ꎱ��3�z��ĳM^����3?�?�(�Y�A�F����:t��X��.F!���� ��F�I�昧o�IBj-��UK�t�~��I '[�W/�ѣR���ͻ���>��b��=lMЬ|�����g�w�k�D��5���.�����F"�̓�#�k�{Mϖ��ES�k���4\�O�u�`�2�`�#���;W\�s���x�c��cU�#+e��O�Y�G����8 U��s^�+�/$.�)�zM�2�u)6Y%FP�]�A �,l/\K�*�DQ&���ti~M�?5�Cx���ˌ�����+���6ݩ�
2�!u 5�mh�X��(tY(e^���_��1���F���ב�B�ӻ6$s��'{6��G!����0�oK�Py���S+[W|Iwc
ۘ�qtu
�����P��'v�>2�h�����sHk��_�y��|�ֈ����]�K� R��6�n"6b��X����t���4�H~Bs����A��Y��Z�S����im�&m�1X��-�c���	!,������	G?'�e�{����LK��/�v���8C��$ƣ}ɶ�(H�H/lKe"�1"I1�Һ�P���Ѥ��;���t2=�����+��"ސ�O�H/u��U���s���%�D��L���s×����ډ&��s��Hp��|2���v�Ҝ�@2��tUO})\[�5�KY>���f�P�U$��V;3UtF��yB�}=[��A�#�)048Ϯ�-�V�Xo[�l .0=�\�Q������H���R".�0^�a{k`�x�gQx�t�?��B�
@p��w{�.�ET&�^ю���N��� �q$\덺��&�9@��B���.=���(�D�C��YЛr�V=�7�ȧv/Ue,&�=�h�$_:U츒YЯP���2j,V�a�VsZ`�q�@Co+��s9~��@��u���8>%T��n�8��a*��֧|0�GJ3����j:�KW�2�]]6iH=�C�|$�����k���՗RńP��L�A�´���)]�
�7Ҧ�{Ƴ�.���^A�Dv��_^V|�#j����s��S R��3�	MV�6�/\��]�)/�u^���T��~"y�R��p�I�>�s�5
*�\�
� &S
�X�%�ᮬ���͓��f�a��X��+����P$�9Ӣ*��׊��ҙp��x m��8��1�;Q��r�(�Nw��؉��4�Iv��hl�_#�G��p�-���[6�sUJ���A�"��£�N^�,��Ա߾8%��0�;��P�\Hgx8h�[Ns���a+aӏL�]Q��f���5�i�e10��8�M�^��=���\��pm�'�A�����|��e�e��1��HTx�hkN����/6��-�n������җ��Ln�o'��@%��4���є��t k��39©�b�؏��˘�"�b�Pu
Ũ�~����T�p�/B������&�!��}:ί�+eO�	�r�hI��g���l��
~��l\��Z��F�~s10K�>?�άO˙�G�ٿs�z_�6� "C��+��Wq?Jrc�b��aHɤ��:�ai�YW/%<�on��(�B��gU�P��^�� ,%7��0O��ĳu<{EbvG`
�����,�5��]��	��� e�)X���;��!`MN(������_$�� �����w�)1���D�z��W�"����K롨�Sþ3ݡhz����� ��e)�_��S�S/��2Yv���lq��_R��v��<�ۯ����e�5��(�f^.��"�y��Cfت�M%�(Ԗ�5ҹ��cP��9���h �.݊� �@d<��,���	��I�E��Nn�w'W��*:�{�]d�(	�Eiwd�m���ES�|*t��F��q(>t�y�SG�ArRaq�[�g��D�K*~��a�� ��:��(��mFv�һ+��s�TІ�j��B��[�Y���I���p�J���A��sBs��Uۙ%���!OHQ�z���J��#x}o7���ɾJ�Ԫ5Y@4R7��V���x��aRX����HTU�ѭ�l´�o���9~(��EB�.Q�0�<���pm5(��g�E�:Y��H���w^����Ս�^�;�4߁"����̱ix���?���%_k�H0b��}�B]�f�0��ʙ'��l��)r�l���{�l�(�pw��>}�2S
���)�Ae[J�&�����zn9����Rj.�6t�K{u��	j�y:�Ҭ�js�M��\L=!��$�����"ʽ�sv$��C�$N䱡hy߫����o���E�����I�]Z+q�r3��LK_@�aU�jq\�xZSyi�٠��H����3�z�lZ֠�:g�k�nA-�����O�Ͼǚy�<aR�oC��A��@��ڼ��\ƔK=��Fo��iY��ze�� ^z�A��+c�l�%M�$��Gr�SyNc4nN�o(�┘[�����YO�R-jkɎ8������yG�;g��%��tsw� )Dɞ&�T��h"�ݠs�qC� M�M��A����!���X���`�*zC�c��'���̹��S	��,^��!�q���{EԱ�l3�E�!J����t��_	�����?�
�f>��A�ԉ�U8�������\%�[v�����;ݍ%��\�1|�f|������`>�2��'���|nȀ��+�eԉ����f���ah�_R}������μO�e���Yi����rQN�����7SN�">���@.�h����+(�n�RW���\+����;�1���O���Gx4��:��F$��N���KׂN�P�Z��-g�_e��=0����*AQ�c�����m�6D��"k�M�@�%�d�8g>(a���[�A��MX����W'��b����<uE�R�4�>yq~Θ�Ԥ�J��˂�7Ĕ ���fԔt����]������[�����õ���M
hu� )�Fw'���@�U qX ���*Rp�A�_��e2r̢8ZS���
�9�����*��M;�{��Bb�豞)&�ڞ@�D/z^���
R/I&�֜8ib_�=_�3.J��ɶ"�u�<{��!N�q��~ -�Sf����/�=��y�SE�6�n��$H���S�}tH�O��!?�'���ݿS��`�6�F�A�L<|/�5�?����9��է�+�S��(��D�З�0��c�0@�;
�U�p�5���H�W�j����%�4��⬁�4c��5j�
y�䷀��+מ/v�����; LE��4��ԯ��BL�����H_Ⱦ��]ϳ��`�-�A4�~�/�Y�]R��:k~�sS��ѝǑؔ12�5�Ɵ�=� �İ��a� U�Ū{��$D��'2��M4�h���Uyo�J�t�0	���o�l!�����;�;��*;��X��U�9�[啖��ߪ����;`��E����2���;�' -,���~�}F�$��[�����r�Ӭ�-��_�ћ��Y;5j�x"��s�s�D�z�^Oz5��	���ٛp1ť+fz6���QK���i�:�G�$Ql̒�ÿ��9�4\���x�V�)�m�mHȬC�~\6<�p�l�Ez=�9�_ё7���6�"�$�Rt!���/D\+���7������Y+{Oe��&��������3��(��~�&=U_lj[G!I=����3���w�SMв7�UJǰ��d.#���������E�$�d���F����5ǐ��Hn�%�/%O�ء���6|n]��	�j�1���zܕL��I\'����z����y�jߏO��DF�k���`��(���f��b�݊�"2��0Z��#����e��4�KOdJ#T��@��t�QM�n��ԭ���������1�*ex��8��w�Ӄ1S¥܏���n�B��e����D�U���k�(kp�R����Z�/��u�6�z"k��q?�"?̭D�pC��f�=&�ȱ{?ϻ�e[]��� =�W׆���3�q�~�ޫ��&�(;��&}��o����Iy$Fp��^d�x[|�jQ9��dO��È��-��eͽ�Cv�!��=�88�v�nl�¯�h�[x)��a�y��w3+�5�������W�u���3R��Ϧ`�A( ��Җ���2|�$��Xļ'd�勒��㴋R$�E�l���8���F
ڝeHN4M
e4Y-�~�
C�>ͬ<tvٺE�C�7�u���ںrk�?��	P}&�Y�+K�W�s$�<� U��������J����e�p���)�Ὀ�v��"U^��ٝ��8i5�o��a�5��9�ԉw�^��;0Yq�y���}����ߵO �ڬe�Pȿ�zѢ`�ۓ[b���R��{� �����5O�'W�^�.�> ϯb|���d;i��Lt�Iq�ѠM�w
���@�p�i���l�����Hd�. <B��,��z��`Ä��=���u�N"�#a������Zg/�&>H�Y)�����r[��T@���!�&t��P�aeWtpM�NNb��CBmSuq��Z���K`�f�Ϙ�n�����OP�S��e�`?X���|X��g=-��N&y�bsZi���2��1�!)�3�]����M�#��K�s��u'	Ij�#{�ފt��K�mOi!�Dyxd�L��d�VH,���X�`j⡓?���;�>H6�����-�����EX���e������c�heT��$'c�RLR�P-"�Z�ǂgz�܃}e��E��T�����6{�rΖ������w�K�xE����hD1�P��
`�p5�.9��qcײ�K.�q�i��r�ǉ����:�] �"Ǵ��R=�ٲ`��Qqř�r�S�	g��^ipT�s�ru_��Ab����.=���g������*5|W�%�KK]vCM3��/V�Z!|tz��f�-Q3�$(���$:�P��Jy>T݋M�"-���]��v�"��Σ+i�+	���Roa^Q԰�ʂ\��ٿM�����(0��r��̋��'c	I�/kfBQ�]�;�BE �[)A��X[�6&�MʾB�0 �R�̔��\������/�kl"�`[�}�t���-6�G�$���EdEm<.i�W����U��.P`��ai�R��$3����V��{|��GaHRY��)�2�ǽ�9�K�2w��ɻJqۖ�R�uC�dt_�e��Q�0�Y��M�7�u�d5G�~,��6˹T���w�X6�DLU�7F�!'�������n[�"z��ڏ�'�[4�ض�+��w��8���g��������dۅQ��!����pa��" " \�}�a���`·��1KY~GM�|ҭ����i��wc@�֩2���~�ܡ���5���=���5��"�xlN���;��܀c�P�,+�ɸ
�8�U�N~�����?mٝ�ם��քWF��-����!��Q�'�:Ky�0�l�tTmV\H2V��MJ�C���f�c z�u����A*�����	�����W��l�ާP��a�K.|�[� V>4���A��̑��|���mEErT`���f�~^�+�m�w)�z�|�c���}/&	(��<�� �w@�ԉy(W�si��5��0Q�Br�O���j����7�,�a�O�%Ԣ��a9��++O��c�H�S��u<`��as韑| �=�}\m�l���!JX�2>g����,�E��iC��jS��o� &;. �Y�{P�[ym�@�Q���ZC���g�5Sі���u"��=���h���R~��6�އM��Ne�+�)��Ö{��f��y0����>��e�]CWqFV"��n"O82�m�G#QzSS��~xmm{�zZ7���6(�e�Y�A�?��Z���^�\@#(�وo;#����ݦt�l�d��xA���� ��7��
�;�g"8&�y�g$�[�Yjj�	�䒊쀺��h��8�s=2��
�Ӽ�9��,6��V现[��4,�8�ׄ;�����2`��ᣪlYS�ʱ�bz���%-+���n��B'�p_jy��5�_�x�jg��i��:����`x�r	�{*F�C��UU�[����E�V��n��Fgj4%�A)������{q��{�<���w�>�7�}�	��D�4\:�Mwd!P�K��a��S���c�T�0�H�|��rM
s'�2���_�~�9�!c��Ȼ�p3�r�̙����Ԭ����2�}<�AN��Z�3΅�u�w_(�h�U�nr.x�BϪ�G���3!�~�a��(G�&⟉�{f�z�<]/2n_���e�35l��ma(��g��Q�� �s�#If6�Uk_��XR�J�ͪ�M��ߟ><�1M���pz��aו��>��p%�'[��C딣�A����͞R�|�E�!�W�h'�����W[�|ν�_�IL��Aͭ���E����&�N֕�kDk'�KJb]�����2pxt:t"S�(`���b�χ2���F�`��
�5��.%��&���E��6f�ɋ�M�{ҵq�7�N1���ZXjp 5.�2�&0�21x��|%�� 샣�9~P�Ϊ���w;l'1E�a��whw���s���Me���#�:m[p���Ĝ�dX��1��i�x�9#4[��%�$�����,�綴!�_�1�U�\%}�g��X�p��'�o�Vl���.zm��6VՇ��y�O����8D"[����W����A�%��O�$%v��>X��[�@�-T��C�%��dC+�U��/����p7��fuq}}7��]�ړ���7&�G�J�Sz{)�:7���2p�%G;���["bzr��l��^�̘���Ņ#1��n��
 ���w�=����.�:B��d�G�t{*�n�PL�N� ��W+d��/��M����x�zւ��G�eP�#s?�4
��/�������c�]!(�-�fe�3�.2�	��+�/�O����򇉎�t��*C@@��ʛqWX��x}���z�k�{�Z%%{{��Y3.�}��X�ίC�����]�
K�Sߦ�ٯ�E�ʤ !0��,�>N�����2��h+��}��CCQ�ǂaC��^�����*��	$
���S��t��aCS&O1]�݌��7�[�?��hRF��A�8���b������۲�a�1kC�c^�X��<��go*`v�R�ݬ�M��=:Q��A�����Fޮæjgm�����Zˉ�@������?��>T�1x|)̒OƸs�.�05;��9ӊO͠��
���~�S��Ҋ߽���:S
t��<-���N61"�ks�G����d.�R|�;�����9� �l��>���9B��*2lmR�Ew���6�T&^�p��'w���'�Lv֦�!�����t=K\=cx����G�U���w	�p����&F��*�!��_U2)���b� �c�ǅ]�C�;ݴk٢�9#�P�x/3!4SO�y(��2�Ͼ�PAcv?\�f��3Cj���D[S^����J |=3�i���/��2,�luD9'����B-Ɩ�F<�ֿ>c��Nh�����$�3t;̄�7��9f�	���t�A��������"3�o�HГ�롸š�x�aCjn��Gv>k�Pp�y���BU�L8F2����ڵF4��o���rs8{��&�N�L��WPR�{M	kzr�<̌��U=���(/��4UN#By�%_]�'Шwh� ��Az��Pʟ���Z��I�4^�|�Tz�����[����{a��lC��j�	9o&�GT7�)�� h����N���&2h�m����_cL�zG^�#�mP@�l �����}�ӭy�T�'$wĕ�T:%�	5���p�d���V�ڠ�Ld'Zu'd�v�t��v���\��k*{^�����ۮ�m]a  ��3l����⇸fcr���<���tQZ�}�As�����1Q�@A{�����N~����B`�۩l�Na���y藥5p�t�=�,ŝ��b8��v���g�1�t�q�e���(H��엤����3�˱/�KA���c���8��o��VH�Ab�۲� I���o��5Z^�8Y��YI�M�?�R�����	B����I�b8M���>q�i��K��݆軦��b5��t���&��߈�M�� SJDS^���� ���t���&����X���Mƕ\q���nS�!~��Zg����&�,�ԣ���*�>��nFq�I�h�S�<oAL�D>(m�����߽�>Γ��"j�$�ox���#:z��
eA�fC�U���RaP �//~�d��[��ba�K�AR���(�x����~J_���rUuR��E��v�r�*����kq掭���i�aH��l�Q��..(^���P�Hy�ٱ��EwK�Xa�Z|Չ=�*�k) ���%r��&]��"*Y����.vG���}E$X��:	zr��zbl>ɟ��yz�9� ��W�8��r���Ye|k	q����Q�LEPg��af�v0��q:~:��:��/�%���L�v��b���S
��{t	��Y2��DU�!�:\o�A4A�h��5*����Jչ�VP'L�L�C#6���#�^B�X{�����cg��fJ���٪�c�h
�>�̲*#2�ዮ����uxV]�$�R���#�����eRY���E� 8W��R��w(H���i�%�ո�,{lX�w��������E��C�3��;ޥ���R��]<��c���N�2�PFfs���[q叛ۈU���?2�M�b=R�VPҎ�7$J���f�V�qoy]��1n���1T57mc�t�s������,ԥ�f^�\T�¸�b��F��� ���4GK#����4sK&I���;B+��;*k�7�޴х��;���'�0�@EO����\�O�
�C�������Q�K ��l���#�^����O\<Y���Xqp�֣-���z��,^�V'��*[����=o�v��0I�F�bq�(��P�[���X���:A��� �v~_:LV�X������4'k��$��o��Y�*G�jA��K���X�G��iz��&��/``�?v~���%#�P~�tm��*�E�N~�Z��Ka���k0!`�:J�7�	��T{ă5��,�������<?_9.3�̴kݖ���Ђ[a��t��D�t% �H������[�9�� �B�pr\	��Z,2�R[��.zS&mc",��x�a�S��i?䨓���Pkʊ�����[I^F1^0�y�a�.�&'s���F�ј������qU./����H�@�o���f����hI��p;ucrq����S�S?b�����5�{��I�闊U�N��Qn2��s
�ɡ��!T���g5d�#�<Ç�K�
{-S���6,X?���j	@���d��1]79�v�U5(��l[������;��P�ynZ�I��);]�ߕxoz��Zq
�J�Y.MM�\O�ou��
`�A�
�jn��[�z��i�����GR�4h�ȬH��sVm8�˿�
C�G`�L�;"Ei�A�)��ގ����^M2�F��tI2�[�c���-��ּ�h��=����+,M��8-ҊɱO�lw[���-��$�M�������h�U��.X�y~]}��Ԓ�Ca���pV��O����
`7J���~�R#b��l���vn)Q���)pG�e�8la)]�O �x����P�wO�����$w�g�!��?��k�i���.8e$?ZX�����1Mq�F�� ����a	�)����_p�P�A�"F;�
$�:�7�ĵ|::�K�t>�z��30���R9�,MH�Zl<q��	J`�0f�>��Pe�=To�2���X����9A�-{ZFZ�
�_8�&�7Q��~��ӑ�j����g-������t�n�<�\��2���;ʆg�KdsF�-�.��܁A�g�ʛ����������8V2�nFF<���g���V���oɫ�h};�0�уf΋�k��fY�C2;��BD��b� �dJ�	|��kC�2?��t�.�ʿY�1�N��;Ts}�n�fg�(�YG����ö�־�&��۫C��49qV5��P��HȂ�����O���؞Y�n4im4dOHD�&��������M�n��s��^Ԃ�%qO�'�6ԭ
�ᯧ��iO�za����U�}����?��p���(��
��̣k���i=}hdvY�I�E�<ܠ�e֯^+�K�p���8c�R�b�h�OQE_paV��Z�޿�W��3ūx{�\Z�~�N���gR�9�������D���e�����d�^�Y���"��N��teBN�QQ:*���|�:;��l��XJ����~��d�p��R3�Z����ݏy{D�|��&���`��2�G��Th��$�����	�;���˒4��&�}I\j6�z����{..��6��N �˥�_�,ȟȘI1���&]��	���XNX�8P���{0 ���^0��0^��Y�%va�\ٺ��.�L��>�5��?�+ƭ�+���jg0�����"7qۜ$�u��%n	�ϯ�N��%�n��r��+`Q�]����;)�6z���'�8�cr ��ʰy��ޜ���@��%˪�hM���AY������.�Oݧ��R�)Fg4MY�̛2U>G-�Sz��m�~�����1�CB�N>W����ю|Yc3�:��*�R�H��[��_�6���&q���7���0�:���X����1�ב��CT���z�ӴI����/-��Q��!VO�p�u�Bt{�J�1�ˋ�"ܦ��bsb�coq>�8ӎ*`
3i���\H��F�9e�� A�m�E=���\�J�&�Ah�X?�u�%�1��X lf."��;G�ef��\P(��q�1�98QQN�m��&*�z�4b��=�f��XWB7�k)ɯF��j����r�\��� ����T�߽�n�;�F寉H�¥� �bS����(�'o���LO�=M� f+����,?g���+8]��ܓ�~�=[H9���E��ϭ��pu�:_�>�"ၼ%�-&��F��fs�e 6J]SnQ��b��9��Z�F�P;؜��z�� \BA�A(�i��
�I0�	l�;!յ$�Ӈ��ȅ�qL�e�Q.�+f��
�����$�z�Q��.�*��Q'C"fX�� #�3���BӢN�J��#�B��*���6j�1�耒뱐躄���{sC��8�́j匊D"�ٽ;-�Ӱ}�ܜ�L߮e��ia�*=�3��,����e�">��;�Xr��@5me�w�4H瘰3�T�#ߑKΣ` C��Y�}�5U,�<�
���ŶC�-�H�@��.���9�!�
�������i�mX"!f�c���ݽ}�#\�&c���d�;]lp��:$��]�p�v�n�kq5�����͐��]��5N���b����` ��O��i�P��X�V��ā%v9%&M�V��JKo�yɏ~�H�/��4�[�v�[��[w���n�nZ7u97#1�!YMRY<��"B"�4U�����Ί�#�A�ާ�H�7KY�ҧԙZg��9�����޴��[��c?�%�*f�r�۴������+i|U���]�����E{��b��.��'L���Yp�{p�w�B�Mo ���aE��8�z� �v�oKn-���S�X%�vh�vq3�Y�,�����i|g/j�FtYT�ԉ���U� 1��MLj�h|���$�H��\�(�I0�$��B�;�����H�5�y�H��d��B��/Em5#�.�6��NW�fD���F[��<��C&D�A�q5vN��E�\�|(��)��S����)�鴃?i�MXӀ1(2�ٿ�=��؇P�lc�8ь��FNdčv�a�2�xјoŤ־�BP��/�0�{��EҜO��Q26{}�#� ���
_�",�PY�D������Nv#�p�Ơ�B�����_���ǣ�U$$V�*_Z���Ķ���8���h���CWg��BV��J0 n��f;W� q��Qi�5M��[�3����.�4�<:>�V��:W�`��'D���Y�1ʋ+�r=��z��NV���q�C��	�9]֭_U�g�l%c�XAq���LވHk_��Me4r��r��yk���?����i��꣝�'�0k�X��g[��$��
�Rsw~����IY�ie�T��}Q�W5� �)!٩���́m�wZ���CN}%s��<ߧ6F��'��́����ܻh�g�~�V�⌫X~~l Ύ5���v��h���f��U�tR�,��Ɇ8؜�/g5���g���AJ[ûj�"\J?9�l��Z�`�
��y�(�6Im>�L��s�U:m�}�v�+� j3�����,XS&O��ZB�)i��1~��Lu��p֏��m'�a��h�_
v��@��촣��6F�Ame�`ܢr�J�vً��f��;W�_d(�,$R�)���A�X9�]���HOa���$��A��R)���(ڳX���T�T�E��֖�:����l��Lu�/�	�������*njP�K��i����i��o	��k炃�L��-2ܰh~с���w�g JR���v-:�K���xh$�d-���Pч�~��Wj'�,-K�x=�P��U����h���Ki" Οj�	uxĜv�Z��<��Ŏ��H��bJ'�q�x�U'S?�L� SR���ÆŖ��n�hX�N�s��Y�M�Gq.z�T����4�`=%�����S�2�X�̔��v� Cd���"�ߞ4�@�����kW]!�h�I7�"r���G��+��S��,��Q귿p��/��|[��״��|s��vnJ,�I���_PuL�.�\F���Ҏ�>Du��S�Ǯ��= @>qŰ�}^�lM R�rg�q#�r����9̒��dWR��X�;�U`��P�r�Y�Bp�`0�D��Ү�7�@q���Ծ�7J���lœ��b]���*�ҡGU:���l7{��m]A�o�� ��9)��%2ɬf����Y6��in�bu8������p[<V[	��� ��tظL�]�È�ae�M��d��V�����}�!	X��AF=�MN�+$�כQ�Fڕ�sH��Uh�tD#��#:�z�e�6Q����4_0�qWru���vn�Egg�����i����l{O4:j�Uo��i�MΔ3�-W.Yi]"��1�;��uI�ih]��c����8ݦ�$[$�� i�ZQ��Wl��(�}s�س�T�3>.���h�1����"�_���Ri�gԪ�ȍ��� }_��,GsS*�����(�C�����]��|����A��C�����������b��U{М*�_H$��t�o��t���,LA�s]�AO˭xݮ�~���X�b_�g$'p��*�*ϠO�yo�-j�Q��^��11dT�1n��G�c`�l}F�����9�=����2������&_����xL���6�$j�se����+�si*���:vv5Ǌ��o/x�XȭY�g����1��Y��¶
�`�91)J�4R:�w� f��5�'� R���>�ؠ�g�k2�ɟ-��1����nb����2J^�%�)%�� �G�얉�#�=���L�)�>x��:Z�,f�� 5b�GMLS4`��,�hw��q �J-�1�5��L���i�wp����i��.GTT`x3b���3�p��(�N�P_�Ul�kt
׉R�boA�_�G۝B���
����$�s��rؖ�:���pp�G�il\ ��AS:�C���nD7ݥ*Q.vX�1�ͺ�a�I)	�	�v�7銈��=�r$�R�/ҁ��R�f�"!Ӛ��/Ɇ��R6�>�6&�A`���0�s4���7B65�O ��Wf:���'m��e��� �X��̏#'��]�!�;Ţ�oG'� ���ֿ<k�Y<�ߙ_���}t�����TLN�ʝwbZ�a�϶�6�7~F�G�&�!�E��O�z�#�Z��T�=+]�K���8����#"�+�Qf<�H�Of�+@���Du��A�=�ٺ����0�f3� d��Gu�A]k)xdy��l��g
��L=� �lO���r*��X��,ӓ���<�}2��g�^N�Q��ʴ&fti9���N�,���b�5�\�M��K���J!�;�l7���ͫ��`��@�K2��p�RЭ+sB���v	 ��w0���8��aey��~i`��H�_I �)�H�x���|���M�zU�wl��X�[��9(g$�Ͽ[h#+�5� �P�[�'�cًl�N$��d�/o��+c�����noX��~+�	&ڝ�sKV��@�.�*�%���U^��B2s��o�����̲� _��`�
*Gxp�~�u�OҏC���w�u�+��G��~Ve��[�$=�`�W��(��)hj�mD�(?xr��9�Oq8�4"i�c(+s:ۤi��a�ʕ��^o[6%��Ed0k;˞Y"����߃���z��tx�]qH�*@�����o�G	�w��Ӑ4l��*�A�\�<�39g_2U�W}���R�\���:ns!Fx	�K��X��E��3��U�-�-��@���'�z��`b�J���i���{
2�:��]2��NI���P�W�'���wi�����	*o?6��7P��Rʉ���h=��y���y�A�S��8��%�C�����A}w��6��]�#��Ě-w���=h�ǁ�\ߑe�+����kҵ��@�W�`g"7�| 5�27��|�3q�`��4T���,R+�u��C��Z3o�'�g����~;Q�S�$Jc-�ɠ�,s�)��|�t<�,�~���>��J}�5�2.8B�[�/�,"� ^�ѫ+A
q7lH�B���o�g�VM�t��Zv��ŵWU,��;���5��m�b���c��9���W�q � uoap��ДR; ��Q�u��:��hO��T��ᢐ-�{m����I<ǅm�FR��+�����%�4��2v���֌�WĘ0�R���)��Ҝ��%Jq����g��J�r*G���jr��Cb��ʡ�_Ү�ٓypGr�1��6��SiXv4�)R
�a����ȸ�k�O~��1��lr�]�2��Y[B��Z�-\y�G�l��@cD#GA�(�4�x�8mJK\f5��C�c���)%����SA��`���u&�l�'��T�.6�̽�~���Y�d%�?���]��iaz�-�cc�܍��c-�T�igg����\Q�*�]8�?!GP*� ��@��*���|H��T�n� ��k�ا���ͯ��Y/ðD�����S`�̸>yG3zg��jR$����`X�w��k�K��/�W��0�S�����F��n���Y�R]��+!n��,{�(�c3L�pE
:,>6��܂���d�F��pc�dT�	���AQ��XM��TO���͛H����?+>h�H��K3:Iq
읹��['�,�^P���]#�2�����1Pl�6:��YZQ�� q%$�x�h5�p�8���p��A�0��^9_�ͻW§G��kKȠ�(Ö����/C6�~��d���Y���5�dE.��5:��u�Wϐ{�k��6|�_2t��"K|��su�q<�(Q�av#D�Zx�����uV�sz��hk��6^�
B��#UY�fؼ+z�H��9����0$*�=]�}��
��~.���m�=�<H� �F���v�1,�E�軷
�9����&��C��F?L/n.�
�d�pA�G���ڭӐ�J�O<w.��2��E�{^HV���d���IƙŎ7r|���oO �>K� ��y�хa0s)`H��k�q���О*Er�Z�qv��#	/���~'A�@�6�����C��'{Lu"@mD�]2Px�m�a�X��&c�5���@�Z�)t�%�7wF
���/��k�1v	��Z8}���?+��mM�У�^hP<eX�|g3݆ܲ1�bk�z��2�k��ʛ$���5I�V�:L:�0�8��]��$�4ߠ|Z*�k	�\��V�;����<��H��z^g�:��8NH0U-8P���l�R�'ͮ4�����y=��<,�������$��	�ո�p�吁H� ��q\���/��i�x�~��%f�⠅��x#Ǚ,]��.�d�x�:�L���c�m}�t��*�P)�� >R���֨&�j�ōB|�I\,7b�RY��<�����ű"v���F��2]���?�r�Ι{�iatk��	8Z ���T���r˺^0�fW�!��3܌�cT��3�}�Y.����lT,clJ{ZF�g�F���xP��6?��L(��~�����"�l����c<�$�bA%{��*j�Q
t��� ��Ŵ50��([R���O�d����Qx�V:���`�%������)/1e�k��uF���-į.O7bQ��1���5�V�{��GS.Rl�}��x�i�mO��P���_�#,U��+�H��I�&pL�5�u��
Z��p�g�FIc��Ǽ&�FqWV^_ֱ���"y���i�8	<�����7�b ���ͦ�MrwC ��~"f�������ItT�H[�jӟ��؁(ND?)���d���ۣI�.>��&]n&������a�M돎	��n�X�r�N���).�B��957�	���7��"���1{&�ۘ
����*�
�)��Hc,������k��t ���섷ҳ������9�J�7���
}�Z����y͛����.[F�F�7�/g}��o[�O/���!�,���i8r�"�������+.�Y��q<�_�6���O4�C�}TTV;ӐJ�F��3d�0��%���O�CM��B�W��^��l�m�c���w�9�w��EU��.l�6�������oQ_���w��ݩo���$'����M���q :�IZ�L�d�|��dI5���mr��h&�Ys��)_���Χ��V����I���ZG�O�П/�c�lQO`��I�K��#�R�{�VV�''���6���e�s_�p��Y��8�p����~���ZS�$0X��4�+�rN r��b�J�A�	��H��7�Y$�|d����s�锓�:O�Ǝp�P֪!ZP�.�q��
�l�b�]�w7`SWxY�78t6�X�XaÁ�+��XMF&y�)�>�f\U
5lV'Ȭ��=yS��ӷo᧨�㨋+�V��_�{��=�JE���e�J�P�,���M&��!�HCiP��ɟ�5%�bM�+�ɪ��us�uI@O��_x,��v�G�,��'d+Dj=<Wn�~�-���_g$��W/$���9�w�@��v�+��*̋���yT�+�.ӛ��X!#��2)&����]��}3�<y߸����Ǚ��]����m)C]+���]5dK��ڣ��:-R!q��;��}��*2,�]�x�s(�����R��w���| W����[�n�8�<�7Y;bW��<  ���[aI�/��}�SY-e��oNNe���c�Tb�9��?�+b.��nqP�'��~���8x�Ʋ!�q	,`�i�>��5Uu�u�QZG�/�XVeN�5��s1�ې������zQt����P�̤���E����p�[V��.I����r���Q�;:O��wXEv�ozan��x�8e_@E����o���{�%9�?���v�Yv�
4Y(�\�۠�.U[;R:j�}�V���<�7-&�U1~
�2��𻍎�1�4YR�r�Nš�v'�t�.�\����y�Y�$��7��~���/{�4D<.�H��(GQǾY�Y�ꮛE�lV�A��K����@RY��溬�ْ*�e{IDܵ�d\�`	��q�^��>�i��@;�${k�F%�Q 5���uq�h�9�0�?���O_�+%K��gc�g)��Ҷ�X�l�Bfy��{iS�m;�G[H�_�.M��^<8�ʍ�>X���GZ�8wc���1��������9�M�j`>�@�߅Q<�����gv�)��c�C��Mڱd�H
�.�D�����p�s���jFG�́z\�����֥ i"��f��T�9��C��V$�hd�8M�ǖ�M`�#�<�2b,QI�\[���` �?f�L<���lZ-����>�(Ȅu-�Ơ��A�bN�ܶ��$���%c&HJ=߽.4�J}�$�o�8��g���m���Rܭ��f�̹�S�N�*ZV��
~.�p���w�[vR���@3���(��sz��bk���X�ahtF3�Ђ��䖲ua��k���X!�I"��6��D�o~��s:��g.?���	Ėm��5��?s����(��L����GG��z�~E�D<��~����	<0�!�v|J��I���wX�ϷB�a{ɨ�M��Cx�.I���?��������D����=���"N������ &=����#�B�N�1��~K����u�-��i���s�< v�:����ylC��Ax�h0��?=�؛eX���2�gzY8<���u&o��ǲP��'��ے�r%�<W�x3�!���w��._X��?��#Q�ߟSg���jj�$�����ϻ�nC)1���A'�کVη�t�)�9(ui|	��n9�!{��+~evJ��W��Y!V�����X�h[m*|�i���Y&�.
�B���5YB�Y�aq
�\�3�.�B4�(7�|8ๅ�c��;��<�-q��a��(��\�8~�y[�?�~�4�.(G6�1�D��ѓ�{T* �xq���5�>���LC:|��O��~1G�q�?������>����5��d��NI��f���K8����}'#d��@<c��^�Fj��T�G�_&a����IC���C�3�R���eZ��)���a� ��|�K���{��J]mr�Z�x��>"Ϳ��!A�{�|�H���9�}#K�|]_aZ��
�q=�.",d��?�*fۅ �2�n�	�<�h��q	�b�ťD�dZ�T��F��<kB,��p�-��hY=�k.�u�y^��	�~By����e�gH�0��w�֕t:&]�Q㭻?��7SP�8��^nz�X��,�)��F�gi�^s^�?�T�=*�w����ǿ��>,�.�׆�';�ڈ����?�s/W��D�������Vs�zR6�� Qf� ��!@���&B&���ʈ���;w�q����py)(i�����$�'��d�X��'�DwW��m(�R��D9�Ʃ�,�na3��C�@]��ӡt�E�ߢEǠ#�UV�]�R�	�k?�r�,�G�ɏ��_��DoݢFTXH�0��m
�%3����j�-��	�Kc�.�67��MCގ�$>3Z�X�L�Kn�hK(���.$2��i'�N�P�LZH���mD�Y�Hs��MQ���p�eI{~zĲ�6U:���>��Tk�������+�h��N�� �8��&��'��E��*�JJx�Z�Z"�m�RBt��ǡiWHϝ<d��E+��Ķ�n�Ҭk{��">�+{�iC�M��b,��>:"?.ֺo�J$
��y�P*�.�&���AG���v�˯���nb�#eȌ�4$jB]p��m�d��~}�>��j����=q��vhx*��F�`=i��cmк1�J��h�ਣ�h}��dt-� ��Kr�ܰ� ��H�.O��v��uś�����x�4�d��M�+���7���	�ذVL�˭�D�h��'�í�?�1��q(���@�N27�'2�y�t��o^1��pvq��^�ΰ�n�A2���!8/�)]�P�J��v���Q˱7���������4�b�k(�ܝ	{1t��5w�m���~~FS�ԅic:�Ix�ג���BB��w3���d��<:���%d
�,��B����M����0��܈A+��� QJz�	�GT�3�cA���Y>ኡ0-3s�����b��N�R���|�=Z4-I��ˆ�̸�"�G'儉�DEZ�WďX��?��_��~'�m�%�sKL$n{���3 �(��w= ˵ĜTJʦt�V��P�bvH�oG
��]rB\�=��PH�v9R�t�J>�1���9�~G����Rk��
>����pCw���J��E��hD�X#~��L��}��xO~� �jZ|S��C�n�bU�e�漁�U�kN����Utm@��ݪ�C���˚��?7�?��q�H��`��%J���-�_��I�Y�k�ù�ɚ��X� ��0%�-��_M㒪ڝ�F�:��
܆+"�փ$��!��Ђl؋|����R=�ú�nJ|���d0��>6��h�|��p:��s���e��-DwF�F�O3-����H$n���f2��s��@.Y�t��$-lf|%ܧ-b�Z�L�*�tj���oV#��W5�^Wć|F�%<�"�e���31��鐋R�F|�#9ֳ���� jz��I��`Q}j9����ӅӒ;]�U�=�AˁrP�6B���D>-�Ky؅�,�4��dM����q�o�,��j�[tFb��D�/=۽p����u�&��d��ov�Gh?���v�\2��s�,&F��7VBB��Д-)��-���M�Q�8� 7��l��!QȖr`���d��S��[�S�����Z��έ/�m���ӂ^E�3HuS�lٱ�s�8����U	I�c���1.)�>��K�x��?��ܛ2�ATT���,hY�u0�g���;�]��I��b��bZ] H�Ei���2ʨ��QڞM�2A���#*�����87�x���<�MGx�=U����)���X�3Yk;{��>�٬�|�����,��-WeL�o�	gEf.����6j�G�D@ ��nn�X���fzS�e���in�8]��	6�[��N��vs��Ϩ�I樳�V�������bCS'���3�Gy�R�G��e��G�7�rl����hxήD� ��Ԇf��

13����v�
a:���{��hǷ�ڷ{|f��zh��������,����]lAR�E5Zb�O���1P"d2ݣ�80����< vF9�
F��Ƅ�کpx�O��]*�ȷ�����r�1q�����	��p�L��/i�S� ��� ��:������%���n��p��Y��	��/o�&��'�%�x!�/�'�?&�i�h����`t.�>ş�+�_��!
ua��C��ٶᮾrׁGN�,U3t�3��1[%� �����V��eNv��JT��`o�4'&�!���:"e!B�LmԖ[�Ǖ¶�us孛E��M�k.���r�uw@�����NO��y�{q2�8l���!gBlGj�!�a>_�x)WK��6A�GF����S�~b���gɪ2�E'��0Ja�%��T<��	�
y��V�kyLe�"�W��揁8�$��"��<����)�@�C!�n��
�����/	�Tͺ`4�nQ�Eʨ\冢 ��W����!��O3���yC��J�ympޓ��H~�`#�f�K��!�ld��Е޶68��,�,�=lS���ɑ��V����V�R����\-C���a�l����!a���#����c�2�G��m3���tqR��&�C\`0��he�ygw�������N��z��{M�E����p￡�<K��q&U1w8�Q*���M���yw9o�JU�k�ɑ1��'�j;�+~]J��`l����p�����IS[Y�c�̤A1�7�P�rKJ=���0g|�f>4����!V�����_�R؏`a�^/�)F����!�6�)r���g=��j��ĈB�z�=�C��پWb6m�A�n�<Wyd�m��Fˊi7(u�ډ������T;f�)]��z�O���$�,�C�:���9H����_����b����b���S�D���D[t�|�T�dy#��_E�^~ڸ��覸����YR�h|'T����)HfV�<q:���}߄�)mԴ�[X�\bpe��>�ֲ2�7��Ō}�� ˑ��o�!\鱡b]��l��v'	ۨ/��ĭ.�'��Th����w���N�p�lѤiJB�H4�e��_T��V�mqB͐>�&~�`F؝>tuũ�G��#�]*5������D��M�J
f�by4b�j�C���;�K�AB4+����h�}ՠ_T5bD*r�Ԯp���y��|����JrYC��:Q1����FȞ{}[7֬�^+���K�"r����i��F{V͢�*<Mli�֋L�ٰ�� 	��SΙ�7I^�o��e���n�kC����#aأ��q�LJ�x�1 �}-
�;�`��ZrG�|7�)�S����_d�s���+�G4E�Η���H7%ᓃ 8؜����o�p�؅z0eQ�@u<F���K/���n?��jb����(��n��_C�����p�`n���ggKꄫ��]u5bs��.Z	������ot,�A_J��i�L�.zA�K�~W)E\��W���i�h��=��w�f�`t0���g�7A�=�ZҚ���\{9����u��}>�%э�s�$	�Y�QT��_����s��y�����e�9ÿQ�����?��iI���>��c�%Ճۡ���v�^E���W�B|s�0�_�gc�Z�i�ܺ�BN���K��TW��d�wʤ&k�w�:�w���cu�8���e�"m�.�~�⒳�ʍ�!m�W��~�	ԠU=;���/�y�¾$#�~Դ�ϦF�Gl?��&�������lf�K��
���Z?��fE���t�h����Ír��L��k�p�FHk�r9��) n?sDG�w�;8��0�%��s\$-���� �8�J!v_}�jB�*)#��X��aa�x�`�Kq�=�|��N�|҇�?�tZ��&������6�S�'d=nO�<=k�v�!�������>#('��˖��?���J�����$�{�p`M1��{m-Q�4)~�;(�P_b��eϓ�TC�Y�P�o���*��U{��-an�֖�Z���1��U~�d�_�k (u��92g��z��^�F���.��H������W�/��Iƶ5T�?�z��qMǓ=T?M���%���d���l�t[=��U{�6����S )V�T��S
���J/P:r�4v�9�Һ+,���E*�˽�O��U������A.�c��Q���%�+a�5������q�'�L�e�f��sX��_�,`��K��4ߠ�{�����.��!_�d��BM�`,�m�����P��+�W�O�?�ƪr�ML`�O��M�"(=���Y��XH�9���"XPi'������=OY��cB�@�^B��S/�*�9����1c��~�7���zM�f*�a���k`D����jsm[d���s����@���gngxE��FG��Zu�(�Q���m��Kh��3|'I�N����76���飗t�;|o��v���׬��а	_D��C,dR!H:�S=����N)e����=-R�E�)���1}�2xgeQ�c:�
 ��]���)[D�����7 8~s����H��֞�����Vv���)xk%rn��y�[�g���t̸<9���LB��tB{��R�/�+��V��G8�>j�Z����9�c,�{3����¯����l~�y��,�*�m~��8� �Fk� ;8��:[_�֊4˭��d[pd������?���LKDn�m2�%�~�C����-�)���yǕ�u�CU�_��S(~������3�Cr䳶L)p����K֞�F����M:P�4��J�}�D��B3' }F����}�X|�C�b#Kzת�Ô���ĝEoȡ�
b`-g�"�m�_7R�]�p.��p6=~�E@�7��yތ׻��x>�s���iML6w͉�y�Z�w�x�[y�B����t�c]�M���\1����`��1"f����n��u���@�e�t�x�[g#�R]�<��0�T<��)h&�b���F�Mg�?^qH�2���p��qbyｽ�T��/���J�q�Ϗ�K�:��\��ھ��#4�+G+Y]��w�0|��RzŽC��n��e�픧�؊P`Ύ��)�?���Z*i1�������=W0�gX+[_�X���sx�8";$��Жqa���|՝
x��*��gN�\�����똝����l�/I��b=�Xŵ�B=<�`��:V��c��n�H��r�t'������[c^%���
�s
�y�Kh����u�vxZ��`x���T��S69�<'���$'�u��zܱ��:g��'[�s�:�W1������-�WG��'�IX
��ڂi� ;E�>���u.��z쫻xS�
HY�j��7�7���(>b]����Ӛ�f�-l֧��ҹ�w-����9]��/-�Q�L�@"~�6��ٶ1�{5!t����5�t�:S!���f��5��|EOT�p
$�T����v����PI�l�ʕ���������2Vj���br'2���K덁c�74�@����g��U���Z�v����FwG�%P�S._	�iф�}�_C녡X ���R_�ϚW���֗_��$����d���+���伦�gkg�\�^��
�4�q�#�mM鼋%B�� /�׆�:��!�1N��^�y��s#�d	5=�
b��BTz�?߭1�f�Ӝ>b�,��	��h��ClOj�<��k{�B����G9w�B��t�L��P���p k�v7���~�6�MQM�oe �ҲB����n>�1ã�_�J"�,�A���ֽT�5����1���!|?��=���5nMS��-w�A����"=�t|��$��g�풂�R5υ��K����!���2c x��Sy���-��@��>�8���^��$�e'ڛM0="�X��1����hfi����1y���H�+���5n���+�Z!DӯE��ܩO�����J�]p�z	$+�TDE�FE*���#��A�4�0��̶
%5���L ��{|���*=��t�������<F�s��;Ŷ�ZtcD����O��8*�nL�G*N��]����H�'ۆ_���|��PB�߮���鄳�N�Q:o��&e��(-8�w�Mޢ�}w��D��F���4!t�2N_�C�����@��%rK0V�z�9��J5�l���Z�{�Ah�OV|�q�u(�Q<�W�bٚ>���EX�IaW,�$!����fX��q��X(������D-;��Rw���>h����7�̟�`��ҽ?:ѸA��10�����B�N\��@ԍ;�?`/H���&��ZLb����Zt./psp�� �C�#������5���0^��a<�J�M~=sB���@K�fzV�d�`ӹ���Z|��m���������`RJ蜵�+�u���)7�*��	�]4�
K��W�/�8�,_�SQt�� �v|��g � �	��Ew���r���.:c&�c���81���aD��&L��{��^z[2�D%)"�x�O��!��9B&�������� yM�[��$�I!
�Y����H��"����D>�,�nj!�`l� }2?�Ω4���
��r=�m�ʯ�>�VQz�:�a6�>e���jbQ^�^�u؞}�H�5rC6?"�y���wy1�B�n������)��( �z��*'�v�G�GwL��_}T3�Q�z؊?v����!+g�앣�6�nX�8��M�w�����t��fL��#��`#��KZE��*/��U�bD2�uU�q��u�<�_=������`. Ȅd&�_l��r��������I����8Ʃ�Hc�ҩ��(���[6�Tė�-��w�y�|«�V^���@�e,�p׽�����*�߹�sEq�?�C��1M3�X]����N���A؜���5P>o�RE]�L7	w�r����Jʝ��VP�)���*��}�N�סF�#�9�49�«U
����\ʱ�c#F𽊝xB���z@��ч��+�b�6��G�j����-���Bo|�y�d�B���T�����9�|�})~�z���G�\v�BB�]��2�ZFl\���Ы��B���&͑��W0��_B��qT�� f��Xo����E�nC�9q��LUom�^���C�v*���5Fy-:u�F�8�}2��ut�y/D
'Fo,͇iN��T�fd2�>Z�Nf9�i�`�M#ɕ)V��y�̔��v��T��"B(Ak� �.���� �����j��1e-��}]EN��#��?ɕ�[��6�~�K�=\���>�5ס9Z��-2���up�h��\���]������pUWy����d ��@�v�r�M�[n�x�Z���#���#w�K�h�H��|��j��
W��������u̇X:��YHuG�>m6q֥���p�z�^Pv�qg��4aH}��������!��1���q�"�ZtT5��	��v�b�6\)�q�h��2�4?��~fn�ع��/9��b&�O�ݬ�L^Z\��1�T�G����ޔ���v���n�:`�+];��[C
�i%g�8���^(!X󔑿�ྶ��`��ZaJ3-���n��O�F�t��#�����bw7�l8�@�珠k�G~(�|"+�����X|2`�;ݶ5��v}��2<��'`�rz?�B1��	9���[�>e�
P���=� Қ4������0�x��V���Ɵ�'��:�)�
r��%t�fq��X��o����x�rx�R:lg����C��d=�[�p0Ǹ���g>�����|*�F���)�#�#�^��T4\۞��	���d�ٶp���u��=�8wI�Z��+�''�L��٫�����m�$jU�kZ�Wb�:��W�cd�E�땡So_��V�9�	���B�Ig�t8`hv�������R3��.n���*�
���\.�iW������z�=��I�-���
�*5����e�����������U��ϓ���[��-��{�V�wd�Xj���d���<qG��瘪��Gw�^]��:�o�`?�.���Td�8{��)�v)?s���	�:P�#/^֐HAb�I���
���h��Uv��_�L����B�)��t�F*�QѸ���f�-�]��t�� ��wYj�A[GW��*�5�m���n�Z���n�%ppW��J�?@sE ����32t��*?��yH�ʬ�uO�\i�J#���,t_�P �S�"�w��|�R[䔔8�O�$ �U���T@{�h�����2Ҩ���L�]��I���u0�yQ��0{2���c����f��V�q�����7����˟��Z���y(}������]��1|6�?Q���'���%GB
D���i�����R�>TO���f�H�<���~����U��#u��h�/봑�*�58�r��&�/�kbˮ�����e���V�*C�]%>,�fh`����sp@�ho���ћ*Q��}J�]�Zb+5�����:$��adP�vK�q��1��͂h�P ��e!2c ��������.�����0�*'l��N�����D~�n�X��z,�i��Էl
��l�=�w����:��"f�ɯ�t
�n������>�et���t�����4$5�hsB��0�OCߖ<_��~��IV���Fզ:p����/y��ϖ��� K��l��!o�AƸ՝�
P�"��7e��aq�ip��� ���K8���X��"J�A~�R��.QUC!i�])��I��2�,��S�(��~t�Zwd�up�5)��Ce�>Gd��tk�6��N�k����v�n:^'/G@��c<���wH�CBr�WӪ�l۪�9H;�ǈJ�O�+���{C�!i�ҋ"m�]]����Bm�s]Q�T6"�cr���h�S�]���,Lp�S��B=�OJ�q��w���|��*p���D�����@�v!*��J3��R��/V|#��K��@(%��?4Ĭ1�Le��on01�g�w�%���	�J�v�L��|ށSfGX#��Z@˫�+���q�o�ff�q]�NH}b�p9@=arדj���i�*�t�`fo���&�<h����2 �F��YspNc�M�;�b�\�c������3�l�y6Ud��\pg�D�y=l	�F�y��T؟)�<����K��]��6�U�q�C�څ�$�i�����U��[�����Vq�&w��� �k�s�v��`�DGǯ�o�l�?@��K�4��`���jd7La�}��� X�P2I��T��("Tg��c��i�Z������]��۰D5����������g_��HOdj��M�˫XÄ�Oۖw�Qүxd�� tya����w�dp�H<&�R�v�%����������(^;�:o��|m��������)�7Y�ߩ����M�@���E�'[�O1��R��8�>��ix��|�*xN�Lؽ�)��,�.�+;��Z��vTb���mV(H]�tْ���K��k�7:m�+�[˃�1�)����܏���n���}�t�n�k����vQ���C�<��7K|�_evѵ��Z��Ub?t&ߒ3�Fڡ�h�V
�q`¡�*���u�u�a?�n��D��Ϣ����yF�0e�D{�slT�
�BpKl■$&`��z]L�(�I�8 ^��I��Z6�ͼa�BIAt��$��~��@t�(��X��X&�+�S @H�(_Hر
A�M�]�f�\;lڒ��c'������\���� ��?%�~}W���x���,�ņbS:^Y��ѫ�%=�մR�-*��y���!�>D�?G�;���k�k��ڿs|�����B�%V�y-^7��9hV���$��+���&H���*]*��H��Y!ݘr���	H��5·����ӚM�b�{�7��O����	c��>�q�R�����}��|
��jVif��4���$����}EE}�����P���|�t}K�� ��|�7�G�ӆ��۳il�\�嘍�FQ-���G��דq�p)"0}l���!�	�4��N�ﾊb�*�`/5')J8Avb�IV��3�﷮1�����bb�*�,C�K���O�­��G*�n����j�2HC욚CZ��B��E�eM�Θ$*GDY�7������� ��ܼ�q���|����	>O\9P���S3��,[��F�\� ��c����b�H�����~ʬ�@��J�����L��р����˝�7��.c�(ڸ~5��JT��o���}F@W����������B��S�'Bh����l;^�F0�f���l�Z�,׺D^��K�-�d ��4���{��y�`����)i�q'%�r��9�*��w`�VX����WX:�1�܇0���
�e:�-88<�ϪX:�x0�늶\���w6м��\�=��z���}������YU�6�!�nNfw���<�0�G����3���hA���/�>���z8t҇$�ޢ���[��g��N��%3�X:�i2��=�W��7Hq� �k��B�
�%uNM5̏��O����w��?]��]�A��l���M�gq�� 6�+�]�4��rpbKQ���'�����ڦ��B$��jO�o3�L)�_#�$��Ѯ�R�j���@Eu�c����A����\���H�NR�ome���=�c�f��s��'�g������a�����	���ťuf杕��h�"���0w��n�@����
�w8�E���|����8�8q�'���A��X��d���̠���7I��ǗO�Y���lM����pH�}���Q�'�@wR=�1F]��Q�P�fd�p���0k��9>�}}��4MR��	Fެ/��X� ��PBx=.��x6nsN"�5@���#���ƥ�c�OQ�d�X������� �M�U�Z��6�����͘���QӴaTdm��gi~(8(l0�/�䉠��m��"�:��?dՍ�܎~"�"&9V�5��E㝋��i�HĘ�aP/��όf�+p4��h/��gDx#Iw3��/W���K�,�>�H9�������m� �[���9-�|���-�U-���Q����m8���`S��(")�۠m����(r�T��&�A�L�( ���\�jJ���4Hvda�����$5^����r�M\���B���Kp��,J��a���i�G�
d2��[�(��� ��T8�j���7�^��ۮ���1�rw�E�μ�CHF��a�5-}��5n��$���D!t�sp��,w!~�#B�V��`������t>A!\
���*�֗���N��/Ͽp�)����Z߶�AR.���z3N�J

=@�'�φz`x���-�k]��+W�š&"�j"o=�|AS�nzd6�~��	�F�k5�Ⱥ��4Z�]ҵI�������+�Y��6M����a��U@	���ZA&y-�Q5���V�ylշ�h���������T�;��<�5�����\�"
�y]��I�������Y��ܟ���r6U�3֣�N/�1d�,�J|�$s׭������y�[�]�����2�K�A�l�a!������~!�=���j�M��13�ݍ�Z�~�)��Bd�^Z����U��p����N����-�g��l�}���h��/�,F�SRX�,��ǄW.m�W>�X��QvI��]�{
YCY�ר��--��"�8Vh�����+�����N���
��='݌j���kY�$��a�;�����l�:�ԝnDx�R��:dGDDuֱ�N�\�/�|$8wDO��ە���%�UaS�	g}�
7vC�ζ!U��;�����2��T
�� LV�R9J�g���ɖ3�5�����{��6bQ�~fT+9�C��9�+E#�d����6�������2�m�5������z�w�j������+p����bki�2�u�Q���X��p��~��[�:�h/�"�F,��L�/��R��wH�tߊHA��Wͷ�=�T׏���d����H���w�lC���nJ�E��2��F�{���&�fW�I��Z��!o�d� p��g���m��U|��3�a�����%�#쒒�3������H炩�t���m*-�>?�O�T]���2T���F���$�I@1���J�F��j�g�H��pA��,���ս�(�>���z���9�s���"�Pb,u������@�"����F��m\7��D.�s�*��ӗ�t��)a�{���_�vN-[�9���0)��:�^��1m�v��l*�v��v�@�&*>�-�PvA����Ց@�؛��~DUdK�=���an��%Ӻ���{:z�A���9-�������x�鮮`�83ѷ��̝��{N������� k ��"Y�>� I���T��f"/5J�e:߈��ծ�f��ڙE�i9:��h4��.P�zc���C���9~u$�P��V4�ֻ}�����W#mq����m���zpP��ef}�(lu=�f�A��}��T�U��	!*��0�����LϋήM��}Ǐ���\�w�:��7�� �C�_�ڊN>��Z�����Gfu2�K.oȲ�O�Υ"P#�/��6����u9Ķ`;���H�#�s��=22�K:ՅN�~PP�χ����;���G�R�d8��'M��[���M�``��)����S�(E���ǭK�{��y��'���^��p"5p_l��c`��(#gR�5�#E���.��	D��y�N��~xm��a	�a�����]��(@�ѿ�hM���q�=�NU�=Z ��������y͹'N�aYl^ðV�=��`K��
��fo��ms
G��C�+c&sY,�Rp�����)�:����q�Wk�12����f�����┎z�U!��큌w���l�\0�5.tX�p���*�{z���n啫rhh_������#q`�Y���}dv{�W)v`(K4H�>!E �3̿��a��Skc�ȔLR����/��$���ȗ��k�A��Ԫt�U��D���T�(��ɛk3;�s��l����wn��h땕#�B��G֎�����'�%5�Z52vW�}I-��"�/���ډ{��(�Ex6�����Z�τgl�ų�l�iQ.���4@���
,L�6fb.���Ѿ��L�$*�ٵ}*R�W&��9�b2?�"-����=�0�l�H<�O1pN	��Z�r@����u+@�(����M>ל�[� ii���i�f������;n,�v^�ɏH���!e���^�G¼��,o_����A�~W�4=�+�O�eȚ��� �__���G�D�]"��(��[�1n߂����B�d�PK�;Z�z�e�!l%4�~i��(�(9U���}O�°���1ykgS�)&���gZ�P�+"4��.�v=Ue[�o�g�xEk�*A��[�������(v}�+����$Iy�D�$5�=)��'ޭѲ!���2�2�"�f��^��OH�)�|���U^RF>�*-sJ�~�A`���a�
�.�^��Z����_����Yl�B�IZ:�ݠ�m�8q�@S2~s*D�g�i�ɓ}�i�?�7H/�=.�5��.����-w�7�܇�p��[ᔥU���VR�T��x�(HQĻ��<٧�뺮Ȥ�8�s\�B̙:b�M
�db����K����T�0�u|~U
MhrV��I��9�=[z��> ����֡�����2Gߛϱʛ������9H�ϱ��ph�]޶>	I�v>3c���ϟƽQ��k�E��@�D7���8x�If���-&6Ǉo
��!�b�� LL���7Oޱ����~�$�,7{�8o�谀���+�`,n�qѻ1RCr��E{���3.�r�G��~�>�7��9{�[UyW��I� eoS/�q��B�V��Q��[��������٠�R�(��~�g���=�(-��Ũf�bo(B�pT���6C�z�9jˌy����e�����	W�WZ&]�S��D!�������"Qck_Ց���K��+̸�y1�cA��N�MRMd�c�VťP�3\�&�b\���7>��FV�t�O��3�*K,��`�{M�Ůk���&��.^3��0�צ�U���ǐ�j&n��F�άV��(	Z��Jq�b���?iA�ϻ�R��[��ք�C3>d��aZ�A�M�I]���N;R�R�`vci�"��lTٷ^
�z�
��ې?-D���5@�o�m��<���a0��&!24��K�v1�m�kuM��o��2��퇺�ʈ�_��4@(�H�m�:� ʤ��ft!m(�ͬ��{�_1��Ƥ�LbB���/�!^*n�������ι��r���)���&��6$�8/m'n��ۅ�͔r-�a	7sǴ�U��W�=ˢQ
D�~�P�u�rZ�&�iF�����e�ͣ}q�]�ݒ��e�P\ĦٰD�������@���5��!��#8a�vDQ��4�bt䈁"�`0S~Sc��G��ZqU��e�]q�GI������m����bU�����=��4���ֽx��Vȉ'0Y�1����ڢ�7.�%�R]�V!�e�㑿�6l ��m?�>��eL�-a1=�rZ�d9�����G�S�SC�mE�}�����2�%F�0�czv_�X]��#��!�['5ظ����dڏӗ�3v�my��'y���RDs��l�����<hxz<�gE\z�Ev��n��/�^q{P�n�54����p��Ñ:�q(�?�]:Z1��of�Y�z���9����svE-���9�����\ �2���z�S��۵MK�a��4�Gy�t4;á3S��P��׋π9���0��o.M6�Rg��۶�M��w.��G�)i���A��ȑi��uk��N�3u��u���L�-"v�zM=Q��.�BN��;ԏ�y�yva���0~6���.�n��_��^���S�-[�&�V��MD"�H��U�RI�{���2v�_�>V��¼���f%{�}�ǹ�歑F�����.*��l#��d6h�c�@Z�e�*�%e"?X�:���;����}�ș$n�t�w1P���1-�*E��ys3I��sA�۾���]�Y�j����a[�X	��.[�k����q�R���^�ςK(u؋'���"NK�s7�JC��N_Ǻ���Dܤ�5��?���ٝ���EZ8g���/N�{�{Q�X����80
����UAVjS�۠d�=���($��7�,�_�̓C�ySmޓ�- ]�p�I�e�
l�_bJ��؋�q9б_J�>}+��N3���/�i�V��'��z�G�j<l�٥�Ul*^#��]]�ŗ+��prw%����F���	�eo�0L�j�uh�o�s�f�B����Y�VР�c/ u���XʒD�y
>�P�5� ��:���ے��@e��VnIw��"����Kv������/�C�/q�4����:��\�Ių)��=m`<�ĥp�XY�����F����r�	a��Esz2a �P�snp��/qD�Dnh�Q{:�	��V;�F�مN�3�W�ǟ	�&��DUG���0�;�5�׬�[�,��GJ�$!��r�d%�|߱�e[�G1,xLJ&&z���̗�<qt�P��	���L�����R-�%�>l|3��f����#QS�/�Y��_+%��22�a�����ɸ��2�S3�ׁvY���es�}�׮���4��?�g�?5t���J�Cl�P �1��XT�,�Jz�����ؘ��j�$ȣE�����UnnD<�Fq�B��M�y�8�eX�sWڞ5�ˮ�Z���� ���.ש��J��e��۸��(��ٍL�B�eÈ<�屣�#�Ϧ�*����V��\�ch���]J��Y�t� ���v�\Ա��8}�_�n5[@���V6J:~�nn%[۷=��n�|� ͹�t�s�S�1�RsU��mr8v���E�����;��H���1D�*����l8�q��v�e�ѭ��l�#Dyz����;.T��jM�N$�6q��m9���� �Zu`���V��.�O1]-7��r��I<tX��dM>�Bk��*_��큈��˲�7������E��Y�P;��Σ���ꊢ��E.Ï}�1��"l�W��3�y��j(Nr	��F\d��ɫ}�#}�[�~ېT`�T�^	�&R¯y��5b��Q>M.n�1���60{4s+�tauP��r���r���u��J
[e:�$���=;�q���!��

	"��H����(�c�E�~k�Kx�����^���[���G����wX�v
��	�فϺ��FU,KBg(����plc0 �C"3���ݍQ*n~U��4�[h#�+�y�2k�Np�V��1=�,��Μs������d$��_,j�=K��,'�M����1���*Mx+���7�h�L�?l䨅�+�b�r�9��8Zz莿 �Auv%��Z�J>�z�|?N�ۜ�u��0��}�1��a���BmB2)��������\
�y��w"<�4`n��A�Y��Z�C7m������!��+=�d�v�>��&������ۗ��e��H�u�*��(�dޅB���f9%�G��r�a<LV�� ���ȡ�ٟ3�ˤs��[��_��؄�E��䲯��@�Zb!=D��_iW��n�V& �1�LT�G�m��頪 EHM�����t�+,STm[�j X�=�,
_��Q�z6u���VJ�+��|{�$�K$v�����X\,-e���7~U�h�'d��/��Z��8�����Ӂ�4M�į���l�P����
����P���&���
�3$)9gfR��1�F�UY�ԖyɜSx8�/ȧS4��Jn!S�؊>����̬��o��K�Y����.sq�%�}��~o�����V���s�p����F�_}1	}��B����"�dT+'�!����yU���Y����`)��=_���I���'��Ŏ�|s�J$�Qo��Xn���J{8�gd���d�� Һ��tk��y����6i�#�H��ט���Âz�,���G��,"5�~I�%��ǭ3 fW��SUcU�@��m�+��Jݽ�~�����%�*&fG�6�D%������4�+�y�M/=��<�aމO��g"� q(�}�u%�����M��1�ym̮m�m�� �Qm}����7����jm�=�gym���?.�T����.d�6b2kn_�q��p��nl�Xʝ�������z-XZ���3��*
�w;���<��9n���+��jP�w�
E��W,�}�|N��q�o���������	����,p�����_zx%�08R�n�G�Fq�WsfIPha� _ge^r�)�Wc���{�g�Z�Y���!�谅���2;�b�85W�w
J�bJT���@��m���[ՅJ���f����v����Qm���R�
e��<} � �5
��td*b�NQy�]i�5�Ƒ�o�M;�8!l<�$h1�HʰN��$}nn��8T���>�3��/�WS�6凒!�!���t��tp� i{��Z�����߽���,��>4r/!c�cQ���ɩ�!"�����Ě�7��|a����n3��n�w䗨�+���:y����ͅ���/F�R���P�����sl;���;�s���@!�`��@0+�� kF�/�0�X�,��R��A)q�K�e�Itr�*DGG����JV�	��"�s�� ��8s�O���hei<�{oJ"�e'?G��� ��� �
Q���Bڊk��1B��O��DE�GGY2�����h���II⅚ˡ�>��NV'�|��*A�A��C�ɔ�KxE�Y���Rm��x��n��5J����\u8�V�) �+�J#]�09�6���S@Ҡ��-��1GhPK�ރsc��7Z�cN�(�:��T���{�gτQWpS�M۰�@Р����5���Ĵo��tܱ�SX�E�Q���,8ɺ3��:�ciz���o��`�(�̴��B�K�Jv�}w��Шljn�����Вo��#�^�3I�|�'?�|�1M��k{%����5��7����`;p��떜�E'J��+�ߟ�E�V%>q6I/�(1O-z�/	#�[)Z�����s_l�]X�{�� �\�
B��Nk����"`��$�a�PKS�����D	�W~(
�6��m�ذ�,�{11��1��F�?���A�ʫmFg�NPL䂱]�'���N��52/ոs�J�#�X@��8����Ph-ݜ�r�ZH�3d��ttX�����#b�3F��-&ЙѤ5,��ٌ>{eb2��R��玤3=2��lѨ�X�-����X|�
�	���A_e/�qh��9��<Y�Uwi�$$��G�K��.w�.���mHT4�0����Q�>�dnN+�~l���x:ۊ�H+�h��\�\I�����:9|���+ak�i�\�Č��U˄-��[X/�u�!N���!�ԇ�f��n�1���of��2��'�Qi¬�L��Pa��.�f������~C�I�L�H^�7�o�i!ԨlT�S.�#YY���N�����v��b����k}`�)���+E����Klq\Ù0��q"��E��7��I�y5\ݲH���*�ztz�A/��
OB�CV�7�N�8f����}Yo�@�f��8o`��^d���P})AC�kG41D�b��e[i��*b�"CY*rX�Pz�[��p��y����[�6���O�������o��6�~�D	�� _����څp�\���Z��>ʧ~i*T���/f|JM7�Y�D���c�g,��&
-��AU�ʚY�
�A���������[n�$�B]���!>�x;��P�;�BPq�X���eXk]4\:AJ��Z}P�?h��e$�����;��5���rD�"~�2��U�Q2�!4�����!�:)h2���e8&�1Yizzun��w�|��G*NMM�DG+�c�	�,�ϒ�W�����ȋ�L��8�)��M���t��S�h=| Ij�e��CE.�i]������還��P����#i� r��!��j["Tx�Fi\���ڮ>R!BX���篷���wawC��y<��>�_Lv#9�-׾/M�(�Z�+u�H���B��#ur����4e�{Ae�	h&��_z���>I*uI��!^R����*WS�ڹ��f/+��= �	��MBD����s�����Ϥ��"��׻ʯ�'^Ц�8�G��mPڌ�����JU���o�o;�����^��BW5��pݹ�+����1�Y�O�@^hWk|��j����<4�h�������/^1f>��L��k�����3C���y�oJ
��%Y���`�+�d?��`�(�4_�hǜK9&=|�r�t���T�m����l�c�>&��8�D�� �/�Z�b|�kE�4$@������g�͌dݹխ�V�X�X�i�D*՛�
C��([So�bH�~0�c2=rJd�5P��=�qG[��� �:�k�����{?�������D�K`�PQ٧�WG`���0�^Lq��?~;r��TC)"$�>u�L4J����ŵ~e��ؼ<���֥�vʎ�'��"nVo�}�k��ť�e�+c��z����z�p||���x�B�<���XT�qd�P)�A�.��5b��w�8k�;����p�S+Ȝ͔��Dԍ�pɨe�(��3`������� ř�_�A�%�c�|�2�ճ��j����&l#vo��8����vM&�D��������ͼ�0Z�A-�a�Md�� �;��4���w�%���x��Љ�
�uroa\���)���Ѽb<!����套��g�K �ыH�C�s���`lU�&*9Q�
�7���`��8[�.8g!�+��ٗAt����	g�%�*$�<mm;���},b0B#���o2�0I26�_cX�&�X��BӤ~��Z�U-�{srPm�
oU%�^����R���QU��Hr��;۷�s0��n�
ѵ	#�c����X�0]ZUV*���
��%1���_�r�JL�ymW��jßn�z��+5��1h�ӝ��֤Fׅ�@g�~'�ع�� �:h��&s�	���:!���S��|�H�-.��h3V6iYO�09H������b��֣m��#�����4c�F	�q Lf^�)��Iyxğ���w<�4�$��Z���U��ȉ����$���1��1Kj�q��Jy86\~���r��#I]�������ɣ| ��������{?{��T�Z1�V��L����Zz{��b��݈��������1�{�T3�._S3(����eh�jrR�n/Cʸ�e'ˢ*E�H��z�y��E�����,4��`4���ర�k���I�;o��<�g�UR�Rר�~�[I��F� AO��;���u�H"��I�����N�%n}�nx���|�����[mw7WEm4��d;�F�8Ku=��p����Nܪ�E2�|��w�۬�j���.�(K�]hj"ؽ�z1��QSǉ��6��	ѻ|q�����D=����@�ܵk��iS�`���U7��n_�u���R���2��m�"��$V}�2h�ہ��w��y�N����I)�[*�iYα�-�P��-�����������M�PnY?]���k���O��DU�����f�C���~��4��h��}25��ux�Dg�.�rk�El�bf�+@SuRF��:E�p��!�d�������5g��T���	5C�6ASKzvi0خur����� C�!q�KP�fg#.���!����}���9�N�{¬jxű-4��{��hHK�X6މ�:p �w�,�O���S��:t�����ˬ1Fg��ݢ��#$����YC�@�=7B$�a����u��p�쥩����H�ҷ:,'���ҁ�������h{Aޛz�,-Ά������Gi쾾}f�J�#T�@��5���1�.�%�A�z���C��r}��*��(8��]�i��7x2Th���B���y%N���%�����|�T�u&�,1�i��R?���h�����{��I1r�� �-N���:,��"B/xO9����E+��;��GO/�!�9�������*X��w3k�(#E2Sː��2����΍e�z˿�_L��5�ՐP��@�#|�6�8�c�x2 ��d�t�3-(��w�J~{���+��/۫@�)Z״`r@�e���ԕ|������8�¦�|���e �z�C�e�?fH�<���DH]n�>5�>���l�C
����?>�<������#��8ecP�?q.ЦbX}\�S�����T�O�EC�\�1�Ҟ�0#�f�7	
��)u{�U�j&�?�����l�q�-�$��� ��V�s	�+/%=����O��hH�b"��eH2���J�5ɗ'��dlI����b+°�:r%��+�zZԵ\�h�Q<�T�hk�W�0ች���]D1��c��L�y'|��	�'��>\�9�w=���tu,�$Z���������'/�<�%ű�q��8܂4�ӹa�ǫ/��L� _�!��c�0l�b|@g���<�`�^��f��"��]f��G��Çi��S�K�sj���(U+�<���H������Zm��݀�L�㞡�΂����0�JNp»LL�_C�֓c#w":׾ȿ�2����� �SGk�Q%�2?i�ʔ�O��R���6�@)B�I�|[.Y�Q`������	L5��O�`V�?� ��Z\0�i=�<ܵr�Z���r�P�Ņ�-�ѿ�#_������{�88�E���&#��}0$�5nR�>q$�U�dK1�m�)B�=���ۀ3���-�;~Yi�,eiJٕIAa���v=�,���B��yG����{�4S5YQ�&Kۜ�<73B�?Z���*�����O����G�y߅h� �q�9-v��K�j��>�,��c|�̡͍X�1+��ʔ�m�xlfP<���i&V�&�B36���wx���ϏX�T�ap���q'x�B@��M�v��4���
�j4��!��� H>��_��3?~j� ��5F�B_��#��j'T� �e-����R�>d#eBl�U�����8�*�z��t� �g<���e5 Kv_vi�����[cUҶͮAKB��;�~eB2�}��f����Oib��ۑS���h,�淛U�Pn4G��tU'�n��B�J'G��kO�-k:��n��&d���������{��)�����7��������M�&9�>Lk�f����-����z\�����F���m*o�#gVw�4�;�<sB1tz��T���R�B mL7�zٻ�f,>���6�O1��e&��AĀ�Pڪ�� D�]�pn�&J�P��.)ʟ�dzh����P��z���@�5��Y��!Z����h��=���Z��P�Z���^s!�?'C���{܌�	$�������];��95�ƈ9��9��Y'��ڹSх���6ޒ���[I̙���tkW�TN�dW��"�<�p��S�ѷ�bA�슋!
���4r����9�	ZH�b4�n�;���H���>;�.=�l���Y���Q�ks�--a�e�X>��q�.��e���Zs��,i�h���G语�b����e�5Fz������s(F��$�5ۜ|�<�6�#6��������X�.���c;H���%����ދ�ڒ8V�ԕ]��6o>�S</whrW�p�;����8Q��w.ж�/��q��X�_*f#�Y�Pm)�~ԯ��vg`�|J�
O1 > �7B���j��.�Ё_��RV3��聕�δ
����I\?EY�]�� �4�.��2��B�o:V�y�yJ�on�QV$�u�K� ��U�����SI�y�����l�##�~�+���T2��� %�S�
Z�3:E/)>��������Q R��;(*�Q�x:UL��5��`I�;*��,d�0���.A��0z$5��)ę�mX�aA�e_%�\�xC�?΁�����4˧����'�x^�zb��?������Wo(?�GqK�W��aY9���O�ª�G���T ��[����W�-�!�Ae�4	�y���C��%�a��V�26D� ��K��C`�,O/����=�t��p��0]p@�R�#{��Gz�PP�h�4�ݹ��8WSNG��q@���@���>�C�Έ��ce��-���*�x�k�3Y�/�h32��5Y��6�#�F�=ԴPׅ4��J��ܰ}�3,~���:��0`��Se�1�e�A��RWў k�9���c��F��S��	��TҼ���MG��PV�tKY��uՄd�ꑍ,�P/�9������\��.PN�C�04u�W	�֐���M�޽���1��L_�s	�]����K۬a����r�᭟3�hwx3$�T�d���K0"�l��ʅ�Qj�/�FM@��Cۡ��\�3�9�y���N�BX�Vj�z�3���+�EI�bVw�u����ސ��Ф�t7��h�ܖI��x�M�����{3�ښ�^���aD(�|3��+�[�9����[@���X�Ѕ=ұ��<�H,���İ���Q�p�ֿ㟍�"JoJE���׃��b9�!?��jV��6'^���g9	���4n��{#�Z��2�3$^�tV5�|�:�9���5j�[��������Rz4�"Y�$�8��J�~F�,�tT2���\���IY�{}�٨"+o����%�zد��5��1�Ֆ,��Y�X!��RO<
��bޅdׇͮez�ǝC���*lxp2�P�~	������Q�V����#��8Bw�1]N]��m�e�B�b�^*5Rr��C�1��Un�?Lu9��?����;פ�,�#V���xu�i'%y>�$� wb�r��ͮ�{�2�\��{�5�\i��#���ɬ�5*�j��NDY�R-d4[�Hm���U0���g��`��h��i��B�,/sUӞ
�B�DM�Qh��[<B���^�~�-/�}I�؎GJ���R`�AN�J���)q9)���kޖ)^b�X�-�9)9^$!���//ҫ�-%c˜������/��/�*N��d5h�9�%W�y��J�X��U���~�"��|�4�fv<��~�64�-%B+=+��g�)���{?��KYȶ/��<�Y��g:�0��Iv�u�����K�G�E�k$�������dk���oR�������9���<�������<B��H7�ώ�9L}����{L�RWw�d'�i�A������;h�����k�OuiL�)Ҭ���q�V�8$�$}��a�>�W��c{�ų2���'�Dt\`FNO�#ջ�m�/E�1t�+/��R뇛�Kv�@(��7E����ݯdw������KL����I߇��Xs��F?)`��/�8�#G�^�㖼+�i	���!,�h̝/��)�u����Pv��i9~���C�Z�mY�g&������\䪪�O
~txrĖ�`�5ngM������Y�?��s�F��"-���`��a^c�a���w���նT�aG8�ק8Pv�L�yE#�N6I��@.�/��R�����GU{���"�/�{F9Kd���=^q�Өy؀����xſ�JCSb���RV_&�G7���W�p��{�������E�}߻q492wd
0U���U	v�0��`B�ph��^�e+u|�6�Xf"���IC�0��-t��d��h�������Oz�!�v7�4��b~!��N���5�D�Q��N������B��<].��:�r�E�*�m�ߍ�;P��9�Ug����5>G "���m��	ە�&i��N�>I���bE7a%���2�ş|����_Y�K�����7짝��SM"������2�#W��v���$��y4�� ���5eA���^^T޸�K���ݧ����8�T�����<��_3-�����~�YЖ��Y	}��
�!!-|�4����҇�@E��m������P�2W�z��[3����\=e��9Τ���87�
�]��I��P	�%�5-��}�Ԩ�#����XuK��CwҭnO���ƚۍ>�*cBo0�Lm�����M�����ii��6�2�h�L~Z+�^Z�YU�Q!]�ܼPMoE��Tu~@n0��`�4e?C���-��DYhv�y��ZAT��B�m.��R����r�K�a+�*~��n�8��^��쉂s�F�����!���s�W�w_�z��-��{��	�,Q�B��]��g�>:9t�p+i��E-W3=k%�r׌�$dh�	Pl;̟ذ�]��
I���nzz���ط�z+��]����n����w"2�Wֳ �4��	I6yaA��͖����cd8u��W��8�{2�����h�R*��ɚ��� O��i�.J����4�%���F�1\D4,k
�G�����X�n̌�s6弲iǭ:a��Ip4��ρ0�~�AyZ�-g#{)�QI��������z�����|�g�_����,��h'�W
�wʧ0^b�}~0���~7���W KU�H��O�Ӣ��"��Ċ�e��۵��}hٮ�r�)��Yr����	q��n��.F��P�&�0��jU�V`9�l�7�����3` �����t����گ���k��g!ѣ��gO���ڦ�h^��P[���K2S�������'��yt'����h_�.�ǃ� m2��~]D��T�uS���ױV党��~��
Q��G.I��[V���+�A���R�\l�TwJ���?���Kc��B���.*��%7�N<���D�^�=�a��6�*υ�6|*�8���{�vs5W��j��U�|ٺ�P,�L�4Z�ĳ���)��;�r��z<�vلQ��Ǳ�4��
�(e��tup���ۘ�*U1>���M����,ym�����F�)����A�O_9}�{r�yw�[������)�~`'�.�u^�_�z_����ģ� %��Gb�.Ax�;i�#���#�"pOu�����67��{q����6�<2z``��� a��r��r���W�"C�e���nT���n�G�RނJ9�@4#��kx�^�C*���!�ڬ=T?Hm���u���|W�կS��	��^q�nEK5�m�A�����GA�]�9!D(G������{�R�����Ē(�l���.��{��+!��w����RS)�8^yH����B�J�{��[���R�
Vd�Hf�ׁ�}�h�U�������Ύ��L��PZE����'�7tl���d�_�:!I`\/'��Y��-(fX���wfò%��H=�+�N�ֲ�U��B�u�B��㘢7�1��y�8:�����qN�2^���<�8/�N�Y�}����f�6:���P��Z���~͟���i�̌�⬆\��3`q�����b����	�mZ�R}G�:�2��N�D�msA��X5���D{U�����!��n��u�W��r� N#��F��t�7ԎM$pL��ǆ=P%��R��4�ϡ�xօ	7 ��x�)_ǌ�!��y�]JR�+�m<�M�*.�d	�vt�|��E�o�h-��㰩�\���'B�����V�	i���Y<�$7	��<�Ɏi�լ0�2ѿ~L5�Kw���(�rX�g�J���n�.#D����A0�(P�E��[BŸ��[���.��;ySJ����:��^��0G-�P�'�W����P+W���x/�	{zn{��ޫ��BPW,����'���yI!N0ؕ괚O1�MB#6`�҆�P>���V�f�D^�/Ї[���p��u/�5v��/���R�}�;!n�,��(�;�Pݿ �h�~^�:����Q?����Tu�$ܤ�ܪx&�Ç�P��J�^��"ia#���(W�����ʿ�
wy$l��Kc�Ao��*�7�H7�y��Q�R�hL�mo'���BϚ�si�]��cƅ��#�>9��R5�~�
�$��BZs��G���L�D��8<g��j3+�E��g���z�t�����YjI���S������N¿�(����j��u+j��$��������f��򰌉�[�Q��յ�(!�X�L�Mt���'P_;���Ό��?K�!� ���F�Fؖ�ҭX���yIP�<��
a����(���9�Ce�qК���~���3�f�*�5l���O$�G����q���G�F�����@j�>����6�����q�"��#�����粲O���_-��P��`&5J��:�3&i"��ۭOE-��2M��yi�#\����p�]�3$
=�v���*�ð/������L�����US��J�����s6��:�@��@�m���	Z4#�Z/e��ӳ�tg/4�+�3�1GZ��|-t�"}���P�i�eF���� ?�� .���/�RWd���N�i��7\B�8�-Qb�|`��\Lތ"ݟr��^�����W	8c�#�����D��cB��������ku����p��x�����~�"��8�a�g��Ia/ılm>pv���A�[&>rg�wA�W���R��}�#�M�#,O@u�s8ƍ>@B,�D����Ƴ>��+����.UI��^
̕�9�5^r�� ���o~0��v�,vG�������-]<'e�-R)ab�$E�D\��릸�E$�<6�j��c&�7_���'<N���1ːIr�񐶔�{<؞u��=�P\ņ�7�����KiS�6����q��k~��8C~����a\�d���ȠN�t��:�R�0I6�����_�s��V��E$�P�C7t�����08>}��H~�����E����[�$�nt�y��dd�D�7�j�
����E��*�Ѧ~�G�&�BXV̘e�����wV�ϗn ����ur���d���������yf�6�}ԃRg?�f�ͣQ�4���o�.ׅ%I��e��nG����ukj��]��7���|���`^3�]rS�s$*,;�<4�a�½�ȔVr��yQ��}c�zA��L�9]��K_2�ʆ�f@֐�0E�������gP<��nĨ�u��"J+��P�e���\�x?��pnSh��W����?> UXlR�E�	 #[�K`kݘ�X�pz�3�ܠ^�U_&,�!�I-"�̈́�(�'����@�VQ�4M~C�w9sDN(&�o���T]sѴ�?��3t(й�u���J�W��VW�گvR�bHw����X�z����A�k9 �&��\�����Z'��H� 5���u		LH�S�Mi���W����Z�j_5�1?������$��8��W7�<�!td����� El��=	LE3�%8$�'f��Q�d� W쥟T3ł	���)�6;��3�#o7ȗL{B��y��1��5�ũ�W͘�Î�OU$u���͘�쓴Ұ��)�x� �SCa��N�j����5�?�/46FhD�Mͺ�y�߆���]M��n(�3���ɂ�6g�#������'�u�N9V���s/����,6XI�y(A��U���"17,$5�_��a��%zߌoT�ɏ&�ئZ���w�y�$�Ǫ`�D�=z+�M���W�{5^�!�1?B�IAX����ӷ��#�V'�,����'��Xcf>8:�nۨ;Ҙ��O(M�	����ED\�;\)���$sZ�����wЪm�PZ1A��)!AK�����5%�Ӷ�����BA8��6A����#�+�X�)���m��)?
H�9(�k�5��*}�gP�����F�t��4�9^��W��@r;�����B����w�HR%�d�h��0p@F7��Y"�( V�i������	.30��%��d��*\nɝ.��v0:�t$��gj�^^m:B�G�C
�����9��ڑ]�s�1��g�#�v0�SxS���$���b��n�;�\#�x�c�n2��� �Iw:�tﰓ�K߁=[�!�И��;�K���
�����5��#��T�7Vo�-"���:�3������5vtY���5c�l��>�;A�2Φ��[�uK&5J���񍡪���+�l���nP�Gmd�dm&X��+�W��*/��m�Z��F�8�?ޗ���yK�7R��m=o冃��:�N�0��r�צ0{wd|3i�p�D�_QPH�7-=�{X�G^�=�n�����H�� �/����	�'x�ppT#2�L�Nw��/����k�AK|C����ɏ��H�D04�8|0Ϋ�;��0d8�Ɠ�N�ƚ�T+R�	U�,<$��������_���OF1��!��,G4sY�/j.��C��g�5��q����>O���k����V�y�Ҽ>|CR�?R���C
����4>�y�̆�Q)�Zq�&STH?*�"�]ABd̢U:cz[�&2V��X.�z��<z�^�#��9ՃX���'���uõ���4�B9g4��L��';h\~/ �FU|��WI�2�jmO���,U��rXN�r���i��J����@����������E�zw"Z����#[�ߩ`���
���rm������}�L�*��4^͡�6�12O�N#e� ��t�	[�eȬ�#lĻ@�>�{FN��U�lC>^���QS�:F:ΊG�3��D`�J>I�s����5�Q������݁��)�cu7��Y�\Ë���@+F}}T%�B�DͯL��>a{����=���"My6�����Rk�
/��܀�+j��Rc�����P�����j/�D;8��u�2�@��/�ʫ�mXB�^��1O:<�<�Mػ��D� ���җ�@];NpD��w�9W�"C�JF|��Dn���w���TH��2p���*B�	c��/q����@۽��s���^k�	h�NB�E�e�qo_�5	E�,��iD�%,�$yΕ�iʥ#g,X��'�Y5��Sl�8STkm�(�d�}z�T�,[��m��?��h��Ƭl�;9H.Y���<��Gw[<G�:u�������xFY��H����Q�<W��:���9"ݎ��x��,�����fo|�h��-փ��'$j��)�5.Ȩ$T@I#qrq�6��WC�pꆐ���һQ��r���v�+�\^_�&�����BóZ��^eF}��B��WLn��AGw��l���K�9K����&�v��c\63:J���3Nu��ܧJ��4��7��(�k�� �<��~���B�ZK�Ȯ�B!Ţ8 �24R�}u�y�zN8�~d�G��nk	og�\�#X�F����թ����� �,��!�8�5��k�B�`f�������tƥ���=�{��z��]�>���پ8G�0��N�.�-����i,�%��% ���m?�p�*�+���Ky9�$B�*���[���c�V����ҡV�X�U�ϙ;���3��3��Ϻ4���,d�%�q{�GňICi��Y4o�!�5��Jo��������2��&��AD^
��1��]
�Υ1b\�C�g���Q�3~� E�K5���B�SKNm�Ǻ�*��,X~�lm�q����)�g����`�$���T�ӷ9�����4H�ݰ\!��?@�C֙א�[{`�%�px��n'��lf�?�g���i�Y��J�&ԣ�����\������"~C����&.Eo��Qi�:��z{����.��wLG+3�9P��@yo��aip�[���D5�l�w,Ӏ&*�p4�w`��.4i�3�Q�뽗��F
S�c�̦��0��c�+*���L4"��"�`ɧ��D2%=<ؖ
]��c[!д��n�b����Ȁ{��41`�C5���ǰ�xϔ��L���p�EC|HĜ�5�i�����.䫷�S�4�a��s�qT��W 2"F���G����s��0}���O~�Ƨ������1(Z.�,��p�B�ˡEZ�OZ��K��_��������8ϓL��[!���'�k^(����v�V�5�͢���q��A����T����E��PL`���j��G�
?���Q�$cp��^�+�Q]�Wh �@��0�h�EΞ͖����6p������H���A�گ%�J�'l����/>�,�8ģnL�}�è
sU�6x�\5]؟e��&J��> 7E�-�ntI��8�7����5%�]���	a�K�׵���j	���i�}|�iU��K[��U�S�R���hG�/�}*|*X¬K��? ;oj9�2��()�;g(��&/���D�V?<-6F�a��ɾ%g�a�p&x�f�mC�Ur�:I�,�*��߅h#�)�]x�|������G�����Pi��N�ʦ��첂�>7�xꐍ`����;M�ڸY0�q�Űs���i�ܠC�k;`�{@�2��6�)	�����������q&��V#om�\�r�R�ZQ��13h��K�����e��v���Q�}R���	���<f�/B�Rd{"PR�%�w�xg�3ڧ�c��F��&�LEz��q��C7��;�]�3�����WjY���R���kd�j8��~(�}=�p�8�����C1�|"�Ȳ�r?����w������ߥ�qޛы�>�'�zc�+[���L�!^��#�����=�h�Ato�Yv|�j�A�O��)A�4����F�uǤ��zGv�����;Ր��ІrI���?��	o��$�5��H�������^ljt���[R�o~���pD[@�lKh�L/�jX�MC	ěy��k�E�p��-Sh;��"���+���DFh#{l>��i@]�uvƺQ�xI|�(#��C$W�mK���><�_����럂��g�wB���[�'z�F�l�"��K�h−�O�:��e ���롏����r��j|�p�2$�z ��\��Oa�}���C��\�]}�^{7�8d�,YW����#<|����E9�*C��lm}�V�9�+2p�Ĺ�lv�\��M��K�W�����
�2N�s@B� xSgY���������XW����=[�7㭖�s��!|sW��Z�%���Wn)�ҏþ�&ܦ��&��!�{�5)Ґc���/�א&���lY�|���Mp՗�C#a�<~�j��RMA�~t@ɸ父)��4L�T2�YD�ȏ�U�rX�Si�B�KW����{ř����0�3����z�|0�b��ῆ�i�j��t��U��G�����w�Q~�St���>qU��]�Y@�*�]l?���Y���#�J6����*�ɖcҤiW�~t�s$�5�+O(��kT8�D������F���}�FŲ����D9jT�\��{��Xf��a��|,I�x���Ͽ>m3�Ir1\��S2}�;��%J�
�᫖�'�()�����rcɯ��%� ,U[�-c�C��3����GQ�#�I�y�*��l�h��tR�4������U��������ls�3g�e�e��y�G����~Rݠ���^�H'K���Ȯ��uBejT��8D�/�dr��6�asC�DQ�ճجZ���K���Ei�8�{��Go����{O¢�ZE�KӢ{ef�/��mg4�>dy}Gf���B�wqHG7�OF�zK0_@T�mYR�tꨭc����c|?�oH�mp���<{��N����n���+�F�'S��;�cl���oaU/��Q���7"���y�KKU�.��?�WMa��7�7 Л\XW�,���W�}CP�O�����\���*3歩�@"�<����APK�P�w�sU��-ƚ'���ʸi`�P�T��>�SQ:%q��h6-�Uf}��V�XUM	Y�=�-�i_�=��<R��U���y�p�}���e�d�=d�N#�J͘����`θ(')� �K�!T��qs�^.؈})�����.�5ߋfk
�nn*�f�a��YvKDp�e/�H-����n��[�t�V湌V,*�J90��8�?�Z��9&:�¨�M�o}��Jf��}{��|m����1�\5۪��ރ�m��Y��D"%`u`o4���F�w6a����P:���68��c�� �F���rgF4�s�=9��e����=���]v�꜕�p^FB"�������Q)��%L	�eQ��e���Wyl��hL]�f���JO4���2�`|��ᅅDэ(Z�d9=������?a���OK���R�.I���F��Aǟ_���E�]Y|an�b�~┩=ݾ�������ؠ�>��I�C &���� �_��\9.��eI���D��Nݟf����v�`m<��`N�ޅ�5"6s,��Ȼa<V�F"A <�Cyο}E�ۂ�\�u������Ԛ����zW�� Rn�4Y�XC���(Η9HN��?|�{� OI��ds`�����l�V�[��^Xly|������4-r���h��Yz�2�w�3<��0ܑ��ūk���h���C�mC�҂\b�Tna�i�r>�^%�e�F.�-�I\R�B��#�Y��L�)s5ԪI
�}���<����3K����8��dA5/Rd���0���|��[s�[à�����z��b�I�j�.�����lͿ<��~�O�tՑ+&>8�"��%���Q��?�D�\Li�h����Y-]�>��?��Wl��Z7:>JW?�&�VԘkd<�-�f]�K�T�>��Q�z֕т"���x�}n��(KOx�C}�8��@�cr� �"���IU|4���wVɖz	!^/�¹���;�r�j+a�E�l�N��jõ�?*��z������%d+9z��19�d�W��$�q��U��s���p�U�9�ԗl�"��6:���ײ���D G�M�$�!���I׆|�+��m�ݵ"�
������"�U��ai�N�c�r�77|��X���h��Uw�&u���Uy̑��#S��q�� /=R���Rf���
�=�"�%@�	t\�@_0��C�sNd��4б=Bؗ8���٪i���r9=X��Ș3�4��iK$3�n4����h4�P����ę�ݻ]D�7r�E��i|��[�7&�޵c�v�������<ƈ�=�U-��{Mz��Lw�$�l�*-�8�n���$x*jXk�w���
̹���y��,�3R\�g�`�]��  4N�Q�2h�C}�)gL
C��6ߣ�N_��7@ֲufe�)���(����s�h�	��XS���j&U�S/U;������ˉ�X�OPU���|}zEbH�"��kl�����o���)ێ�$�0�_B���_{���i1�d?7���q����<� &�-9�!�Ի>|QN�Z �9ƅ"�\t����Wt��_\�h�A��/W~: ���"��Ώ�{c� V(�*w��2C<�2P��! ��6i���ӺMd�=�fJ���7{��$[0!���օd�M�8��#CMÙ��N4�q�=�G�/
��D���-ijQ�2�����$ɓ�u��E��oz��Z�ןy\��w�E�ĝ���
Twr(<t�� ��s�E%a�NB3����ٟ@�3��l�:�U�9��(��Ï�j�(�H�A��,@ɐ��Q��	)�ktv���H�V��Hx���4��3?��e�/t�.�p�����ifp�鰾*q�W�H���(�������ak�iV0a)���+PQ���S��ɐ��؝�:�dEt�kˍ����m��8<U򠿝�J״b���.��8`���Hl�[���+w&��`T�ǘ�"�Qxs�1�dٜV8+��~3䕹n�e�?�-Y��I�2s���`�r��jnED�������!��h�{8a��{�)N�x��i=?�e�O��r�U8�B#7��O񻌊����� w��#-�X��@ඎ��t^�`뾖�D�KV�C��zU����A��X�_�~�����+��|=-d�U�ȑ'�H����Lq��b��� �p�&��!��|[��V��R��$�bGv�,U����D�q��$�#��d��y>��&$������,�.���ٯs��su5���+�[��^�mݗ���6�j���
�`������C��ޚ���Ut����}����1�u�x����;�3*Ԃ��	�AR�[�/+�7�C�&�,	c�H���G2Ys�͚v����!��9�p�iK��4/�rT�a�Ŏ�VaG}���W�F=�RѤA� �>���+�hT57&�%1����#;
��c�Wb�3�5��un�q"�(���@���&Q��r���S�䛜ͮ��=1�(ֽ��5�N����SӲ2<cB2�I����e�_�3��8�j�2���t��|�/�.�2�R��Da�iy@�{�b���Q.���Ѣ
�� @���4Ƶ�����¡�a0�G�[�|�5_E,��Ccd�bC}O�75�k%Yř� 3c��S���ԝ��ڬ���H<~������[v`�O��p�O��/�b�v�p��s�������s��3����M����U�t��Q�_ep�-��W1ǻ�;��D߫���(�+8��codͫ�A/n+��?�Mo�aLz��8�&�����R@9��F�)Z�|��>���ۢk�Q\j�ET�^+�2�<��z<���T=t:���5��-�!�����t�n4z2R&~�����qN5A��Ɍ=@�F~��HN�$Ry=��e	�*%�7��!*�3X��3}�!C
�Y�����4�`���St�)�v��L�ݷ�X��O����X�M�^8�Ȗ���I�Ѫ$z�/VEx�O´r�-��p�������� ������ٿ�A/�&�I*g�77%�g"��ܧ��-�Uj��D�5��h"��A>L�(������+y���K�չ�Ʈ6d��:�F)����ɵ�|L��fՁ���|�j�<����d�
�&<�3�˪8{F��D��W�RP5���j�*j��3t�}۠w�4�t��<W�D����q��(�߅Q�.���S�}\,J$V���m}��֝;2r�e�?�������OSYe4��ZV�;|
;*���~����K>��K��j�2s�HT��R�9Z�;�9�!�s�X�m
B�1S�?��&,Ю�����*>����|�����X��j�ˇQ	���*
Gߗh�R������"t"�l�ڔ���>��rs��~�Y�:�������Ր����x��aY>��
�4�]t�b��x.�U`�pX(�f�>�k�q�W3O��[bI=�r~~zo&,{��\8U��v֕E�(�'F,�78�#"�ħ2�\���}�	��E%<L���f���b��$[�6��t�[�ة�r�e�u���?�)"��݀uD�������A~���8�b�J`0��P�C{�ȿ�ؖ݉s��9���MG���dI׭iF������g����ɘ���sV�QY��R wT�x�a�d$�1k�-�{��0V��x�,��B���~� A;�����Į����
��nZjo�w�d.��4i����Ҡ�������4�+]7mQ����ҽB���R��W�A4�ٴ'�I�����}�\��U0�R$�^|m:I��Gs.҈*^�`��w���|aR<u��c#o��\/� *�[�(baIVmg��#�����t�j��A�����ozu��4CA�����&^6��	b4Z�[IvW���Qr��v�2��)�b���F�mO���럊v"�~�P;O��h80t�rn#ی�n8?M*�^;H��u�ҝ��M�g5�μ���Do���Ι��H��%�w��
����״sk+�p�{7�'G6�Z��� ��A��HVd��Fk���h�$��"�^� h��\�"Ó�+#u��>�
��Y<�a�L3�q�*S�v8~�-X�9A!MG+ӵXn��Q0�/?BM� _Q6�ߩ��Q�$C�6s���$&�bLI�aq����HJe���qH��Z+u������]wF��������;�[[�՗%�喊i�	����9�9�7ly`�`�g��jC�,�Q [l��-Vo�:��!G�%�	 ������w�����f���������bAV�;����ס�"S2��=Q�w��/"�Hq�������A���x��A���m�<��0����*��W��H�>CA���kʔ�HWڷ���ڳ�ڪٿ�U�U����
i���2^ ��{�q= al��C���~��݈`�H�SRk��X��2�Ƶ��*{U2� �9�q�V�nÊ%�5���mR�,��DoF/��e �Ĕ!�J`����/RS�_�m�����v��L�X=�O�ʆ#N�h��R:�#>���	�������=����\�m�%L��"@���-.�`]�A�士��-���S��Y�7/8"��*�K��<�����2M��>�u���u�
*�g���F.��υs���5T�<�6T� G�H�Ey4"��ک�E��ھ�F�tBs��ˣۜ���WT�]�X�H�X�4a��qt� �67��qiN�ˇO����bY�A<�"�uF�H.���k�H��m��bq�̚�`R!�~�I���OQ#P5��v��ӏ�&2bv�i4�#;l�;�ʈ-"B8��XQN����2�ls��[�г��[i�l�m��	�q�	���=��:�e���[$�詖�S8��}���'�) �q�eg�[s�ׇ`�g^�V��?"Hj�4��>��Ra<v襒:�������6�e �%-��������p �gݳ
ݽ�P�1l�!�!��m�T�9��k.Yx��c{/((�vϪ2H^��``V��$	b� V(Y�^P�>%E5D^?��,2̰�r���p���Z.�LS�;W�J�IdAw�Μ4^)�����ϋԍ���"q��f��"QIzi���:8�q�75�slڪ���n�A>���{J���X��ӆ��u�)�ؒ7+*�S����Aܭ��j���](��P<r�ǵ%�H�d?��.	��n4�Ɩ~=R�v���d��XU]�A�;<	2��T��Y�����&:��3_R�!r�\w&lL覮�Geêc��:و��i���<JR����l�߳�5�-��.��8I1��[չ������A"�M[�J6XǜiG˕�<\��h�c.TZG�]�V�]��d�	<��xקJk��k�f��	�`&��K� חX%n
��΁����п.,Nn�%Y��"б��?��`_�Q�%�h��ћ�ʪL���b��y&��f<�Y��6D@Y�3��Q�m�k� �+<�u?CxÏvo�l& Wї�a+�MA��C�H�#�P�%*��}��&����c�,_��<�t�E!sP6#I����R�����^.�7��,������ ��	vM��*�����-DѡA�g+�vP��ےwO�"�R�o*�Y
4{ޘX����T=s�׃� ix�F�O�^AH��`~�?Q7��Xi����B$~4��/�^jȅ�ĿT�h(����&��a�ĸ�á��T�D���>�(06�,+M�*�
�_�����0�6&2��ɫ�(�����l_>�x$��gL�:VWt"�)D��ݛd�����S�KLya�x�u�ǜ�<� 0�9/�V�iXxP��F�TXC���1wgb����L�b"E������P�2����h�M�#TK/��q��$���m����]�0�|�����1gs���fG�j(�U_�6تt��<�-��g��8�,Q�<9�n����r���Ǧ9BV�Ӱ�f`:
y/v�Y/�Fw1�T�vg���LE��"l��.Z�K�z�x�L�O�iwWScZ���f�1��$��X ��|����L��P��)h%�=�e���4jP㰌�.3������H4QKowΣ�(H�XY��Uqȕ��X���p����J-wBY��<:�wĐ)�uɯ�
���"����IZ��#���n�ٮ.i����W�Rcm�@ ���GXY�l�tӢ������W�uwJ` ��z��K�GCv|��5����	�GxI�t�>�G���_�)��3P�b��h��E��Y1ֲ͘�߻U��e��Z&D6�����h0���74��<ޕ��2D-�b`_��闹�n��T<��nT&
�^�5�69��e����UД~ֹ��v��r����x�$�( ���~.�j���f;�ʼ$�;$ �xS��~J�㏷�v�ɩ:�e����)�����R��ʪ���B(���M$�����~��/Қ�|]��'�1N���>�2\��?-�B����+���j1����X���WЃ�/���TEZ���T͵[�&_����
��I���]k	Z%��f��0���:AI+	���ƌ��J�.���/~m{v'+1ꩲ*傤�T3�!]9Ύ�!��V����:�O����2��qZFf��J1�[���¨7Ɉ��A�E��̂���9�>�m.���J��o&�vtOr�FlFt�j� ES��k��^6J���w2O���֗ @E�.~��� �җ��'�o�����J��8%C2��:��6��̇1:�
n��~8RDk�#]�����xn+���<MZP,��V��P��d�j�����ns���u� f����g��p��-���8Aݗ_�z����v�e�y��=<P��H�s�����B���@���=��ǀL2�n�3�q]�۷���C�$�Y�x�=��	㹑��|��S�W\��N3��ݞ���$��tи�-�ϼj;��=ӷJ�s�,lCG���Sᔨ�3�����(*�Vu��h������ͪ6�w,,���F -�� �=�nW���(L�`X*?hX~1��hXC��6��	�6ꍢ�7�m�ъ��~����#3D��d�Z�1]���P����pZ�'ʷ�����%!`Tn�:��� �c��:���`j˓�y�=[��?���5۟�T:
_�f�y�>����B���r'�}{o���3��P'��RV3Y�%�qq�����j$�ZE]����եT�'����<O8��wN\�[�HK�#�� ��V��r�^�!��S[:�b0|�_��P�f�K�S�u��r��S���T�����ˤB)&�RƱ!����-���h�'x׬qbb���m���64��
�߭�!G-ӛH*�k�$%��0�a #��C��l?f�����9��u�|�˽2ؗUNܦ�<��ah���{{؜�^���hI����_�f�W���H��袻%����j-��qMi5��y���/!/=ct���Gʈ���T����#�Q\�{��s��<�@I���<Z@X}7�e�֡���p�G�7�8S�eo��Ҋ�~�t�cG��4�ύ�P�aW&�k�&��A�[�������"[<�;�N:hy�?l_m�d2�f���>�w�$ksIe6g[<L��v�I�5�_�[�^���a���J<R��� v��:P23l�����ߒ�6B���t-:��ҭ�2����m�v��T�*�B1轞�e����,�i�Њ*�Df-L�p�ٍK��z���~n���h횜=\D�&�1����y������U2";V�~������Q)������%I�$\8�q�~>�m9����T$7���V�?{&	?�>�x\��ɇ)d�e����h��t��ۭI��7����,�����2�@,��$9�C�q�C�<5�����?+�L�5�)%�۽��i_�.�;&� I�v&�Tb�uT3�L!��I��9�麄��e�/����vC~C0y���@W����A�3�H΋%o7�~����)��PZ�v�N��2�շ�DY��rSl�R�� �/"8o_lm
��Z�Vq#X�a�0$d�ȧ8�!��p�Ѫ=S�7� �����d}RY���mN*���O$k�_�p`P�bv�� s�%KuX�량~P�y�)*��&Te��2L��,�L&�,�w؈�S�i���X2���j��=JB=(�8���`���1�܄�/#:�����׹T�ӻ�9d�z�����#���e$��E�@4��������/=�����֫Zw�$G��ϼ�D��Y �p�7�W�(N@3 ��������7bnr�i{-E�uI��{���'G�D<)�0 �Zf����:��Gؽx�vH����������h�u�>uj�)������l%�\�o��y�����v_E�;r�M����	c����Z�H�sD��&���Ȳn+G_�\z$ Hێ.ɲcܺ�}���U>c�O�4�2΁����rR�Q������6Om���h1���x��J���]+��-��w�ycg��[�����-��=�x��Q�]6��3��]��G��B�ęA���w�&j�Q��4�kq�/���'�0�-�a�pM@�%c�ڪ1�ɬI��"̤�C�,V��,���`�|�����8}���A�ӳ>C�c#6c�,�i�O񿱶F��K�V���t��y�
X�q�}eH���~Ӿ0$|�F%��S��X��J7{���7j��' �-怙�=$9���G��C�DQ��5UwI0�u� �mH]�X����
!��kB�������I�E��ղ�.���:sUS���㑲��~���Ia57usF�@�� ��c���jk��
B�|�4>�-���-�p��vP�I������_UϸɃ/�j�S�S�\aG��&
�:T�.Pȇ�$���T�'Z�b� ReP�q�lP��ݘ�b�A]��
�u(5(Ga�W�%k��:J�f=��ob��í�&]F�Q1۠�8�
��tև�n�ӓlNQH�	����4»��>FR������ݻ�҃;�>�KY��[b�g���2>���a�o�p�S�U�U��y;�0O��Y�!'?mp��O�pM;�0�G����L:�����ir��A���/ѭ�,�+s@�W��Cmq�]M|X��o"�`��Ʋ���Z�e�ק!�a���V�<��������R�0���I�`y�K��4�a�L���=zc@7o&���e�|��
��m�I�#��M���eſs�M�Ky�]��
�Fk^$ש��B��iQq$�G��M��PM�ڳ(u��Q#&���µ�õ+j�N������E**�bHY�y~� C �Ƞ���T����nP\�~	�æU ? $���"������"�CXmoN<��yV�*�iz]���'iz(���2��ԯm�2߻��,�S�g͕e������%��_�Ȕ�h7���TZ��\��ï���}�H�8�Na	�?�9�C
�=o�iA�57�2uE�'�Èk��93��8t��E/�
���r��,]4�EYxt N�p;@�)��Ӏa�������{����$���
��5����	̤�s���g$��	�nw'�ƖL�KZ[X���סؗ�J��f{����,e�CG��bs��.u���VS�2��#6{G��r�<s��%[
����]$S�X'�T���oZ�r{M��yr(�P��w"M�/���?uq#X4xP�r3��#��YG����|ڛ���j��nvm+�w�=6��Z�*�d3C�EJ�5��:�%;!��;>�?��O���Z`�Zۉx ړ��މ(!��6Y���X9	����m�����0�� ���$N���\V�BB ���\�zŕ&ڏ��9G)/2��3}��Ve@�lR�.c�S��E���;����c�F=��չ5�����X��hȁĳ���J���ʞ��A?v9��܄<���^�ZV���=~�h��>��?��c�l���s=�\�Kr��
8���q�L$�2�����J@;���<�gϞ��l�h{�Uz9�vA��X�VZT�t'�7w�7;wH]�n�Sd�t<,�O� �w̪�����cuڜ���@sQ��;I'q��`��9v�֊���x�u��h���x\�`��` ��\y���(#��:�f�I'v�ΐ�"��L���3��q��>�Zw��d�Ģv��g��|%������"�}��Zw$���[Lh�^���x��b�s�MT�*�lh�#�YC31ElH۠=����6|6��i��X���x�T(),R������Q��ϘLxI�&�����&�5�Y�'�d�W�q,J����:�,�pנ�6?�n����.���'�p :]w�/l���p����|����\��p$[��VIC��X�,R�S7Dz�0G�ra
R�0�\��Fc<�4�p)D<��:.��(#�j�Tۖ��_0��U�S�?9~߰��R�ܑ_W!y�+B;�=G�1�����s v�҅���S;�昲�����+̤� �@��v���o�bX�6,{V-�y1��Pn����b� �-�Ӥ�h��[j[��ۡ���6)�N/�tY�c��H����5�}%�/��ٛ��Nq)r�N���G8�"�3?Q/�*��KX�{,ό� ��)�^&�Ѧ�XR����aoy�d����u��Wh�l�����~�QřZ���I������<ƼK(�ҝ��y�0�N��P$OMwv9b�*�$
������?�4��%��X�ekG�<%��96�}�)�* �'��i=Q���
���� �k}^�p@���P�S�$���ʁ�Mty�ժE��%� �#�o��U����\��������4{��"u��ƁI�^�2P���j��V5 ���E��׍.V�/�`��ݲ� hv�����)����69����੏l�@e݂��^�`���&�0�͇��_[1��3�p���|��໳:1b5M�@��������Oi5�Su�r�$�����pz�l���E�y����T�	7�&�8���~��Z�
s�q�UY��̓���	�w2��|�^�����޴���nQm�$>˭�������5�C�!�Ў'�R<l��a�t�4�c�.�~Zbm�K����~��I���m�H��8�zb�}���)YU��#|�	Z�dϪ��!�:|�}`}o���+���(Y	
�O�B����Jt��j��On�
!�m����ľE+�n^(��b�hEAD�3���c���4�GN$l����Pu�o��rt��V��DY5����_ǵ��S�]�	m��K�(]�Ng�N�ș���z�y����K���LT��nm���\����RMi���B�8B�v���Qm�Ƴh�,e!'����>����1�c��SQ,Z����o���-�@�I��ĔƔg���~G�X��L��v���+��̩����.��re�5���U'�Ή��Y�^Z�)�L�������`M�8���H��-��xiC^�ȞX�^��)K�_曇n���GP�����ge�q�`s~����� 4镑ϕX��g]�ę�g�`����P��>�^���{xM=!V�L��-P
��9��b�p6,��I]Y>�{:+4@��w0�a�K�t�(�Df��M�կ��n��䢦�X��V{�,j:�yǨ�A��)��&L��~�5@��/i!i\�l�����Fo�kjeV��܁bՎ�j����P`���_IvV1��*�o'>��-�k��<T7 B���$��j��'M4\�e$�E8HRn�P)+(S&�pG<F����y`5B����=�_�h���g�ÑO�+Xj�@�CE��|�Cc���9�,'��T�*�j$=���mo=�$��o�&_|�6<C0�3���p�`t��Ўel�ƌ��zKH�O����o�T�-V��^<�9����w�^j:,\����ً��ryݕ�Pqj��MP��!��C�[��--x�W@:(�>n{��}����e�����3�u��V�z�D�7Ɖ2Ͽh�$����ҞRj�%0�F�y���úR��>���eO�dC!Y }��ʈbc^Y�	�/:V(�����v!�J��|��了@+���u\�1|��RΊ����*��r������y�6��e��@!��@K,�����,�s�����m���2$�kĝ��Y�+��)����M��3�����J���Lz����u�&FjDg������\�� p��&��82��~j���_�b������[��X��I��6����tHe�4�����W!)c��\Ĕ�'tA ��,�6��B�T�ː�M��Q{����d ��/}>�L��N�B����N�i�[�V򝸵���9�'�Ar���i)���'���W=�ߧ�,�N�4�PD�
ЌR�^Ca�WP0�<UQ��u߈q��$�"&������HR�_�9�&�#��1\������@�X%!�^�@����2��z:SR�UG���ް��Rg��b&�pY�\�R����X�W�;f��������u^�8��������P`�jĢc:I�\ĵ��
�^�K{��)e|~�ɀ��m>}�E  lD��"Ѫ���R�@9���|mC:��tn.�K{��^�}�������B�IV�vy?��E�`+㾘׼�OX�Ct��L=�󏿸�n���%$!�F~�[��!�5j0"�2�'25�x0�Vr�Я��A�\�
�P�%����NK��"��Ͳ�)zW	q�#��g|IH�^%ۯ�#_p�),Z����p��l��:�n�4�_I
7y;���Ω2��M��e�^Nɪ�B^.�]#}2�������?�	�f�������"��v����̯t�<���1D�{�Y��`,Λ��j?��<T�)0�'WV�Td�΋��.i�x^)�u[vCYC�9"uvg:���ݴ�nj�Qj),��{ WD1�`��Y�hhx��?�܅ўس<!�<��>��G�G6f �����<���.��۲��F���8j�o��`�hE���,����~e|TS����M��E��g��Y1|�x�V�xDu�eJM{�IZL�t�ZiFv
[��T�_�3���y���^_���>1�����o$�F��xd��A5����+]Z����XbA�Vp�u�C$`l�W=���0O����2y�?n���atqΙa�����rR{4�.�1��t�.����Q�k� 7�e����;ܯieͤ@�.lHTقЧ��u;��AG�j�e��R���	�im��cf�T���	��D�s�OĬr%�"l9jg͛곴��P��2���\��B���'q��v��:�ys�>$�n��3.?�?Se-$9&���d�Lޡcf�˩����c���c�G|n%�9 e$�[J��˫D��j;; xbj=]Ca�����R'�n"^�y�C�?����R��Ǐ��nr�;2^M��Ŵ���z5��c�*m�(�8]M�b�q��U{����=��c��2�Pv�ڄ7"q]�A�]O�������;���7���#@]��j��r�S���@e��J�S���@�/'Q�m�ucӆp,}��D[HCN��������������2�rB�R�I�#��d%�^O�������w�+.+$�nTA�>�^�a=�$k/�)n%����T�Od5M��&���2@_O���x�:�	w���c�+�Fꐃ��;���.r����ևg�󉈯_52���ؾ���w�yI��%�F�3d�qAW^FK4O�Cp~�,1 �H����x��2�n�nP��M��R>�h%M68���p��~�2{��#��f��.�7��,d��^�����0��
Q���4�/VD̄�<�PY�?���{��~x���k���}��L�� �R;�Dˋ�UPrkݼ��1m=��p�˨����.�Unٲ�k��i�j�"���KKe&8H��Uz�ݍ�2����������b��8s���q`f>��p�}��y�kY4Lj�uA����pgN(I ����Q~��/�3���CxEf1vx�4N�Ku�h�p�&3����T�Thz��X�% D��-�)�y;���vĆ��
����7��EVóSvqR�D^䶅C��{�Cu~s�8������W��hN�Pπ�F�
��L����W��<|E�Zsu<����X�g�5�x���!���6CTQtNG�+7�˻dc,�?4�<���"�~��f�.��7��Ćp~O����� �����j )�:�d��76� ���"4��`Ӳ�M��'N�0��F�V��fSh�и��w���-�A�u�ӭӥI���ׂ���l�m4�B��ո�^��^����Æ<<nP#vA��X�v�ph:_N�u`'u�	$��4����0��aR?�=%p)�/�$y�S|/畫}_�>�����ņ���S�KE��)�KPc�Wn���E�ʝ��l��١l̗j*awC5��Q����y�U.l,\\�������bu����V�5"t8�;��-AUz��T�"IA�C�����,��%]sY�}��u	93^o��4��U��?��1�����k>��G�U�Ɏ�.egߚj�I��)\�#�L?j�D|z�y��������Tu�������o"P�܃��9�{�T�/"���u��a���L�g`¹Ռ�n�ʤd�f�����},��GtO̢f��-�E�'���UhR�c ӨQ󞸔���SEZ��n��g�-�k�R�|��o�ٓH>����c�}  	�w!a�7F�n��^�`m����jܞ����QY�c���H��-u��EH��rQ�k�99#.��S�8���IM��2Z�haZ��Րc���nO�\?�!�&�,JP�{��=4��iݍ���1�^Ci�3B|��� ���+�s�}�`�o���)�r=Jb��S�8�����*��Pw�u��V�7���%kZ �x�O�)a��+�>����<���0�#��$���A������nن}�{��%�:áf�����s��8Om��An*��ɓJZ��|�|x�G_-���
%{��:Lx��&�a��V�
�g%B�\H{��$�v+��U�L��R�|�FC�?>?#�H�s����f�> CŋI<>�*f��'o�vu-�q� )Φ�>��1Ⓡ�A� �2z�!�3h@�WS_�XYgd��Y�(�D���V�0�]�J��v���e5���	jx�e�`[Y!]��7�1�o3�����j�� ��������5��ͥ*p!���G~�U��&�,��J
�ǁg�85%�����\|?I0�(�hF�C&���N
`��4ʨY��#��3��r�q.��U��dY��}�?j�Д3`��*>�\��[d�0Ʊ�- �#O'{�����1j>2��� P���#g�+�ac���!�&�w9�U��9����O��*lH*��plX��Y�����0���������݃���P��Z�>��Ws�B��3 U��/'�j�B�V��kWg�lh�w'?�yO��F��cD�hj�/M�����^���ޟ�E}Sh���.)���s��G%�(/�Җwgl�Ba|t�(��Az��&ٔ-O0&�:���E��o�U�v앳�e�œ��^;.��)�b�{3�b�.�*���Q�J�
v�
��B�eS���y�̓�jsЗe����}�@�̷�����L��l��hu�Ō�y��w)-�T���[T�g��,Cʪ��=n�Ԉ��m����!��~^#I�u���vx�&�ľ�;G�7/e7�5Cr��?�8 [q�h��~�#������q"�oG@x*�����ks$-(t'Q�C2��Hq�y���碼�l���t�!qj���&k�*R�� kD9
(˶���I�1�yZn����Kڭҙw]%L@?��)`^i�(L���^@Y�޴�"ӄ^D�1\��;+��j$�/jO0h��u�#������x8:��e��h@'�?o;g�K^@�� �K�p\����J�ܿ�\���h�u�p"���|7'�#��W���>�×Xf8�kwD�M`uq��OǪH����b�c���q�;X�ݍ�,4��"Ξ�w �t�HӨGM�n[ߢ)1T&~;��ki,�����3�i���&qX\bü��86roy���v�K��H f�� �\Ժ���IFk+���:{
�	3oh��bӯ��%z���2�%�H6w}f�M�a��k�CKk;L��������`��J	�����1�f���@Yɢ�0�o��
��{�֝B�1o��/�c�����u�֛[�ޘ��.�Z��_��o���4�0�&=Ϟ��@ʉjo �������v��g��aA�u.��Et�:�tr@O*w���\B�
����ۿ�{��M����+*?�}AÉ�.Wt��qÁ�?sphĐz�z1���Ev(i<��g�ǜ\��dzDF,����Syy��5�R�K���jl���C�wk.Tc[;����F��zeI`w�q��|��ڨ����KћaR�FO�c�!�i�6��%���@���3�Mn�"����8F�T٪׻�ۢ}H��.c���ݎ����	�,��TS%Y~�P���R2Ȁ>��]��Ӧ3
,.�)3���狌��M>K��`�h&�E��m���%6�8BSOD��%��4�h�H��뽺�<���tlq�q�S��l�P{�S��Ž�t[6O�B��쉠x���eCwt����˔F(��jM�C���n��������`��Pij��o*B�M���X��rvE�	S�l]��Um16�VZc#ԨՑ��o�mD̚"���v�?phL�Z�EN/>��Ӯ�fQ܌3Q�wU�~�I���v�O�A��Δ뎬=ʄZ�?�I'
��Tn���C����ׄy�/M���3=i]7�{�el�������E�Kf5$����t�]#�a�r��S���p4	��.��:�%�k�r��H�)����f R� m���D�:�-�d؋�>lR ���]X�{��W5
ϖ��U��F��TY��ε�{q�g��x�@�:%|+i���/
� �;&Vc�R��̯Q
��Wb5����|Y��p�\q������'��s<{�^���O�4\E�-��p&N�H;d���f)�VA�Dܵb������'���x��+c�����Wٵ��"ނGc�8�~\P�,<���P1C��%���B0�e�zԷ���a%!R~Ԇ�M s�t(����� �J��V�0Y�-d����j�C�cu�v��e��3ߥ�F�n=��(�ꉹM���;��Y���6R
��>
U5��K�e��9�?�S����,`om�o0��-<�˞�|i�YXV�r��ܟ�� ِ����մ �)%h}��e!���V���Ȣ�$�nfئ�u8.�O�*����D-�����YM����>M	��-����Hע����OL�"�+�����{��o�(�m_%�/7b-�̈́�q�J��[���Z���鯐=���@4�6�=���E1��[���]i�)�wH�Wf�v������8�+�2��T�u����ѫ�i��\B\��8sox��o�,Is"e�r�V��Q����}��>��c��~p9C���u �);2��<�]3��ڥ�l��S�y3����z��ΪSV����[�i��!#����a����N����H�����\n�"�Ǌ�
4y���0eŞL$(�����0Ie�Y���������~�g��CXK��fm��r�>.H�r�Kŀ|ı%�� �?����o�������s&Ī.�֤�Õ��_�� ���{�z��y�֘��3�^�n��Y}�3V|������s}&���Q#2��$_N.R�;'����W%��M�/��A��q�+�8�$t2����d�T��R���-@^����V^��1M��?UK�D���6!�e@>���}'6j�wQ�[��Ƚ��I��FO���7�U�4���ꪄ������pvX����6���g��������8�k>RȊ�Es،�Ɍ�F����SK���F�&���\��&�U桋�������9Q !�?C�����ޒ��U%=��
��~�c��S�k����ލr���&� 73�-��G�	��4�Q�[�0#E������<\)R
���PR	T���r��+��>h#�B�ɫ0H��㵹t��*��P�ǞĖ>0�L%~����Y�-?Z��ng��oJ�v�R���X�*��&�{j�ýU���eݤƿ-GC�ˌ���$+e ��8{#�p�fI;gD� L�(��Y���6�t�G�ktg�/w�q�E��}αT�ڷ�_�~r�#e�
$�!�0(�Z�fJQ�.s��ɷ��4������)	��,�~l�ko"Enf_�+h�m�w�d�iĎ���GV5c��oƠ��8i,�S�����KH�j�b%߈�wéV@a��o��95p��^.oZ�^mgΨ��:�(�Kr�xn�D�|��QnJ(�(�_+#�ٕѕ\G�h��#�:��g���_rU���rP(��ۭ�Z�ܒeY�"�<%��y������4��膥�[�$�RwY$-�)�i/,���>6OՕ%��d�4r�`�R�{�{����!�#'/�S�f֮Ʀ��o��7c��mo&��N�D�B#��p�9]غ փ�?I߰O�La0~�gC�o<�D�&8`0:DS�����b[1����mp,�7uں8�J��@��������KT 7���!�,���^�"�a��EO���|�Q�n��vjI�Xd���}e�vg���������~QQ�����r��1~=H�[B~��C��8��2Or�;�����=��"m��ٽ�I�5WRL}9���������[�ǵ��@gi�^�ޓn���/�Mhjr��i��E���V̉k�`B�WA|@���6T��z�2��	�j�	
;wu�:*�e�m#�xD��rK�2r��_+#�Dgg��F#L"rLm�?�v�x�	����&�09d/S�d��+�_OHS���9�9��ZX�)6��?��3�B�����aIe��8�X7)�GH�����<��)���ĦN��	�Ѕ�i��j�s�� ���Ҭ~a�.$>׊�wl���l�?ٸ:Z���ս���$d��˖]�����	�br�i̢u�h%ڑقf��t���M�.5ZF��T�P���}u
w	����5m���4o�G{�u�/��]�t��zh�R��ُL违*/��z������r�T��鱁�:m�ה��Ǻo{�o�sq�����n���DE	�<��	[G��I����mhld�ñO�R���z9xN���V�M:���)Ӟ9s`;.�і-@1a�,8k�ܣL/�R?=48���+3T3b������[ 6R��S����\�<e�ߑݼA�����QO5U�L���b K`�є�BT��,�`�!Z��8"z�>O(P]��+�XsW7�0L������8��o$(� $�T�_&$�ulHP|���rW������z	w��3�����H�Ň���� �	�	�nmϾ?�#�N��]����ĊJ���ǃ�T��Kkn���jP�)� �JR�J�uw_�������xɀV�{x͂:����2�uО@^���m~��}��0���@�TU0�_T���m��y�&�u��A�J�_����Q.
]��?z�x�7M�N�"t"(BqO�To�����ϳ�A��a�������!7q2�㠽�w�g�|��Y�]ކߍ%�5�4���԰� �&����{b��^�
/7WG�Oƿ�[�9Ӗ[��Dˋ���O��7�LBO�����S�t�@�P��V\s�P�&���mG]��}K?>�TO����L60���0t����d��'#�E5��_>:ؐ�����; �(r=��JV���[)�4�T�v�I=l$����4�GJ��z1ݚ&z�GȰ�#� TI����Q��e��Ҩ��D�+(0V1:� �p�}u��jL���j�
�/��Hp����;n�O�Oh���?�[�ݥ�NvV�}�乐�L�3�8L:����>�F�EET t����>�D�����eN6��b��>��)_b�Đ����r����sg��w(�ߝ,�q���Z}�h��,�6�d�OS��D����*F6.�;;A@2ts�tN���i+�+�jH*jQ}�Vބ�p��֠� �~�\���: #O���q��np��~f�i�ޚ��z�1�YW/*hN4+�8a7u�41ji-�l�|�:nTniM� С�V�:��
�@79�1z�:��#&6|��'�*�	x��d3;[��>@c�q��PH{P7]5
�^�'����3u	ơ��6�׍�_t�A��O�7�s�!?���j���}z��.�l�"/S{٥"�v�E�TٟE��X7���jLQx�)y�q1d+d�:gH.��Ĺ_�W��\�1�i5⌑�	)2*�s�1�*;[��n���p�0d��m��$YF3���jQ��$�(��Z�(��1��UO��"�%Q�L#f�D�<T��eL����:���R{hS������\�Wj�RS��V�\"�r@A�u�x�n��g��Kh��e�w����h�m�Аt�iL���6�X�/���ɿ�̖h���C��@f��]�3�:��muܞ�h���V�7��;�J�do�S�3�16�����#;ab������7B���u��_�����Ez��x���0��e�j�a�>Z��5k�ra� �oݠ�Z�M1U�0�w�2� H�
+�˾��xَM�Ne`�f/\�%��\Use��Tz\M�4��
0��R�T�7�-�I�����?6�X��|SY��OȠ����(��mS�Ρ�'X���#�&̀�m��{�p�ܘ��5����`d�פr,y� o��G���>��X�:�+�E���'�`�	�|_�VyAj�C�b�.+���s)/��lp�資 8L��%��@RjH������=��	���%S���h�b,��?d̔��lC�?Cp� u�0! ���� l�A7���~"?�'A�_��Eq�$Ad�0�C�������t|��C",%��Ԕ^P�2�lWT���(<�S��n�I�
F�d�3z��WB�a�!elτ�M���]�v�%������՗�}l�<yk�r
 p2��K��kѭs����ƹ0�<�b2c9�W��)*�S�d��/X~��l�E2R� wf][ӊ/�J��(��@�v��g;�����s�Bf5�3$/�͕:�����C�+�¡;�ٯ+i��Q�2�m/Y7��C�0����>�T�|V�.�\�l�u`P�3�lP�Y�
p�15rPtq{��CiBFv\S�3߻�=�Am|U'=�e;��y7[�������2T��j7rd!4��r��D-�T�x�憟P�-�ϥG��q�.�'�R�G>�;:�q-2�����g�x^9w ����$�ɺkL:��`�-E�W�vE���e��A�ຩQ��&�လ�N����ŭ걜n��d ���K��ּ?���`�qJ�<U�_-}��>q���w^���{�5Zg�
!`��C�a��(��#\Å�D�r�LH�����4\�$h�bk4nr���&��Js���§��i�����d���	lc��#��D�<#�iE�\Z�h��Kj���58º��5�B+7�=C�'Wcp�� .�l��Ծy��q��F�R�v=���H�l��C��K#*oO�a��+�4�%�_��Ny���"u�X*j�I�������T{�'xR�Ī�l����/�י���a���^��,6F�hǥ�P�����ƙ�-F��c�E�>�������tv4���ں�]k�éE>=��h .	3��S�mF�GMA���ȞJ�m ��H��Q���4�Ѩ���^��/|I��
�N���AyZS�ڞq�f���/&LZ9r �i�p����Tm�s�uCES�S����I�E�:c���'%O��y����%.)�Z�VU8k3���D��qӞP���0�����T��T��eS�A>��t9(�'�h�	�V^8�.ȟL%�<��f���7e�Ƕ�@��q��"�,�z����.�q�L ��N(��+P���ST�۝�hŲ{)w�$n�䟵�j{�rŲ��Τ��JE��#Q|cn��1��˿�������%��DT_�X�Fxj�_�=�Y�� ��C�>x���2�_:�T����������syuBB��V�=���t��w��d�9��r*����%��b��2r���*�����`�B����E��T�>�N}n��a�3j��/|S��a�5�`U�SI$>��З�/������/D��ڸV�����Q��@�%-!5�lX�'�Sl�/ 4k��|るK}�C"�!?�4�d��A�Z�c�SF�y�A�(#tF���]��;��[S�ߓ����[q�+��tf5y+��h. iƂf߱y���%��X�QHw��tv�15�zU��WM�t��s�y�w?�B�i��`�Ӂ,�A�Z#�-� Fr���*B�f�T�&��p+:[��!�Y��-���Ql����qp=e�f���^��6^�d^���zc�rSѲ.��q�MOJq�;v)X�+2�5eC�����d0��3�np�]c��FޣE]>�DZ_��oj\~&E���7T�"��E*��C=#�sO?+F�y?�Gm��O�
�����o�+�Y.�K�,�C�v���kX�Ox?��F����`/j6��������J|��^�g�p5yN�ʨ�i����ND��
ߺH��1��o��jĒi�57�F,P\S�*�*�� ��۰��<������n� ��^è�B���(��"��\y�L�p��fV�}���;p[:t.1�%l*�6{o\���9�/�Ђ^�8+�����y��XQ��.G�2`j��o�0����9�2�B^y!	������8G���7��̪���ԷT��N�"�%�	�#��[a��b�=-}�N���J�@
���Fy2@�0q�Ҵ�m��K?�*��u�m��ӿlB>���$(��)�5!�h~)�$oV����]��P)�m��c.�RA�����4�e`Ə��k�#�@\�?���k�n�i�-Q� eG��O:v�(�.늗����L�(=Wyob=�c��Pt�.���{Z;��|;)��2����YX��S-���h�6�N�@�t��e]�>���
K��V�>�q[�X� �ΚG¬�M²�Z���OR+F�8u��'��gQ�R:;�mpߒٺڶol�!	ȼ���]fA<a`An��e&P�������r��d��a^�14�Y�͝�_&��#�����h�J����1o+�K��|g��)��� �R��0ڠ�H[�8yuXv \j|
�3%7m.hBF��w�ݺo�2�nH�.±�Lc}B753G�� w�ˤP
1�t���%:[Y	
�cq����s.� ����C�{�������9�%�}�J�:卑���5�|˪z`�`JM��Q|۱�?g|�3��Cw~�;s��m�ܹ�!!�>�Sr]^׿��!�`�p���l\�����z"�a~�v��^��ȨDŹ�Qw�^�iة�._��D6Mo�VԪڠ��X��$�5D���h�(�K7��$�@�7�!��8i��H�v��KU��2�4\��h�� ��K�[(5�ƿ�Z^�Hg��c�Kp�K�����E�]f�W	�wᚪ�xXsz
4�.��a���1eK��`�_��@G&�4-z������g�9�6��~�U�_n*0Y?���v�����T�`�]K�i^�|�bȃ=\-կ#Xa�I�g1��)V�5���.�߰/��x,iX;Pi���1Q���u�7>=0��2V��IaTs?�����q��
� xz�m���	�����[PG̹i�m�0<�1�ZU���Ha,�EЫ�YɚPrfT��OvU:����IB�$r%L��oE�iP.28y·@1Zi�]�-���z�3|#�L��&��&!K�� ���9�{�|8,|�q&H
�K�<��?QH$}xʈ�e�^�5A4;(��x�2("���߫dB�v<���E�j�Y���T{�,��,�+��)�������`bL�̤"f����F�^�'��d:���=E���+qk�.?��Z���x��=���a׶���1�9{�&�"�G�q�>!�6��4�l��J�B�:̮�٩Mo��U���k�f`_ I7��n,�!�}lh�g2��Ǿ���H=4���j��7���MqW25���np�
��2�QfS~8���!&��`lv^|	6�!>1r;���� 5��P�r�(
%��[�No P�j�yn��sf45)k[�_��" �?���E�_���X6�,�鹱c�����?)�"�k��h�W���͡x�KC
6�RUm���[k�Q�-۴�Z{����]����B���gYap��e���P��!�������ܕN�D8ZT�g�@��l��D_�qH�*��_1�����⢂���X�= ���!|�>���9Aż���1RL���@���d�Ϝ
�Ƃ��6.=g���8��ST7��s��=�3�;�å-�EvS�Hv�ѧUkϥ��<�
�q
�K�$/��P�a*�g�H�eRV�ܲ��X:'@i܀�p�8N��x^;y����:5ʿ�;D���݀~W���Jˑg�yP�j8&!,~���Q��� � �2����OF<#VCaD�����L�e9E�?�I۵�_�����/=����ဇ1��骻7�LC&n�9��(�8��E��P�����6ՀKY����w��2rط�li6���d�"^`����m�0���A��`�$���Y�ώ�?X�Nu��6�K�jw5?��}�!#�;4]�1Z!�X��x7W`+��Yd}r�����˿O8O6L�ړ<= TZA�mH��>�Ә�2�,�,�//'�K
, ߕ&X��*>��/R���p*�]C���%�� +��j�O�����D+��iKlN>I�ED����_N�P�׊?��X�ֱ� �%�إ���9���L�d��)v�ZNv���˗&΍�{2���ۈ�E>7��ߴԷ�~��n��~GM~���!H�Bi�Bc�o�Xy�yfY"��ry��C�ୠ���%�VN�����g����;���bw�
�	V����g����η��B��%o�`�I���FՉ@�����|}�g��*���"Q/�	���> i���*�' ���"g���i.x# +X{���͸��ɳů_��S'�m�` *n��]��i2<?f�_�P�2_ʞf������^$9h�����T�pʃ�g	ٱsl&��T�-9��4o)!�ʇ��v�lXV�g��������
_���"Ԇ|m�ݑe��@�/�g�=l�3� �P5^�=I��L��ѳi��-�=M).*�S���Q�7�D��c~	��[/ȏ�j��`c�/�<K��8Vb�)}��R�a��¤�3������>�æZ]�'w�l����-���#A�,MZi��b�*�~�L��S)ÈNA1�M%C�v�H��� F��g�l��K40>���͈���L����M�R�,i��kf*��5
�R"�b6��#��$�9+�Di; �6���s2��܋�:���"1�j|�`�,�Fd�[4^k��h�޼!8�HGgb�ye��.ȸN(ߡ֘in�C���oe�˲�e�ZR�Ͽ����t d�F�R.P9�<��Qr�$�^TJ(�qqG2|�P��Cv�`�1��	�Č�&���w%��쵮u��\�$�l���ҁD�O�k��:Og��/�}	b�]�����s��vu�'����鼋$�$� �,�1�npȨ�Pb�I|[~ٳ����͔�#t�/�<�&�̐EW��]"����!\��1������b�ާ�Ȓ��A�vt8͊�x��t�� �d��c���OwâOX���� ^��"�����ă�ƪp�w,���N��vFrnN7���2� S���u#ms���jH�{�����.)������2B$#��n\��OU�q~N5��c#�-D+x�2H�X��<k:s��w"A�h�$�C�Y1?�a�G~�,���0Gҹ�{��3$ϓ	�W	H;T�
��"� �=�;����u.p��uE	�4b�w�oj�Ya�ȉE�V7p��ܟ#!JÀ��;4N�E�YdZ��ήo�4�Psh4��_ےyX�.�� ��Sa�c�+�$�4j�y"�H�j4��U蓔:{=�!���.�ܻ��ܥ�}��j�̍W�r�j�V�蒜b� ������@��u�9M{3��"��H��Q-z��_*�ii� ��W�Imu'#�6�V,�)����,:�����i���`W����N1X&ջ���=�d�5��++���v�3����F!^�
O�=��>=����6 ,iT܎C�TN�Mj����ڵ��xZ�8 (�S[�(�ue����z�˓v��Oh�n�����Ro��JA^DkXقzw�V�d�ݫ�K�\�~��p� W���հ)��v�y�h��N�ӡY�<�j4��ɦ�Ԍ	��ᶎ�o=QQ���n����M�(�Q�܅8��M�$���|��<��>>�O�$�?+��@�X���Y=��Eڪ&������[��HP��� 3¿)H�~�Ē�1�RF�Ϭd�-|�Zʨ��]�d)G�8N�t:��|����XW�6�b'�#���`tؘ%w�_uOP��P+���Hl��*܃�`�"��<e>_t�g�C�Ak>'{�&r��,��݉�r���������"��ᄣ���Z'�qO���w-R�� c"�c�P�h����|�������aO��Emh��m\5'T8a���}����F��΂���Oz�E>��ف���G�S�#��/vl�	�dur����\�߬����U!<Y��d�I@�;N��y��)K�t�v����7���s�鵕��=�w��������bB?�|�cd�|IJ~H ��B���%��z��MZL\/� �c w@���9����#*�U�je�d��$�@\L>�Ҍ]Z�O	�S���L�R�g7��K�q31�q8n�}5+=���;��n[��8J��q֕��%RF�2�PZ734J�B�������S�=vSfFH���\�U=��@~��0;p��]@L�(���G-���b�xk��y��D�[q8�HqJ��f��
�i�ܰ��b�{��!�\6.���1�����̽���������ߤD�LV%�uA�^���mQs&��ⴡ��k~y���ǖ�qlP�5��F��Ļ`��}�-ZNHN���%$9[��БR�t]�뙩����mZ��w�����Q�e�O�&v�o7T/�����e(�F��D�� MKf� ��yj�*�
���e
н�����f��2"7ɏF�2K|�Iڢo��׏��BREo����&`�:J���ibH� ���<jאm�3$���B`�Ĝ�7��r
e�ܐ]� ��=�F8T�RS=Vhx��>,?t�7�7�,Ԡ:�+������4�~���6n�æC��]�3��M>��߇�{�y$* �I��?wL��HnP��QQ�o�ʶ�_~��%����A<��i���Ώ��"g߿�c�/���:�γĬ�3+"�G��{ \��<�u���u#��A�弳���1�j`������P��+��	���}Zkn�)4x:�4�pg��u�]m�/D�O������b�ʅd�б�ګ	��?er�1��z���b\F LM��Ŏ#@7�o<V�R<s��	 n��p���n.p��M���ܵ���j�h���Τ���M��g�X6&>*�oFS��2���b`'ZK}q�3���؀6��/����	��.��'�5 ��w�5e����vw�2<�nq���>^��FR�A��4�Zϡ�&N\�^�D�2���rh�x�a�a�[��8���w��q���NCf)�O���@��3�Ł扽c�
0��j8�߆����C�y�%������\�����l�el�Q���:��.�2���m� �F�6|Y?�S��¾�]y~���'�����q���uaF��{�h���VD;��I�F:��b1�͟7�i�2��TZ���u�O���q�{����y+��{->���Q��D���x�_3�Q� Aj��µd�[�u�JLtgå]U�f"��'�YX�gw�Y���o�b�W#��ߐ_�ka�R$��V�$;�h���l�2��0ݳ�_�(�����tu^lOOy=�0�Jp�oJM�߱n$r�����t�i�◖ 3K+g��A��X�ni�B�R�Z��S�h�#���)Y�����Q��������eЦ��
޵鲿���I:��g]R����o�����[&^i#;+��
3	�jZ2�r	��W�OP.�J9���h�#�b����=d�Dk��a��D���s_&B��i�wm���H��`du�D�{���v �׀d �0����@�:���#3�t~K�(��t�m
T�8�XP ���c�%yT�,;�(�1͌�(
ީ���{<� H�f3eBc=X(�1I�j��:եd? ��<d%ư2�5�N��D��^�.ՋlR�g��My �=���$�K�������@<!��@�EC�s �:��~�ү�`�G��]�|�]�M�F���7�#��C�}c��fVʾ!�5��ת�,Q��M�������[ީg���ܣ�`� �[�^ѱv�pU�~ѷ1�t�C3%
�;��L7f�� k�� f@�����C:� --��+Le��/�x�*���T<��@p.y�o�?��
��p��毙�,%�~/[(b�����w-p�p�@����M��+��Ƿ�X�z�[�P�
b����C�e�7�9�#8�O�ӂC'�9!"3Ö3/8z����ӟ��|����߾�En��O$s&V-�]j��W;�z���h�UIڛB�m�e�v��p$m�-瘒[E�W�Xd��{��	ۯ<�(��XI�z��3Y �ug�M�{��?a����8��V�"^�?��#)�☑�����lW��}c����%y�E����;̍iwd�rY�6�5��n�̟��Q��L�A��������ٙ:�d���ʌ�{��1�PéHMp��F�c`4ַ>׳ΙEҘB�.������z��(�F|Mti��Un	Q�i�iFG�� ��2��,B�t�nj#���'���񪑠 �|�2I�ȑe�@���j�=���Pg���������j7���f+��e��7�Ɗ@��cMg"�U�qfٺ0���B�+�G�������&dƅ�r�9��:���4n�����
��!0	�t/��#Di���im���)��U��.^Bh[�)Ҍ�؏Y�!�V�P�7o�P���V����i����Ά	��ޑ&��O��Z��(�H-�+�)�ECQ;��4H���#���ᭃ)
���5���j��֠�m������&��G>��9�O���@٧_��0������R���	|kL�7K���oZ��Hm-W���Ђ�y��X�.3�-����:�G�Рʒ11���^9qu�-���D.X+$�sK�&���C�֙A���)�M���\UM(�Ь��^ތ�x�ԗ�0E��د5ł�Q�Iyx�T�;�d���O�M�`�� !�]sT<�F܏�����#E�-}f��cO�����T�S.�TI����>�4#���"x{27�a�'��}���gD���0X>-�~������9���O�
�C��0�:H2M�brX'��,�l\�����=�|>��f�u5���/���n!�L!�=�������c�}�s���mK���̓�eA��AR�n*ZC�����1�قa���&{�j��u�=+#7���D�UW���e%^t�PdFwT�C���",\꼨�|eOQ�ūd���R�ך<4�ʊ���6�+���w͉��>�~n�.%L���b?ȱ�.�ь����K@(��p9���xM}ێ���M�:",�q�^#��V���7V��r�Hk�!�^�L,v���?�%�ښK|�����pxO��lK:5��Uw1)��-
��91,���$z#�p���R;�������h�ʦR�ׇ������:"x����g�� Q��`�x��5=�H:|��u"�p�:,����2n%*��������Uo�0�[OjQ38һ	��4x��j�=0���AMPk1�n$6��e"UHQ��l��d�+�>Ǣ��ٖphF:$R2�}��;6�L�Р&��/��O�V?t�D�S뇜,l��9��N�]-Q��<M�c�����|�<�����kaѾ����0d��}�h1|�qE��%U�<�R�H�S��Дa�T�t�0aڗE�n���u����z�+ ���u^/�D!F��: �G���l���g>a�Y���7f�8��r���
'BHE!�0#�>0b�����M����K��>���G ��t@
��o��;p��+4��������)T+*�c;h�L�9�t4l�EFQ��'�A``
���T��RR$���<閖�֔>f��'+�-|�l�*r�4����C�'T����qW�q��M 9	&*�����u#S�B���r3��~Dw:��)*W��r���o{z[9���tW6�hM���ѿ����w`#vkX���V	H���/�Ũ��br��s�9O����S����˝?�Pm�;zze�����gē冼 �d+D�g��6^杇���B.Ȟ�c�|e��K8�aKW���#A:=�&o��Q��;�N_�ta>�� �����l�p�^�l�h��\�t�ȗ���'����?P灩�lL����Nlί��I�:���0�-����✖-�[�	��Q���]���bM��v��!��8ے�~�+�Ν�UO���"[��p�\�V�����d�b���v���t��b���N�K�8A_&�Y����A(����k�rhw��'���{�/���tk�S���<aG=��I�'L��I�Ec �|��D;�<[an������z	�tb������"C��г ����6����t{�.Χ?Ӿ�~r�O�����7��f�R�tO�q�����T��dK����hl��Y�A�S���Lk,\j22 � ���̸@�9���xn��fC�7��)��������v����9oK;l�|��]�
&�
�[��C3ES�j)�Ǡ����_1h�Pۚ�*@Sʣ�z3��$ٕ�:��U���������q�|�d�zFYp���0J ��G��>n������eq�0'��b_�/.�fT��[�w*�w�n�EcLd�1��N��>m�crP��h�(@��g�����&�����[�]�z�r�ȴ#�-Ԧ]��v7��G���d��\�k�2W���5XH?�I\��"��i�l�0då�t�*oB�/Q��� ���J2��,�2�����3*�>�\�}(��^]�Ó�#@�}ǯM��
z��#..��~lv�K���U~i�a����ٖ�dmi�/X�Å?�	[j�k*�]�4�I��+ֲrN��f䷷J�饑�E)���-
���O��T��� �������Y��p�	��4���(ߴ�xϧphюp��l�����l�0�fۦ"����i��u�t�cʻ2}����s ��Qecos�4 �����a�������x~Y&qx����_��ҁ�g1��`��d��)��u9�`az�G���j��`^]�1�
h��A*h��)~��V�ϙ�}5y��mu��(��Bz��������`y~�ݕ���k������h_:�Ӣ�J�X'2,�&���	���R�o�����P5g�䬰}��(�:&�˻=&*z���g:�� p��u��g��)GS�C~���b�$JV�*�e\���̑�ް��VQ�6����u�ҹ��g��7�:�m��y!�W|v�4�"�qk�d��k�$XpiD���0M6���l�]�K�V34�o΍4���f!ޟ�a`|Wlkؖ -Sٿ��V,Jx8��(y���4�m1�dRőlQ0l���󋾃��B�H!�x=��9��������.���d^e����צ��9�iZ�h���]�)��&?kq��I��L#��Ն��?��
��ג�?�@Ý����^/��G�H�]��������;C�n�0�/����OE�J�&�8V;$�*����$�t�Jh�D��!��U�A�������V�>u��[�������ގ%*W�؁�92��9x��P)��qZCW�����Mp��r�,�����f.
*�*X�Vj�h�/!ܯ�8��1�y�F�����un�V��:n_[z˸Y`����,x�>���m2��L���i�9zs��2�H�H"���]]��<~�X�߲�����}	�5�F銼�Q*�?p}J���׬Gb*��DiO�xQKԛ�et���sY�2hG`.,��엮��X������Y�T�i��(���Mr�k3q�1��R_�x
�:�\#v��������N�M��%8���>��L*�	�	)d����Fln��F�#+���Kɵ;E����R5��,t&�������ҷ�
R�峻{�d�F��gk�or|T�ayUH֚&�FT>\���:\R��`4{�Yh7K-�UAM�N��9��� "ep�JG�������Q�'�a�:��"c�j��6�}Y�τ�&@�ל�M��<8f��i# �B�O��'�*�eM�(6��\��p�6��ʳp;��w� sP�|是�s˓�b��#�¤���r��J\�x�'��[v�H�ȳ��&U�{�-��.a}=�u�r|k�x�����N��8��F]��2�w��ѝ[8>/��ُ*G�����t1Ļ�͢Չ&�=�7�$h��M� ���P�QC��X#�����U)�<���H�o����ܥ5��_,��VM�s၅lH7h觶� ~�Pm��?����9�&������-��l�gZ����[�O�����i�k���"��g==��s0�Oc��y*̓É��{<��,���S���J~b��w�	-��3Y���������ʱ�3ԟz����M�Iv�Xg@�&�!jٶ�#.V �Ng c2��SCҟ`��ZE%&�P;�h0:���ЩnC�M9���!_g��v?(�l�.�92�j�C�f=�v�"]Y\2E���]6�a�/�=�12�6������P~���9|�ƒ����ݠC=>�MP����C��Гx��L۵���|���':�;$Ś��X��G�E]��sɬܫ�8��i~x�m�Ýy~ S��@�KX����L���d�{�&�/�* K#�%s��C����i�ζ�����E_Hc���S��_�zOK_:����r�
�l/��>J;�� 8v �V�^�=>y@1��F#��A0m1��F̸�S'�S>�um���/��K�A]�(�l���)�����v'xD2�S�$�
�_9u�؉e��˔��V�`���}iށxvx�~2s��s	N��ca��'[���;��bh�X�^~��z�L0"wV�z�}��E�b�"�w�\�S�u18��'��/��zsY�?o�ad��C
���hT�
7����#v\��.����mK���w�Z8a���DK��1p�!" �N�*�'�9�8�1�6�_�gD����N΅(�~�0�,ڳ�$T��4�q�[{� �(Z+0C	`@�p=��
p�+�;N�:ýaÊ���6��Ɗ���@��SB^�ڠ������Y��ؼ���E�(�CXqb���>�%��43�d��HN?$��PkVo���|��V��-��hpN�e�4�nI���a�|�P�;i��d�}y��t�IF���/Ey��˲���[�����"�c �����p�Jl��Ć9����T$)uL��W��9�V��X��b�d�oڿ�i5sQ�#x�!����o���|�xx��MB#�F7���.���m	�ա���J�PJ녵0+jT�x`n���0�����{���·�i �&t�~E��]��{��b�T߭V�D b��u���nudk� ��+G|%uW*��'Yh�:*B��U!��U��5�r��!�U>E�lE�����omYH��ոV�O�T$k���T~+�PU�S,#]�xй� @�37e����}��^���m�3>`��Γ�YU6�s{яP�I���l�s��� xh��P����A]��F�]�5�b�!K��_%�O0��܄Gm>��������$x�L�^��B��XI��	kIJ0��c��p�N�R����a��ݯn^����=>,���=d�5��Ҷ������ �6������§B%��c�<]KGK��t��C�G���	��8����Q��5[ǋ�:5���o�yſp�d��\��S���s�9"<�R�5��BΙ{��.�:ݼ��O�j�8�?N����S0�
r���aS�l�
V\�dPs
�Uis|W�/����ɓ�đa����C�ƭo&fA_�L�7��N/��P!0��ԫ`�x��I�܆�Ќ,E����������5`�=[�#������כ9](�Yf&�,̩��p�Ղ�Q�2C3��z��xpoh���
���4yX�E�I3�(խ6�\{u��z��P�^�����E�� D"�M��,��(m���3�Q��f��{�P5��
X{����Dg��5G(�8� ���<DH�Ȋ�XG��R�"=�|1B�A��+��'�����b�������%	X)C�5�_d&��.�,Zp�b-`������C�=��в>\��_#a�o�����ܤ�̇�œ��q�tG����{�(�h��*�Z��e�g���s3�!��	5I[v
��ܗu�Pm�s��Hw�����ア_Y��1@�'�&*J� �Qdwe�c��-�s���=,1���|ui7���&��;��fMff=W]���]�Bmv����E�Q�g��=��-L�E�T�iCL՟���c3�V-��w#��G��A<���M��D9;��yD���^#�y;��M8������d���Izr��o8�\�KL�]͙�L� `�%�jb,O$]{죟�P�^�LI��˻XIV���;=;��Uc��J�Qkn�ʣ���p�M#u%�?s�9��G�����<W�Uo��r�4��?�-:�r��;��թqZ�I�7X��3�1����,��W��[*S;���<%�B�xBpXi���z�<�������3X�i�]�ܒ���.pGU�F��/�g���խS#�]-���w��������E�*ΟX9�'B`w�fA!�HI���U�w��kÇ2��f#��(�-D�V::��V:�p2�+�/�'��E��}NL^�/���y)��Q7�w��������$@^��ꄵE��߾��~y�6`���:�m0I�^�U��6c��Ъ����޾Sd�~��Ȩ��L���EZ53���b��Ȓjjx&�7����I1F�%@o�mb��A��f`A�2)��j�$�����4�曚\�*+�%��U�r'����?�<�檺st2��ґ��SB.X�ER����y��Y)Cy��GKA���@,��+b]|@���v��?j�O֟��տ�P]���4��ܡƊP*F�y���<W,#�x������s����q��z
Cp��T,c�i�C���;��i�x`��l�M��xVeQ��o��֠frB�V�*�M�.��"lG���B�c�L�`��r��J�A�'Օi�"���E��3�e�k!���`����[HX&�`/;�3;�yeb�J�$�ҹ�Kc.�.���/AY�U�����yt��AHjNÙ�=`��y=Cy�v�#oݍ6�5�!dț�����Ԃ��w���<�"�/'(o(mCi�,Wo��#-����>���?g�ּ�������uW���P<! ��!�6!w<V8��?�cD�9"@>�_�^�L���1#���j�����۝.�Jа籔3S�Ն��&RLD�Y�G�A'�������/�0͟7d�K�,%�S?h��-:�2>�֌�Yl���.^�baz \k�W��~�Lڢ�o�}�E�#�Q�Bg!K�y��@Ԩ���RĶU'�Q��ᬉ$��A�oU������g�U-sm;��ZG决��
e�r;�{�ܖh�9Mit�ؑ����ޱf��=2fC3̝c��Tz��fq;�~����Yc�&�r��>�p�e�f'�Wl�9����+�X��)Xȸ�^��/�[�b�
���5���Q��� �[?s�v�?�Z�D��{���H02|�#�a���A�q�:�f����ٯ��1G#(d�O�R��W�0��MTq!���fپƢ?��QJC}�@�Zخ=`�:8�.2n%��翜k�#g�FF͊��S��o�]��Bl�uU�O�,3t�2""�v��焍"�0�.��=�H������{��22֒��l,�,R����zw.�/�CM��%
�3�����{��;������,Gc����İ`'�T"_~��`��S��wК����(���v��͐��d|
4��W�������F�������_���]ՙ�����բ�$&��
C,�A�ce�E:۴JF�=ίGç���U$�h=�����@��;��-����u5�O�!�FrN�[�;+{]|$�u�I<;:��I�Ă���%9 `�8��x+�c�]�����L_>�^Jђ�"�I\J�JS~��a��P0��Qc2�]��X��V� �J#\=���#ʉ�m�up�El���H^-���X"7w�W�t����.��a(iH�o��9]>X�.��t� ދC�
*�ʲ�s�T�:Է��]\�%��	K��g(5
�υqpE�C�"��h	��VН�n�~h:��RpY2����\�9��X�kMN��4*#uys�H�6&D�2P	�?��hu���g�u�����jMd�4?@�!� %�#�\�c��:~�  ���`���ID���1W�����L@�ߘJ�>��/�)�K��a������3?W�N�����<4Z�{b���/�)�mߢ�>�3 �NW ��m��N�
,��쑟[���}m�ы>�{;׶#�i�>kW��픴���:,��&r�O.>1��~{���_	�C��cl�&"#�+���5�<�A�l&��R�Q+B?�N�����m,���׎ ]~�=]���$�6TLJ	X��C�ǚ`.+�\ ��␱�8����D H������A�fܠ	�������Ԩ)c��)�,U~[��5ed��I� �t�� �F���vK�Ш!��Z�Ʊ��zՔ\4)C���Zn���~s�aN�`��������G2�[͒�t*�Ǖi���ji���D$�0��=��3u�_��yC��m�k�ә1�j�������Q��
���=��%�N�{������}�w�	l~�T��G���Ii��7�O!�>� F�h�n��#�XC���M�gݗQ 2U3
����w:�=�Z��=��\9�G
�Ka]x�g���p_�/�? �;?{&��8�rk�Or�DR�qo 10z)n���g\k��H|\��2��t�I�AvG�{;�#u�#�l3<�_\+���>Oo�Dz�%�캇�0?N{�`w��2f��2�e]a��:�_)����f��_1��R�7�O���Ӡ.�m�0�Hj�t�����j%.TB�k�~3��b�TD�U���hrΡ_�;l��?OK?�kհ(��#���9h�B��,	��N�h��k@����(+k��0��Jh|��iP��|�a��U��kc���5�ඝȼ�%}��~h��>�l��I��|��HB�w�?��>x��`F�xSIg)	e������8��;ǘ9%�r&��C���]i�DI��D�v����V�*�YB�h�>�~BW5�cƮ`i���,8dd��~��S�M��Q�Lx�u)��ɳ|���
����ƾ��<,�d�(;aӻ`�d�K�Gd}J�����窸+GA���e5��`�_t�ԕ����;~�\�'{���.�����0���6漘������؊�Z�_82��-' (n�����`��326,l
���q��'��:s@{q����;�|�d�^��4o������՛�.9y��[���#o�wً���x���m�*f���~R.}��ӓ~�ꂸTt������Ԓqݾ�S�	~���|�*0���Q͹���1ۋ���_ u���B���{��2;)s��~�)�oɅPȼq>�ܕ��1�c\]8�Ɯ��%|���Njf�1lZ���z{�MS�KU��La�h�E��e�s@u��M}�2�|*���e�R��]�0�{�nB�$�XL:e2b~��������s���?�>/4'_�P�Ѵ	�1z��,��[z�tX���7�������8�[x���(�I�z�������m�3{bq]������tK
k����p�6'5��j���<�D�|��]�<)�1 z�΂aŉ�D��X�2��L}�b���$o8�6��o�+Es:�穿{,�Qh�h�>�")�>�nkq�b����+�cA���p���\�1w��ȉA��`����'U�]�@�ϳ�R�$
g�8$�̈��9�+�_ՄS��T�|��3�@ċDr��2GR��l&���Zv}/���>���;�c���9��(}�ޯ�/kN��j�Zd�~��Ck�6��� �.�8I�
�+�y��<�R�F�S��<����^1Y��S4~2Y��0QjFi����;�M{>*�W}0Յ:�mÀ���1/�}���
�Vm|^D#��÷�KocB��b�/��!dH9.�r���fن�h�wݺ>��N�s^m{Ww�Cw3�^9��m���ׅ�}r��1����b�-�$2q�5�mY�5�$9c���Sى]�����A�����G�����M����1��ťN����w]u%C�6�=��Ţ��0�9�͢���2�	*Z��ܧ�jU���-��V���βK��@7ǉ���:�Ϻ�~���81pG�Ө94N�R�z���.?�w~nb��-��r(�;5da��=�0Z���r��p���TL��-v(-�`��(	��6��Ky�+=�ʖ��b�xܱG�)�p�:���&����l�\��a!x��0��77@�4��y���,e�K�i�r� ������\
܁�n��_��{�]֧A��i���Q���ӗ��q�rr�_�?��M�s�����h�t�s��?�-^�-M<"!�xPOd8�5��['��%��=�W
ڞ!�t
qZ�85��YɄ���*�d���8���A)���PI��*����74W.��k�L���S���N?��D[���ʀg����V��Shs4s�tj�|��ٯ]�絎=����33kڍ׌��y���^����*p�� �:
mn��ٔ����Ń)�������eu�(m�H\xR�s�r���p'�J���q�l�g�uI�B4�ob��CrCO�a��V���^�����~ܕ�d8�+�f�JN~�1?)�!F
\A ���<��߮$����k?񲲟����M��>IB�+>�#��(���K��>��M��S�\�)�qb�����4g��,B3��x�?w�=�M4�1�k��6;!<Б��]�؀NHAy�I��J(�'���ň^�e��%	wL���9�D?Pq����������X�<�b`J\���+��5�b��z�8˲é��&(oQ$�7?��+yp89Ht�5xHbj��&���r��aGZ��9�?�<�����Y���.@��jG�b(S6�fyw����n��?Z�X\B���C����˷�V��sD
�/N��3������������H���i=�s<���Z!<��Nj<��W��& ˤ��י���G�9���V��O,�g����|��<����wj���?_,���麒뱭��d�e�Z��:�	�;y*뗐�)��GT�H5g��u1̽&���b�Tjbbq�� P�)!�iJöސ��<���ש�vE�R��mTW��Z�[o� l��|�B��ߑ�yQ
b�� ��Z¬����.n �}u�3���)0(��S$���Mb�%8Bφ��ji�dc���#���P��8+��Ľ���g�!�I� �2��L�>:�~%����$����.+�q��o���y�(���n�y����"�)�Q��Ř��_���[yOzv����3K�����`��'Dg��asK����$�3f ���]�uc���sdo��(PF��J��$u�%v#x��nf4͍��D>�������.ț�'-Wr�ڞ�������;��2����VU	2J�0��0r's㑤XD�5�$��N����T�%�0l��S��ϑ��	�L�h�b?<�-Q��᪷��H�r��ˬ�/s�b�"�dtz�I�Ĩ��|?5(��Voz-���[�nw=���J| )�F��/�i-�K �.:�{<%��y�]hS`LcP�
�K_�z���<C:Z��E	mX|��8&O��.�����\�$�ރ"��,�D��'�@���w%V�ͣY�]�@t
��M��w�:Wf8�@�)���X�ZZ�[�c�D�Q�a��Pc�j-:w�H��y���/��� zA�|�u�<���2�5�W=�
Kڇk�F~���]%�|�8|����K_���5�/-N����D��n���1&҃H�AH���5Y!�����_ '��٨(��f~�f�H��(�py��Q��fZ�G��F�܈F��)i�����%/�q���dI9�hn�H�*�>[��h��� ����'(�%��__�-��~:�yF�G�A"\���V5�zQ��8�g��n9����u�7��0��o4h�l�/�y�F[2�$�8 L=r����r�֠FG_\I�I�>���d!\�;�eP˴�ŤWf��X��x$d��Q6��%����8%�y�,�8�)�����D/3qo\�Kbc�������if�+p+�R�X��v����}8�˘�nh}_��V��6i���Q[H�΃^�aS�W�UK�,*��0#z9�i��$��q��3v�4�Ÿ���z`C��v"�˦���[�ںEL�����N��}�hH۸_��O&�Vp��A�8�<�F��pF����B�X��R�J�\ݏ�׾B1ޔ kq�g.��z�\�E����@�AC�UK{}�Yw�=��5~��А+Y��8��
!�c�eͣW(cT4T�����1�){��vv�9�K��J�tskKJ�svZ�ӆ������%�x*�@���P�=7����T,���c�3���h#O�MH���`�cIA��:_
O#N�B_z|�'�>9O8yȡhn��$�W!a�������qɬ,�̊�Q'٫
����ޱ�R���>��H�o
�x5@��0#�'[�e�y���Da[~�R�C�6Ⅼ�=�
�sn�TH`z8
_��sz:f�lf��R÷mAJ�R����4~!��Ys5��k��('���͜��Lw��[UJ��2����b����|���3@%�ej��B���\mZZ�����sR�M@)P����0�㙃jz)T�Hu��9c4
�%��Ò�W�.��B�����;
*�cw{'e�M5:�[;��cOG)�C�2��WX���ik�P�����q�� IM�2���:~�>�D�4��(�9vIdzAc51g��xr5����=�ɗ��kg���CF�Q��þT���G���(��p����"�8Z��t9b���L����\���#r�qN���������.B ��"�}�J[g_o#�Zx�f�I'-S��;�޳Ld����!;�%���i��,��`k��RRe���: �o���#��`6́R�OmS.K�-g��b/�%��j4j��"QR�D�Ox��Q�!��zx��hjk��x��YD�MB�ݒ��F��ښ���`�<�s3�&�`����O;���nU,��1�5&8TJw�D<���p�Y���X5��e'�:���i.���M�=x�.��Fѳ�g�$Qt��y� ��Y��Ñ�-��y"�j�c��n��g�7��J)�In��>B('q@R �[����P���m!��=��=�K����HU����}#��A37zQ�� ���4c�'�,�R�9��?�71�s-�"%�0���_W�7
ˎ���DT0=�_���l��"5�m3L�ó��N�(����nnWj��� ������+s$r�Ǹ�Οwm��Wt��3^����x�r��c$Sf5c��1�~��$���`���A��$��C�⹉c�N�Vy�wYR,��9���;�א?�0'�n�ub����D�6@�u���a���2�D�V^-Ēsi�$I��|���]�O��O:� ֹo���S�P�=B�8��ȼ)V���t@��<��}�:i���@N<<c���򝫠���ScI��z?t&�zx��"��ծ�Ll$dT[`��H���Qr'�������%��sTjb�Q�ɿt��p��5�D�VL"9�,��8�ɵ[���r�	� pZtb��.@��we6h���$��WNN�¡��|03��نӮ�)�a�AW�D\hAΉ���;\%O蔫=Cnr�7v�0���_@�$�5n�U.<��p^MEU�#���.�:��0��L�U�F+@�G��)�G�̫`�Q?�:��͑/��t!7��%/�(�	6�2*}����o���N���I��mb��Zl����C����><u��(���=�[	�4u}C��Ά�!���O��E�f�L�s����@���+�A�DGA��H��w,4�w4H�Q���u{��7��<���8c���9�����'Ab3$���"�y����,�-:�u�j�v��������k��iyG3"�,�%��F�o����i���b�]�=6��8�VZ*Ŝ���^��Y.*��!��h�9GPh����%"�������-e�֏Y� 3{�B]���\�JnUWV�6�AY�w�����;P*JG�Du��[��w"ə�=t�4s��d��e��G�F��ŧ�"�>jrv��������
��>+��'���O!f�1�3�����_Y�G��<m��Ia#�.�!'i�W�t�j����@v�̦��Zc��ִ�3��a�����_��*�9ށx>8��ђ&?���AB׎�;㽬x�Q+��߶�|g��|��z��_�� �ׯi�2<f3V���q����H=(��Q<�o�e��7��X(%��7R^��?�jz�X.0�o2\G�ϼz�]�X�������i������b��1Iy�r����ꉝ���$���>�9@��	d��B�tZ��"�{�W�%&�5��m��F7q���e�o^��+甾~B�P��e�3Wi.�Ƣ#�<d���%Ur�||�ʔ��
*�}�Fb���[��VR�vLQ�� �(�Ub�7��U{,����������/`�b���C2���j�>���8�ϱ��PN�#��J���f���d�/��3v�MKg�T����c�GM�W�$ٟr-n��h�xz�������M�<9��������tI�=LH<M���6����v���)��E���x�o�~�%������XE����E��~FUjr��p+���K��Q�;ܱV�ǲ����Y�W�B���?1�u�["��]nVp�H	�(��0S����,��	�C��?��Q)tK�X��:|V��c5G��*55�������h�*>���+��uLų$h�JS�oZkm3=�:�Vwd@ݨ(�I~|(G.��½U�/.%��I��=x�@���"$`mܢ��ǆ.7x�<7�'"��<
Э�)�W�/�l�es{A`ϛ|��2���)�QN��ge"5Z݅2���W]���}��?h�����Z�%��D�ήV©���?<��
�n�P��[�sM?]$���6�c���*����l�螫[݌�!E����4�V�!���ԖS�O�Y�畛V��2j��	s��P�RKz~��5bN����L�8�݉���mY0�=�Z<)�E�m��z���5��M��E�����&X�U�u2s�O,m��+v�
��{%�ህ�D,�+�x�{$E��_{>$�nS�(����P��`@�#fj��4Kr�E��ʂ%vCOn�I��U��F��`���A��l�;� �oJ����7ug j4/��G���}�J�LW)��rp�	�����X���;`<�H��%�\�� 1S��
Ix:�D���e�&�}���ӎ��7l8��{`���������D���fDc$az���ݛ3��GU��	�ix!�$�\���p�es�v2��W�ó�j� rLvoC9�2��o-�a�N�*��k���Kd��^h� �h:y��w���j�kd+��/���KJs#�����J�����ډ�3e�%�����a+Lz���䨹�A>\"قj�W&	��|e\��S�� ��/$+���}A�@�i!P�y����<��b�����GZ��&��x��J�w��lk�U-׈��r�A����N/�!!S�ҭl�d,��qGZzV�Ƭ�(�hVn��0��.v��UEi�����4P1-�rv3�� CR� 1�r����r��Ex�>�磳M��,��F�pJm�A��,IR���K��ԓbp[&C*֚R-<Y<y��e�D�2D|Z܃���㫐-�io}��fL;7y��B�&�r�=�_����Tλdc�ҋs���![Vni�AE�%]�s'[�xΚ�ऽAS^�S�24�����Td��
�aVP<:����V�͑2�Ɖd�c�fS�}c�<Sy��MO������Wɒtq����_��lr��S`��c��+]�!޾��4��j�-�]M��v��0t��ۋќD�<�+��x���z\C�]cD����'j-K�V��E_�����w�j�`7Ү}��Ѿ�*	���b#�u�$U#%��7�_O���y�;4���e�?|aۗ���n�N]�� ��S����i%r1�r��ȃm,0�"ڛ�۽
���;��l ��7]����b>���8�~�_��ʼ����R߆i�h挰��'����uV����pW"�,!y�l̜���5�Q'����4��bQ19*�<l"\�B�<�O��ܘ�a}-�S�O����G�{����8̈́3���]$#T���?�upƻ�Ձ���+fh=KB�a��g�C=슏׹��V�ox��d ZS��fwl�=��)I�Ʒ@��d6ի�vhQ�T����޼M��?~~��t��v�Vl��W��^��X�u�λ&{�2�⛳ޭꕭ�����2��������_��8p�Y��M�8!�U�M֜+��j�/a��O�*h5�u�9S�o�Ha����I��R�u���P�&��"���w=`l�"�Ww��FP������5�m͛�֑��VnKC�O���S�FM(�>�ȯ����%ؤ�O��b' g�>�,i�,E�Lҏ��d�X���?�`/K��ekRi�t����tf*�Wo�gA�pxI��m��s��TkhN�۪��S���e>���6q`���dH�I7�z~(��%��)��a�{������pF��0�@v1&(�H�J����u��O�^�[�C}��4����N���>,��waRP��j�A������)"�����E���<���Ő��R�@`��i�d�#^.�;mĞ»M���� �W��=P�m8�/(�ɽ��)lƖ��ؑ�V��:��G�Nh�&MV�ԻS��ޜ��=�0�C�`�	��g1=M�q�
��J�o�ɕ�֏i��z<���,~d�h'	�����kpg������%9��VZ���Q�)wR���@ @��o�(�?.,W���U�kl��%�0%;�,�ԋ��јQ�!"��仈9km�A;��m<h��z&�Jڗ��ş�)�7���Ku�Gp��"z)r�F���G�.��;S�7�	]g�����ʨ|˵���R�����m��H�R%]��q�D3�ܪꒌ�������� �C�P%� �o��}\I��ɋ����0�$����� ��w+�~[�2u�N�O6cʙ�����`i�$�ՖD���=�0�`�8�7���x5Ի�G�n�v�ʆSf@co����9��m��$�A�2����9d7b���Lz��FQ<��D��Z#hŨ�_V������OFdq�'���hD��s
	)gw�F�x(F�X9ϧL�S�LD�$��G�כ\��$C?�U�<$��nn��f����iu	m&eH��!��j��X��Np���d�~�~���ӯ���V��j�IUj��?'��Ce@�)Lv�p�<�3��L�䇿�{�����T�Q���,�Q�09��#���Z�\C�=�V4Wu���!-��[%$�b�F[���A��_��C�ꄹ���8T��;����9�(��a����:;W1j�� �. ]S�U��U�@)F�k6��P�b����+�=�fS���I��)��OB*G��V��q2W��z�:M���nQv&<��M���B�
k3�k����6�!���U���/�d�9"��^�8hK�N��%���&�h���U>��G�q��/���
o$���fIx��V�0�>�8Ðe��UK0�ǿ=�9���;�?͵MtG��c�i�S�%���,cV����x   �ZNl7��u���"�8�g��oШہ�������F�}8[^@���͔,&���Y� lenr����d�4Ԇ5��1�����p�x�����9���%t��<jGc?����S ��F�&l\�>DՋP*Cؗ����a�����]�(�w�"���� ����H�9���B�t��=��}�fuu�I� E�(���8ک���Α���,�RJj&��hd��o[��������c��ᇒ�'O���#(�7O�jL���dbGc��=0����X�`��%�H6�s�8���[���y)Q��Sn�Q����`Ww�$n��J9��m:��\4��j.��c[�X��` k�f�y���`C�tj���*�1�Bf=(B@j�t�y]%_�&��7Tެ�r�ڀR���;���k��>�����7Y/g���(z��?�6h��Sd��W�	Ï���Oo�`�(�T�r��ޟ���fD[��p�ɿ^��B�EkbX৮�O^4��b��y����Q��j���6l
�̃l����q�@����'�Q[�
@��Ɔ�&��3��T��#ؿ�o�}�l�Ǜ.&-�}@җ-ÿ�ľ�JG(�@���d���C3'��S"\�6l����}Nd� H�T���
^'ClHj��SQ�c�"�F3O���i�5fS��Y��i|vc\lk73�\��'�5dv3T��of��y1İ������~���4a�*��f��%�p�*H�ۺS�̟||z��L0G}0~�C���D����*�jӭ4���jgXuk6�^��������d�ȇ8H�
�Gf��K�n�wC�i�]hh�ԯn���\�V���7g����\p�և>�7�*�Եߋ�&>_�����A�$�s��٩TpZ�A�]����Ϝ[h��E�7B���y7l��:5]�1�=�{a���a�!;d�#vS$�F�������D} ݱ���LW�͂�U�U$���sF��xF�!�}�M9C306/3�s���Z	n�`8����hP:8tg�����^{%n�	)�'Xg0-���馤Rͼ2��ATS�:%tݒ��Y�'�ggVx�����%�������V��x4�9Z����� ������a¤sR`}W�|� �"Ƕ<���֡it�o������٢�h�$
g�S��FsZɗ�N3sܼ��x����5��^[J_�HF�P� �QG��3��b�_�����1q��dK�;�aӯT�<��K���^�$G>ly�u|xu��Cm��H'K��p�wD3�.	�U���y����m��U���#���jɩC�\���X���7?�%n�2+�p�"*� �t����~V�H�,��)D�][�/���x�t�Fj���":I(��5/ q%�>�d�� �l}��W�o5]�?��՘H���?�����U�\��Sn�o�w�O5@���M�4bِ�իR�gvA0�����J�i��L�	x
��i� �V�aPl�U��hL�~Y��&��r�{GNh1�v](����T�2��[�{a��X����&{!Q�3R�7y�	h#;]�ؘ�����)�/
s0]O�'���F�=�#�R��!a��#��m54omn��_���ek�o`yJ+Z���6ה?}s�.x��0�;X�`��fh�q��ʥ|g]�~_:U��n�愹�s����F��V�sB6^�QjF��h������'�Q뤈4�j��tF/�fb��2$,m:ы�ڗ�������L}�,�"�S��b ":v�zǝsD�����+ގ�����HNO��d��M]���#���B�B���l��s�
�K�Z^��,m���Y��5U5��xO���f�e�z&��$�����X��RP���J�~�x,;�����#�	:VY��[��h��������8��/�HThh�b����-�S�A񆄻x��s�2B��if��F
?�[��Z_��c ����0����k0���1%�Dс��#�J�^�r����+��p���U���+�8��Y���4�q��v�{Y��*�4��%��@ +b_̞��K><�X	ɠg���-l���u(�,��O	[����[�=ܥY���";��g#��W��k�z5��ѡ&��a|wI����*���~j&�'e9sf���T�1�����=����t��[��ikRK����G�~-�MQ��*41P%��(}OA�4�+��Ta�L��Yò��I�hQ��7��s��jũx�.	�W(�#��
��3����V��-�Ō�O3q^^�9O�ɔ�;I)�e�7�E��h/��h���3Н����i�Ԏ8k0a4�=�V���/9�������>�6ǔ ���T��V�{ؠC���Do���/ש"p����Rr��'�+��<�S�b���L��(� H�Л1�s[Tam��@�7x2��Y�ϕ,������LMk�Q�
4x��z�o������.��i�Ձ<��K�7����D���Iëg����͍z_���x�p������X=��q���/GC�)w�����=��X�K=9�!���e1W.q֧�u�~E�?����f�M��Pu�#þ(%�a����ܛS���#q�<�n^���~v%i�L�"쩩m!�dBr�7�F�9?M4�Cq�B����J�a��b����B���?���~㴛rZ�������X���c��,��D���/Aøc|9����h�����S��e7^
fn��H���B�`�,��/GZ���.NqI}/֋I�@<r7�jb���(�1BG�5l7�7u{��>�i��|���L���ē��ؓ���o��&o��6��sl*�~���OHt�6��'�-�gNHŦ��i�S���q����X�ҽJ�D�[�q[�:�d={�8`ސoh�U%,ٷ z�T��&x��a��ԖA�m��(�w^��5��|I�_�@^n@�vj�g:���&��p�qHs;��{8��,q��P/3G��ㇼ'�mܲҨ�e��VC@�H��ݢiF6�.K;{�5lU���1ߐQ��+8Q������hCz��a�M�/r}:��+d�:
&�|�;chj٦�y�254���	�8.*�������6�{C��^.qX�
9�<�;��\���ˣ�s��a(�/n
�m�����G|p< �Gf�>�N;`E��j�4S���)R 8��Gd;{�9�j�h��_����NB}7�|�n\r>��2'!�Rl��o��7�Z���>�T��LG�
�`���XF(z�hf3?���4�NoΛD�ɭ:~�ܩ^��i�2<K7X�<q�Az���ŉ�����4y��4�9c'A-�;�j��ns)B�Ҫ=���~�g0E�p�=�3ҡ�w���^�#�:�u���������c���&b&,�&A&/T��
�|nw��G� h`gi��k�|��iy��P`�߭�"K��Cf�H﨟ZY��$��4�� �l��E��vn�Ti�ZV)1k�H�8�3(m	��l�
���I�Ku5��Xs�@���8
�x�^3�R��L� �?��IJ{ט|���g���h�"�� �ʧF������z�^�XbkQγb������C���r/𪨋-G���=ے
Ɇd�ϔ�����N߄�\��x�����2�Gs���6�����M	v�N%��n2Yh|@�Uæ*°�2�XV�=�:�
z�YkN^V0�س�ە�|�ՙM�I�JIg?��j�~�g�y)F����Vl���y��3I����@NK�n��W�'4b�.��n;�o*���>_n.���ڵ83�j��K�d�K2`�j�ϊ?a�͎l�(N��k@te#;�OY��%K�q�����U����n��_�@��mB.!��[oZ�i�%L�_��Z�
JЅ�|,���Q`8��H��js�䒠�B�3e��@T\?�h��X��ً�ۂs�T���q�V[{ˑ�.Q��N��H�ff�dU���e}u¸����)k�L�w�����X���X��@�����-{ݞG���Dq���{�Pp0�����)��=�����գvO���8����
�
G�u�=��`ȇ
�I���>`�*��AkVI�g��7�������17�n���=O#>��@�S��]]s��F��>�d� �Y�	n@c(f�[蛄.r�~+��s) �ьt
�.^h���j�H�y��C��O��_�k��}Fx0��嚅�0s�!3�dt,�͓�(�+!s�H����DK�Z���⺻���Mk��#��1/��Ј6W/2�2����H�Kf[�Q	��<��gE`b��&��}ނ�=`�H���?�Ӷ�4�������kY�)z��W�˲���_���C:��Q�=PX|ȻG�㏖[�x�1�-gP��ϛb�8ͩ���Bݐ�nPhY%4	��^�4�V]�	�5|{�Qx��K�Hpw�^�9�䬈.���vrF��$�_lB�5E{A<� ��:�n͝)ͤ��?z���ܭ�:T��߲e)��Cy	��j�8�ivLC��ԇ�3 �Y2Mƌ�o�>�L��� _���7����g�	�wq1V1�Sl��5��ۚuS��U
���ʁ�:d%��M`J�)��ɕ����oG�õ��X���V�mP������ޛ5�����n��a��}��5��:�r��O��Ŕφh[�_��4�QR(nZV��#���`�g�>�V&CN�ޙ��ؼV����c��NQ"nM~��y�V�7G	��Fy�Ja7�x4훡�H���V�&��p}
�a�u�TD��H�8�?����I�!{\��=pH�3�0e�O�V�F�*�/V �5�e流�𬪂�R�e�'}9��@0#V�j9L<\06�O�0��B�2�.��`�R�q���6�
�)/�A_U�F�n�EY�!'6�j��'��~/NtnP����!uG�!�1�8��	D�,�n��H3[�6�����J��a41��ڝ��@*�T0���o����7��O�jTY����Z�k�b��^�ZZ�I��t�h���Q<�Z����,Ȑ�AG;ʷ#�C�\��h߭/(MapVX�h)\��7&��7��QҐ�̞�/ڎa[�W;�86Bz�	�����*^}��/1�KB<[��Fl
W�/���}!��G8�����x�tkѲ]�/v��xX0�@HO�#h_�>2�kߠ6�6�,�
�2��=��ݙ�َ��Ke�VTy@k�[E�JY� APT�����*���:�0h�1�������|?����^��k0�UR&�i���(��*��՛ja-q|F�Z�6�;�!Y���AD_��r�E��r��q�����S��׸��-��+49���Q�n�L<Ǎ݂��"��R�K�B�Z���<k'^�Q>7q�� 7�nCtG���8�x�J�9/�#i%Qj+j���F� �IԎy'�nc���},K�@}��DL#���Tflw�t��T3f���{k^�OP0ˑ1�������� ��U����I�� ʽ�2��星�$��'f��G��"���]3)B�?�*�pXE�����;��h�id��W�2�03���dd�V��A��_7�.ŷӖ�*)����`w��|C)$;3n��u��g���B�md����:R�9m肳�jRC�Ð�����1_y�=�/Ƈ�׿s�T*�P+a**4�[s��8����
_f hN尻"����J咍*�W�}bh8���U�LF�ԗ{8��cS*8��<f4��OgU:��$WD���-��z9�gС�Jy�A���۽r�������z$��0d����Tع=�f8@�݋��@
���bn��$/I��e`d�|�� .����k���;7��?Bn�Q)cn�`d�r�°bΞ�&ys&,h��5~�Ipa�V����P$~x�!d�MrU,,�9Ƴ�)N.f��-��x��΂�\l���.�tSnlʇ���}�c��T��U�}[j����+����A��Q�zBt��e��@=���ד�H˽�9'{r��|Ct����h����?���ȼ��j�X�9S]?�̠'���^̐9l��^	<���'�m\0Q�4RU=�q��׿��QI�h��\!7r����SY}�\����C'RN8�0��7*�l�k�t�_�Y1��$��J���ߢ[�j�V�\�?R��l_��N�g��{G��X��G,�
�n�%��Y?&һ�
;c���En�*��\G8���pA'��m����#�?3ځ�E%�|�H|�5�bG�u���4#�Qcb���\�Hf��&i��OD��h�tq��_W�b*:���8�������t{	�8L:�b%>Ҙ��0SV��:��I&�x �([X��Q�W���%��0(�_L��H�l%V󶍒I�=�N] 
K�1�-�0j�NV�f^���Q�"�U/�庈H�����V��myB햕|�{�_>8�t-Ér���d�� �"�rDKJ�F�2��f��,y6bv�Q`N���e����9 �_�l6
��[�ͽ1��+fh���"�h`���Ϩ�_�%�Ֆ���.�y���1����NT
��l#�����z���3,�
���:Kx>��qZ0�~Z�R���ο���r9��]�𗡽1�ɡ��(x&�#�\ˉ�j��cgl<	̔�Q��d�;X%ū�w�\:/��s5��[���bB�g��$��RE|44T���Hь�R�3R�a{j6A�P�6Z%���ݤ�kV��5��$\�b	������
���?������U�x�*_�}�Hz5װ6��%� ���ոbr��:�q�F	��+O�)UBӦ(}8ųk��L�7nѧ�o{��i/}��(�C�ݣ�v���1��.R�h\H${�Z�e�� �j���o�f�h��t)��;T
�3\�FK8Y/D���V���ʾ��]`�Ak��*���¡���R��KЮ�4�e�0��\��=}l$]F�� �`�^>{|ܶ߾Wf�E�]$�8uƨ����Y�,뜞 ���83P^�aT�^��_��1����lO �}��S�0���i��P8JA���rO}�st�Y*��N�92�!�E�����4��� B,�����z7���	�����i��Y`K8�+����%�'#(Y�9{���d�'��fۙ48�>k��^_�4��$�lv��D@�l�'BǂȚ�h͙�a#3�{��V��P=��/��C���(��س�4@����t�g;7�������v�O|.(;}��TƝ��&��%u�<����T���@��ěEFn�����9f]�y����<�r��Ѣ��'�Zdr��-�Zx�</b��u�]&i�y"׺��Uky�?�k��e��f���pz|
�D�B0�*��	'恱y���'`�M[��[��I�Ӈݐ�n�Z�6��N(�M���Z @�&c�D���X�6/�M�F�G�?�++�0��
�wn��Q{��dZ;��}6�w��//]*��ge�ƶ��+EL�+��(;���\]�1�[8�k��H_��R�;���hH<)������m� �wj	z��H,�U7��zr�3���4�FdΖm�w�Ǽ�3"�\��l�$�[��Ni!�t��n�_wBX)�ʲ1�cpM�Q5�-7ZLwK�p����2��Ĝ�<xi�ˇ Y�2���pV����'|�>����mF��d;�t�V��!:yD`jZ��V�m�p@�t (�31T��A�*�8�:�נ��������k��ݪˮ�PAݖ��c�)�͉\��8l�]ze�#�z��l+`�ǵ<F̸ݸg��R<!X��X�dkGv�I�$��Fz�/�@FS%1�2Bt�AJ4% 3�|H9�g����f;xNO��~ڂA=h� �������w�9V��V)m�f��l�ga��'�ge�J[kL������S{�!s6`^p�	wC��F\���U��sr�߹��0][���ׂ����y�8vp:+h*Ue�@&�o��2]E�{8��?�ş�qyz �B�����*CC�dENk~�0e�$:��T���$�W4j���������j��M�ux*���Į�������'�/��tY�cE��M�[u,"(ƛv�mP���``� 	�:��` �R��_�si5
10��j��v�L��"�x.��1j~]rA�$���#��X��p�g؄��݅�=�x������	\�A=�NܼKnG-Ї�E�0WZ��S��HʍG�z1��[�z��L_|VG�/v�5��aB��:�v]�Y��|�|�ZHB��x�9r��Ye�['��:�}J��-�ӏ�zd��b[(�R�}?g�����6��e���{S�i�5ص�ɭz`"�e ��p.�<���zXGh���ta�٫�>�R��Ջ�x����~�ZX����e�$�"�)@'�N*v�q{�2l�f�U����}5#�D�Y{B?�^Y;O@.��D/
�qţ$:k!��P�WȶA�����y>�`�<�����WG�v��pf�ݥC�'	�!�r�b�{��xa�����	��BC��s�2����)z�8m�U��@/���hA˥�~L���ؚ`H�%��v<���Pl���RM���& u೏�B�l�U̍��j��8Y
g�ˢ��W�}A*a��r�Ǖ���D�{bF��"0�4��m0+���֔ $��A�߇ý_b|��U 8�#CuP�D��v�R�4��v�W{{�JpL���X� �<ǭ:�g���9Sd��R��I�=��������T�^�>����?҅o��'N�"��I��˵�!����5+H�i�$1'�
]?�l?��J�c�u=���$�Ӻ0D�f�j��
Kv�J����0㜘��S�s!H�r_�a���;�R�%���]>�S3� D7��VpS��۬��iu�NqO���i��	g+n��4�< ~Y8"Pic@N�Oш��lX��g<;
wz��M��VK�㖜N�̋�i?����΢hu�eD#�7�t�(��q�Ȳ�L]�����v[�%LX:aќՀ|iw��b���Cjn[4����7��C���*���b�!�f5�\+��P�w>P��@pRH;&Ah�t�s�[�����ր�w�C�f&�J/$�8v��T_R�G�l�'2�Xi x�%�t�����웊ӆOq?�J����`1b���~B�\<4�a��d��$��U�g�ƴ�f�W����r&WD����>�g�*�R}"U,��J�9DQ�o�qw6��� 0����>!Qq8l��Y���ʇb��	�}@_����11���8%��4)c�\��D��nՒ�@,7N�=?�LKM��S�̂7�R��d�Yu����m4;�x��o��a�<�ı~E�a�64=���g@1	D��Zv*�M�熎0o�g~`��BڢU����E�&��1��|~�x��{FO��D��0�ov}Bj�I&oϗ�2�m�j�	��m�섑��s�R}ʻ8��+&Ü"T�Eʇ���z�J-��Z۾��sc�2_ �4A��aަ�4�%���9�t������y�X�i��P0�<^��hύ�qB(ΣXq�ƛx� ���@�J���^5�h:δ2�S\��螐j���C�ֆZ:��v*#��������8�f;*	5(�雲�r���F������!�Y�';"��$)<0�6lm��A=t�X���.I��u,w�k�K����6ތI��5�������&�7�y�'�O0�d, ExѸ�x��3�������8��J_���iZd	D��F[�v�"�h�P�,�y�bԍ�OTƆ�<��}v��*��}�޺/�ΰ��B���?eє�w�h`��|�B"�����[{�ob�V֋�k%�eB���o �HhC�[ �jJh���?�Y��K��_���TB��/�X�XZ*���`])���{i��P�s���U���%X ��@|mTbp���{Y�����C�b+������8�z/,�lo20d�21�b�ȠC���s�/+)>y �?��s��஢��Z>〺�Y��4����7[q@�<��)/�)��%_���?�r�;y�_���"g48��}��E��,�L����C���Qo`\ht���/����w3K�C���V�ژ~��"0j^�S.��-fX�[�X�T*h-���`*��F~)��w݇�.���j�~�?|J����8�r�k��,�biq���
8l���F��K�|��ٹB��0�&_��:���v���E�C�-(!-ބֳ��G���Y:�ei2��w�Z��@ T�<fèN�RЂV!z挈3�;��L����7~Whp�XqWA�%3�!.�~�rl_M �L^��D�ؒ��J!��_�=�6vA
��CtfA����ŭ�{w����v}��G"J�k?�A	���p򩙩^�+U�����R�}�/4�gP<7��m<�<�:�BW�,�%�Gr�T#�C%�@����.�'��㾳���\��5���R�[��g���e�+��s��)��++�I�A�֚�H��0�!`�wvQ�j~��z�c�#�U1z�z<U&�^� ��!sȴt��"��֫,���!V[P^�	�n!��뛪�׳f<�0�a<��������f�[Df�;x�����_���ug���l`�	Rw'<E�{:Y��aK� ��Ǥ�<�l;��&xVR���a�ikp�����G �	KCӑ�e�<fU�,�T����Qٿ���q�=�Y��g�(�Orc����Fk o m04���/�/�8hT��@U���h/Ĭz���'��N�u|�?!ٛ�07�ZQeI�甎g'�&���cW�����r�h%�Էc�?~����Cx��ӳs<�-�vC�K;q���m���v~��ӭy�#��e�c`A��9gF�{�R���M[�]���B ��>e��j�/���tg������(-��, U��?Χ����K=��W��3ېT:���""*�`�5~���Y��0�=!�����v�+���(�z��}����%G��o�� �z��d�����ivU�ģzMN�����w��Z�蝑[��~ĵA�2K  XW�`��(�^�+:��l�9�e���qV�+�y!��!^��pK����r1�ĲYúH70�F�X�(�4�<'L+`��&i�����t(e��j����y�{3��+��S(�A�H-�J�w��5ϊ��r'V�P����v�D,
/�t]��o:������\��^��S���1�B�X���=	�����DRÝ5��U�ba���kAy 0�R�\t%ć����BB7rȘ���z�&�TK�VZ���喐��G���9sĆ̎��Z� u%W�X��s��SIC���$�-Q��QA��e���l]�٣yg�p��^��tZJ�Wq$�p���R�l9�s����})����(��E��V)��U/�VA�ũ�q��="?+Fs�ݏ8|�Zx��W7�/j��!]��b�����j
>8�0�CV����׾�� $�c�a5q�&�۟�@~ae�Zdr :R3LHo����͠�o;>��17O]Gt��v�L��o��a��$IPu�m{��Q<e��:UUC�4G��*r~jXud$]g �O���݆�v6Ծo�#��P�>p���G���GU�kݿ�b��W3MA7,QFC� � ��*�󹆸�L��S�����<5�rl���L�jb�������=L?�U�U=-�9���[�j���]�urX����	4�=F;4bR��ٹ�C�5?�,`k�c'm{�I|=*�?������|E��	��Z��%ڹJ�3��^��OZ�(+�I@�p�+�V�7��4U/r��/���-�
2�b�����E�9��V���dD+� H�`]0�߻� �QϢ�\�.�2ıG+�}X���AR+�7y�Z������ �i<�����痮����a3=���@�ģ6��AQ|c��L����؛\�[���)M�kf�P��d���G�݋c
��Pm���J�a�7pH���1]�n}�݋� t�g���q ��~)��;����,��g	�NΠnx_֩�X�ktF_sT.�+��>m_c�+������85�?W�2j�%�"�Y�Q��a��ٛoK��W���,,�i�ȋ��w�|���������=#��|/����O���pJJ[�1����]^�0܆��"l��[81�F���>��9� v���\i��t�6vd���;\��	�m;#�	T���� '�G����>��㢕�|s�bb�#x��Rg���.Lq�̶x���!$�5������OXŴ��.v���D�%�������Q+�!5m���2��Fg�ϴ�Ѡ�5��d���H^f��f�GA>�	�Ǵ�?8��p�Ŋ����]tt�H� b��e�3�~����2�]A�┙�KFH6�[��*�iF���;nۖ:ٯ����Z�\r2�����3OxEm�h36��;k�4� *��X�Lb���܃F��Ƀ},���¤Y2�؊�}(�5V}r�}W1�I�s���4&
²;��F��o>Qὸ�{Y-H�Mx��Y��Y�t5��tt:��0����)K�c	A�K�{	��#�>�׹��		w�*	�/�f�d��	��"�>Y�0�z(���Ԯ �8����b���=TYPͤ�>�鎧Q�(�)���LhxG�h��������5{��o����҉r�&c@x�����]�5þ6SEZ�]:М|�HƊ�%�ϴ��6C1�'@E0{����?[V�=!$7�\>�o�#@�=��ʯ�DH�%�i,�����>Rsoi�t�d�yw/qF;l�w��7�H�x'f�JN��X�r�4��a��ԉ(tӒ��.Ω�;1y��/#�q�~����l�jʳ�-/B/P�	���p�An�l���JqN��V�瓣�y�ou��L���$�Д��b�q`,��(�˺���Hfq��9�������,�[W<���^�1U� �f�Yy� )?��(s���8qb�D��Bp������M@�Bܹ���"H����i�����ea��iU�H5���H+8���b���!$KM��М��)�TWl��@�����(@ƵyK[<xV�.j# >A�S�$jR*�K�Z�+��q��z!�a�%f����_��: �����>\�p�^��P�5�:���&���IB̤V��r	:��tə��AW��XN:����eJ�c��+^�3Y��M�J{f��k�~͂"B5	�~Gu�]v�蟙x�/���8PѿϞ�̮��������g��z�+�F����i5V, �\�XSs��\�?��$�]���le���Z�`�h�0��|�*%�_�����e�i⃂8���o��Ә16�(v��wx��"24}���[)Q2��)[��͍�>7�$Gl1n��BF?��>��������K޾��˚���wʒ���t�z��k�;
�
���Б��YC�<��GP��6 ��Az�]FoT�Ѱ��2��Cl��L/���>���p��AdR�0^�!�<,a��"y�n�w�� ��ohT�iqA5>2q��>^�5X!����>3��t!M[��W �?�U5ǔ����/��OR�E.�/5�j�
Pn����t%�n4�����'�!��$S��f�8:�U���Mұ����,_�cD�ѱ ��<@��Gj��ێ�rW��W*�,�����3/�r�^�j����ƨ�n`�8�� ��:�bP�>����Ѭ���Tڻ�A�ˠ��O�-&,U��7|n�a�Ĩ�C��"������a�gs�ܼ�yV�\�m��
�b�5'���	�vԼa��c 2�5#5Nd��ޚ�;w�W�7W�A�w���� Ə�/���_~�H�bH�:���M �}�nNH�gi���؅��ſX�Z)�o�>d֓NR��x�=|��om��-GE�(f�?�C�* ��)`0?�����#�I��sc��~�U�t�\�';Ika�G�ÍӖ .�ԩ��*,�1q3��|�z�<
�`c�r#��1�����B0�lb�ԘH'�Ȃ:1*��»�p}7������dD���ӿ��?���7G@�Molk3^�rc�6`c"�E�ok@�MY�a�{����Z�����Xe�nJdt�}ͮ���&vAv���=�H�Q��Ѱtid�)����4�Ed�Ͱ��>�IB�E��5(\Oџ�=�Ie'qfhEɤ�W?�@锊g����T{3l���������V��Ǜ-�XV�o���^8�$�˨]��Z��P<��]?��gBGW��"�ũ���Г<��q��
���7v�3�S,t"͢���&Y��6�@X4qg�m�8N��愎� ��v i<�>�\A�Q1�b	Ɗ�xkHXK�rϟ�$�ғ��%���4��Bg hH\�B��[7
���T5�5rε�b{���ѿ�]P������lZ�����SOwr%���%��Ήi@�5��M�Z�z>W��q�+�eJ���w���j_v�E��Rj��2&3���Y��tY�F4���VM��@c�8�fH�lh�i�#/�׬-	���/Z|f8��/�(���0���i��&��)I��*ͩ�yiڳ>��(s<��*�t���yN
򯔥xW*m��Ix`�_iS�c*�G��ǐ�b�E�񹁩�'<RҀ�*�W�^z� �����Ks�C�z��Y�w���I���)��r�c~$�(���1�eC}�MkP�Ӿ�A0_6��Mɻ�*�/0ґ������n���I�JЖ�lsW�}?}N�Bdi��\�y��\{¨i�p�X#��@}s~�����b���9QR����+��}�z��f��Q���nG�ibK!~~���B~�Nr~`؛����Ο��DLL��i͒�+w����S��p(��\Q}�yˌo�zU.�V����u�NQ[ȢyW:�����jk�����lj[s70p5�`cN�����ir8�~I��>��0����i�G������%�H�d]7�p=�uN������7��� �\��C��Y0H+(�0˛IUnl��[��C^���pjM��u%�HN�@���7��,�o!Ԟ�fm���!�^h>�ݯ�l/׺Q��NE{��c'Y,�m��� ��#U�$���1�;_QI�V��N{5qfD�s{_-��ܣz���"���eN������6+��f�'�M3J0������$K'�H���G��޾���~4?��$t��Xu,���]'@��F���5
t� {A�Kj��J��� hu�_���mG�D}*�T!�&���xBR��2i�Q�I� Q�ڧ���ޓ��el!�'��@)�H>B�]��2�rP���4�A�������R�{����]�������y���E�/Y�ݱ�u^b�w歞�w�xwYw�ƺ�<�l1j�����#����>�u�+��$º탈��	�{:�HwS� z���;;K�$�{5��6ۀ��Ի��x����kb����6lfߙ���4��!yW�dc�F�ݦ�]��
�������.�`-� �L���LnAv&a���]�Im�:��7p겴:,�����l�7b��ĵ���b	�KV�g�Y�.b��aY}��k��t4�f�$[y��9ZC����W�"�ϹL�.�G��>H�~sXt�N��<����qr�}ʔJ�o��VT`��P8�풵����k l�f;������՝��ئ�9����>q�2�����ԎQ;r�̿�%���\ X��o��dL;[N��>^	8����V�3�Y���4��F��/o8h���>�� wg���{�W� ��8���$_��s|Ѻ�%��B�8��qٔ����:��������\��?lET���<�Җ*\l�Wq�=�Ƈ��x�-/[w�à��
�2j�s�'��U��bx(4�$��m]�Xzn��C1;�R��}u��U��^�ߦ�e��G����ܦo2��]�`�,�n�ޱ�N�������7A�����lЕ�S�yl��0�uԝ��&��ֲݒ;D��F��{`���Ų3�"5Y���ds���"�D5I֬܎��5^b�e��b	��a�Jtq���"�U���:T*�:S.�c�;��^�Go��.6�~�	�L���)����z��0r�A���j�p����F��PI�G�/U{��n�D���ٔN����x�����Z|�Ig*X��@����47P� C�v�Y'�tj�%ߞ�*D�A�o�Q��7_��/"* hu;Mv71B!��ȵt�*<;���xz�����*(�v1GM>X sa��1`(�D5�<!ܙG��'[��R1��&��*��j�;A��M��Y����T%���U���I����~����?y�����07dNN��I�o���_�R�A|c�T�y��#�j���/��{� i�����E���w ����b~'����B(��XU*hf�� H�r���5]c�w׆�dR$�_���ɩsN��tI�廂�$�-;�;���ևB%�Tf����g$r�0�FQ �`E��gv���f��cBZ�[�	]��L5H�uqA���'����`D��Ｘzz��3�UF�\:o�E-k-jo?�\����V�(ǥj�I�
�G ?�=Pd��k��[Փ��~��U�����ҒISS��-��C_&�"��j�g%7'����x �i��,��vB��{�o� p��o��ʰ��@�����A���V"����(�:�rF����@=�����	��&��c� ��V��J�2�!C�����������������Z0�!Y�J %�|E��5\ħZ(98�n�*V���C_��ݲ�6�B�mw�:"�N �(�c�Ƨ ��%�J��e�ց*�؆ԣ~LV�?I8mf���Q�Yv5���-J_�/��Rf����/�t�X7�I{g�ͷ%%J<P�U���s�QߓB�7��|ކ�(��C�G�*�����I�����>9�t����K�-���])a������Q��"�/��F
L�QnpN�wP�~d\꿹�!]O����}#�e������7� b@f���ud�<*�	4t��c[���Lj�D�� ��!�@wY���)�\��D���5�W�:��Kp��om�����s3$>�s�8�謆��c]�+_���Ԯi�RiZ|�g�%����>f(�蟇��q:^e�Ux,J� �^}��bm<��>b3k0�KW�My�0��[+"'3�6L��K`"�d�zu f��f��Qg�,,$��^+�앋,2��ǭ� �m��X�/��
��ۇ�0��S��mQs��ɜ�;;��҈N;r=cL�h���矪�Y:�g1����U�C_�KR�_��qy�|�;@/=�2=_Bi0��"<ФäYM;������v�c �� �Z6L�����8��g�o�Z�,�J@M�,��CZm���)�=��ʒE+"<%:D���
R��@9}y����b�����[�'��s#G���U0�Y	Be�rx��!l����rAݿ�5V�
���o�`_h=3��d��j:�x$�߭���T��(�{_[y��Z�t�����ꀙ�N1=4�Eu�˳^�����no]>
1�A�q�-v��|x	����[�AjJ���67��H�<����ޤ�v���S�r��1�7��G����W+��h�����{�V����aD����D7�:�̡��$x��Q�JW��)2{4�H��/l~$�6��6��c1��ݡ̶]��bn�zx���c�a:M��S5�L�5�4��&����d�gh�^����y31h���h�Ʒ�l����$�I����	'T����cl!�S|ͽ� �j���*������{���>����#�-}T2�Fz����j�l5�Kܾ��>�>E�KO��ˋIX��V����H�b�E<�W�W�{f	��l ��G��h	��_�$*���YKFHsƸ��J�yis�l�01chI�ۛ���7(����g������E���|�� �R����7��OFiJ���h%��fv^� S�{��d��8�ZKR~�~��B�Ch���'�\��p�Or.���_%��`�����ܳ��9{J%PFR+���u���"x���-1��r��Ӭ�Z��>]��ƣm�D�E��i2�t+~�^-��u�V8p��Y�G�m�?���cck����e��GY��c��
�*h�E�}������>#?�|��Dz�}� �!�W��+	�f�[�pB�D5M��,�Ȉ���n�]�Ǝ�����ϚI�42��f��}�$�J����J�J'�y�PS9ZP�E�sI�0��@�^��Z��#�PGq�>}��$���(_��d�'�aǼ�Gm<�E��<W4�Z �9�F;�h�0���g|Ш���
�8P��T�0�"�8M�VO`��ІB��_��E�c��܆�9�|L��}T
(�k�v�ʷ��>�2�B���n�<��X�
RX�N�1��̌ᇟ\��6�ԫ�>q[�{E�t�HԑU�s�*�s�^8��'�A�SC�IDM����cFF�M.�(�Z�X�o�.�`6DIA;@�f������쩀�84�X�D��IL�r맷|bSI�{�#�C���b2T���i�,v\E�w����^��}�5�ڹ2����j��n:�U�	{	����)L�]�	��O��5B	�*��v<������{q���I,q�����P��-?5ҳ=�z�[}�o�T��R�?ȃw|�ʳ	��1��<�{o�|��j�[����4��H�Ć��יE������`KM����vb�^&ў��#*A4N�q���5�.K׉��ķ^a����9d,�|s�gy�V�¤�B����{I��*w�%��G��Uܺ���!幸��d�&ep)�O�������}&&���_�K`�'#-�R7C����� �o�>�M��N��\�o���c�
�]}q�����2�z
��@��b�Z����[Y3�r�(��'�c��_�=��v[�-��ks�uz��$4���g����i��aF�6�G؇@���%�65k� �ݪ��2�L.�R�8Ґ�Ű�����#wF�o#k�HC�Me a���8�%��yBn�i�#�:�>�N*��~c"{�Yx���R�hC_��N
Od�����8Z�+iK�i5�Ͷ�<��CCS$���0�6�3�}\O�������ZᓯTD4GX�Q;)P���ǯ=�b�� ��i�ꅊ~l�Y.�?�m#��Md�N��	���X�{�0Dh`��o��9���I�S-������B|��߇W:G����6a���>߶�P��DكOU{Ω6�7?�G�bޏ���u&z�Y�е�>�>����e�|�+��Ӭ�
B�Z(���1�=x�C�| 2i��S �	Ґ�R�?��!�e_��1�^`�-�If0�@V5�Dd[nu���  �	�[��o���ui������ea����Xo���06� ��Xv�(���c��u�䳭l�\Wq:A.]S��Ξ��IJ�D��q)�j����8�.	��6	_=���I9V���n�s<ZZf���)rɕ�yZ(҃K�����G�ʦ�|0�d�+�,�{�kѐ`����´z��$��ݬu�K�m�^X�5�b�����E?��s�l������:��}�˳v9M�6��W�%
�p�%?F/⽆�I�ӝS(j|��8�,&��"z�N^�I����y^��t|3:-�w��᧲��&9	I&w+\��U"O��2�RS>�8�t��s�������Ѕ8�'+��I�X��ٛ��ڰh�瀍�&5��`�%�����ǭ�
yT6~��{�{�ܳd����Ί@٘���`4%��s��s�9�r�]��5˻=G��SvF������	U��9�&�)L�y��E)�kM����+�Q#�'*L]p�m��3�E�)�p��h�� N��.���y�]5Z���S-����Y��ҍ��S܀��`�%-�v�O�r�Le\��4��|��5֖z�����e���)�2��A&�A�SK; *&~�9pb�O.�	i����aS���|�Rpނx�W=�W�`M!>Ꭓ��v_�~-n�xvcV����Q���>���6O���qv�A�yU]1�c��z��5F��J���2���*�:�Du���I�j)���Փ��l� x����΋��Q*^���$,o���?r���w���� ��8a�{^J��gV�n�,^`:C��?��垒mp.�z�fA��Ţe�Lmwd��Cg���+����p�d�>�T�_�l�zS�+H�V���f�!O��H8V�z����Li�qjیh��QɁ���V�#E�:����i���K�7���嫴]�$o�nn�ۡgK��
Sy��&���	���Ivp;W8w���k����	���J��$ĊN��ClO"d��,�D�X��d���آ"(m��ķʗ
uf�{��-�ˋN����F�g�^�^2_�#��-c��Q!b�LBW��)�U�hx�Z�p�:� �:��z�5��G�US��~\T��zqU�p��4�1<���3�����6��9�G����S�W�lw�v�m��WϮ�F�<��kX�R1�-�?g�u�����qV�⺓�AV���V�^�ټ���Y�ȇWH���&�>$����d,y��� j���{ii||Ip ���;��� ��&ю��`s�m�Jk&Ս�7y~��X��njWYB�f�Y辀�Ցlܣ_��o����9�0�d����)���or��/Sk��\K�[ٱ���kPaʔ ���6�('�e�./D-vj<e�g<'��e˂�d�A2��s�̺��a���P������8�MTܐ4��#؞'x9��'�5F�jJ��b?�t�Cs�G�dK�Ehj�N�$��w娝�*��K.�,����BE����@���N6,M���d̪�T��/�V�����1�?��$wx+SA ǅ�p|�X���1j��&����g
�	����a���t�tq��+�S,�/mF���$_�AEE[�3����	[������-���G�ln�y���7%�B���B�{�W�=�Z����INy��t��	�4�/�|2SEA�6���&D� a8�����Mml�u�?�B!�p�7m�fr�JR�r�zn�_;cp��|����}�ǧ�a'��mf�u����犐���D+�f!7í���NB'S!`0(sØ��R��!ߎE|d"��cI�d�������]7>?ym�]H^�}R�
D��8���@��Y�P]����g�DǢT>�����g�+E���+R�t�ӄ*�+|�e�k@�M�8��2��2�K��sera�(� �0�W\����:3p�ΕG�h�1�B	��Ra�J1��]Mzt���,g��Q���ᜦq���b�΢G�.��!����-���=!A�ĆD�9�蜒�y-Z��1MB����Rg�76<9��3�-ɓC$�):}o<�y�M�N�)��n_�D������Q��)������(�;�����C��*��'��0ٽjFZ�t�b �_y��5�\����O���,�m�&SF�?�q,eȸ4��-��>�&5�D�>�������J�+,_�@sz?��1B�_f����ޭVې����^�Z��^���jJĈ�.[7n������oS�1ؽ��3ӚBn̴���8��M�`ۤ�׹R����2� ��բ�E�p�l�r�.:�A+���Z�P�<�f�Om�4K�*�K��'
��Ҙ�5���.kl��V�����x�b`,_�K&�K�f��l~�S�qa�������h�(��0%��"f��Z��l�x�V�츭��|����*�>3IhK�h�*�)P�Q���̅����d'5\����=V����G���N���Z>TB���|�9$���s	�#.��'z���3�ɽ�-��p{���[,�.sVq�W3@�*�1X>�f�%�g~
 e���Lba�b�}a�v��o&PO���02g�ѩ������"���J��اL�ǐ�v�9< �k�׶/%��!UȭZp����M�B��n�pr�/�5���C����P��-�g���#/��s7��d@��{�K�A��p�FP�X�Dzh�Bld ӧ;H�I�g�X#��*\�L�v�Cƪҕ4��HMRL��"��[ȳ�U��"e%��8N��ʒP�vΎ?-���Fl>]��@�5�=���>���Sa��dg+4M\����<�E��}eY���mZ��<3�u���(�܍/X�y�,/��gxm6Ϯ�:x��:�!�k�� h/x0��F�6Y)`�kw��lL�#�5�r:���ˤ�* pe��?����y�7>ݝ�Bv<��^�`m@4���Ŀچ��Mp�V;Q9Լ:���oX��wE��I� o�q)C��4T���Jy�5`t�S���<,v��w��=g|���tP/�l��
���E��葧@N���$J�ۡ�����@�G_ض���?��\CX�}�D��W��zS����B�K��w4�mI��O��Y�+j��]%��2z�z&�0�ZRN}�W�E���I�T�� A�c�[NI2��X⬠�1 �q|��M'�I�����@G ,���]���h��O`���H
�4�Ǌ�t�FmD[�4;�n\x�?��V~`�ȟ�S~�0��}*��Q�N�I�[IX��!4�S���0��n8�\a)0+�������<#x�x��4#�E
�'���|^��i�d��h�W��1*;�n_M�߭�릜�8ބ��巰;�����P�G'���v��5����<����sў��@�$Tc�pV�<��ڏp�bWSCx��_}_0����Q<���^���~V^�>�ⵤ�o���j%�~��$�!C%#��(��l����s�[5�[�y��-IA�J(Ů3�{xw�ָ_��y�ڴʡ]iW1��eʪsw���0&���c�q<NI���E������-�7�|y#o����z/iM��U��K<Η�Q�b�v��+��q�=ݾF��#����n%J�b���fS�Ǧfr�p���;����ޝ�(&L�n:�^)�ѕ�t��-z �])EԤ݄�\�lE�bÀ)�[*�>�����p��VZ�|D�A2�)��.�LA���0q��j�\�n��<C��_` ��⼥E ���P.`��; �Õ���'Һ+6bxi44}$�6�#9G�1j�j����`��r8�2l������܍X}�D���E�J�c(�C:>ch́c�Iz(\�h^�e�V�Y�"��	�W�N�^'�☺i�U�l6�(a���>�ƹ��)Ka�A	���$����Ǔ��k��c,����J��ظղ����}��#��%����CR��S�';���auNO����"wg�� X @���!��D�Ǭ�-f�.Cf��rڊ$$����g�SL�;I���ŽE 2�N�V`*��9�pWp�E2���<�����xһD��`ct�x�y<?Tp���c��3�0����z�b��/˘ˢ�AG|�:���>5�ܝ^-1*��K�x�5$@�P>Dt���5���z�k�@6��`�6݄M���������B5)�����&�N��>W���Ax���]���2�Fx*�1���HOX=G$i�ǎH?��~5ܕu�Mpz�����e�<��U��
�7������������aV�ǌrԱ��������[Sd"��0)���W���	d�k�Q�x���p6ɝYP)Sx�� ��X��Ի�*���e��o�Js^�F��T�w����U���rr�#o;���̿��I���d��R�������S*�5�է�|%@0,��yKZ�갅�������6�z]�Y�[��]�SӲ�y�H���J2Le�331���	g��b(V�N��q�m�_���s�=G�MU`����St\��a��*�ކ_a`"�U���H����I�P>�ئ��9j�;;���ލWV+���H�d�2ꆛ��3lm�X³#���l����ޠZД	�����x<��Y���#��߶�ȡD{���D؋�e�A-.�S��yÛF8�lU[��Q���� ,(�T7���|���]�C��;ʔ���c����n8�5�������\�{�V�E�P��A�D��\�CK�մ���gr	è�EAc�>�a�_[�����ˤ�߶��޵g�̘�j����怆��95.� ^~�v>$�+J\�L��ۛ3E�s��� ��nP�C��>���By��#�Y��k�
�����UAĳ��Q!q�:��[�cؿD#�1�)ݵ��`FBbĩ����wP�+L��ku���nޔ�Y�D=��9dy��8��7$���
Y����'d�~]���+G|$��F�B�r��R�W�i��]�P��y|��'���+���� W��%�tG�L��{/Z<ѝٰ{P.��zw<Y��9����y{K�gaP���!��K��%
p�@	��ŀ�0o�|���@��:���B��hl�����O��0���R���>#[�8�Z�w�'q����w�?�ݘ���;(t@��v���H�+��G�]��3Yǔ���0�ɷ}kGg����<��ĵ2hWr0����_��c7�c+�a�V{�+�z�I�����q8fӦ���8����²&&Į�t7������J�ߵ�������1��:�>^-���7FX�KBҳ�!!��HLh���{C-O�=���<��nE����$D�Y�����T�&y�h9w���.��0��"K�2�ތ���J�TDB���֯H���stkF��^��o\�����w�2F�+s���ѧby?��P�x^{I��`���˔�~S�ޯ�ɤ��̔�P@v��\�?,Ď%Mk�'p
H���%�Q)�m�xWhT:_�z��h�"��e*8�~��s��׾
���>��?�Ø�wz����A����E� mF@��썒�0I��9�~����H.�o�/���@�#i�~�M�4��P���	m�������BE{k]��/��ԑ��-%-	�ЈXV|~��ۥٜ�4{w�~J�ݸ�T�dd�A�O��M�q��Ąg�:���ѽ���-�+4Z�߶^�C�,������~m�l�s=WHo��D�D�`�ۅ@��pX˘�!���[�7fU�d�2���7j�f���k��.8�8��1�%��q�gk��1�C /Q��~��v�0m��Z�V�W�@e�vG��?��?�Ϸj�Z�"Zֺ�j3�ܼ�|�M3����IE��x��P�]�Dq�o���G�@�����.@���a��co���ER�����)$�����"�|ŵ�O���#៟˗�����ɝ�!��������E+	y*��^�@�������7�����*#������4}_�����	�����'��s�q��o�,�aP~Y.$"�)b*�|hT�|��U�V�������#)>���:�oۅ��0�����$��u����#j����~��QK�#SOMj��<(%~�ק��J��Υ�y�¸�ǎ��˙�БP�*�����]���+o���CM'�̎e�9�"�潊X��4�tP�"{1�^&���2��l/zTT���)�)����:�0)FUD{��R�>�#z}��(U�^��	q�8vH��j%���.��0��_��]G�H��J��-3'P��f<`��� N�٩�9�]��8��S�]g!���,M{���Ҏ��Q��+�/������҉_3���m}�)�Ri4��K���p\5q�x}I$ϣ1_�A�0uC�ڭ�^=M0rR���b.al���J˨��(�l��6ň��[���;Vk����Nn���B��G�_�� �ɑ��׊�L�ҥ$�n��M����y�>>R^D��"��8"0�H�=����-�ǂ�OHy��W� !.��h�1�x5Hх0��O��z�J|D�P�0�gz�alʢ6�<dvW(��m.g����������;���!��n~�ۇ.|CX�!�K�_�� ��)&��g?��a�5,'�D�y/z�3z����-^t䓾t��_E��zL�� ��_owCe�<��+��-�A}[T���V-�,g0�s�<�����P�kWQ��*�����ޛ��,���HvZ�9����_��( )�.y0�4�<�QU��xJN�	!F6�U��&z���>�,�z������
�T��U����A��ፂW:ؽI��*���i��P�Oy-*�y����\%M���NJ�ޭ؃y����}5$ﳄ���;S5Nh��H+�XE ���Nu6d1�A����}�v!�u�S�XlT�x0�;8� ��J���]�p�M�P�l��x�#X�qiJF��|bֹ�-�hP������.;% ���ݞa��;����-*h$��w������L8����GrZN�d��ƮG
)���A�������NX!!n�,|}����>q�XM��Q��Ui�����K�e4�Ó+P�`��A$�p�В�=%����]T$�gͼN����hq���y�M�e��m+����Cr��X�h�������K��̋
�\��,˿h�vz���*C��7�0˞I�C�a���L+$%���0Ht���\R���k_*�8�Ȳ팤>����|f����j�1i^�L�g+;���j�~�ԫ�q��H}���/Iy���E���eb���*��\Բ5����ߢ�����yv�?���s�	|�h`�֧<���icu����|�M��9dϻ;�ݱ�J֙`�f;HH)����z�.���ڧvN�֧"�F��bYNJ~C�ޢ��� ��n[��W�i�5�db[��7��x�)1�;HY�W��&�N��8?.�X�տ&�xr�;|W5^�k�Y��p%�!E�hmR��y�%�ɂ�+qb�����/�ɝ�@ޞ�OW,��PH�Eٳ���Y<�L����+�j7��D�I�Y^d�Km�74-wh��{�C��"����9}F0f�C�_��9�:M����_���3�v�\{�v4�[�Y�"��u<���?E(���gZ�'W��8�cz�K���|}lFɖ��Bk���K�^��u���2l�3����?�r޹aOh���+e��Z$��	E���{��v��m��s�bn�PR4ۛ�@"����J5�9I̋ӾG�p�%`�"���m�^�2�����i���4wIF�� X*��T��6�D���`6#� �9Ըc�z��֣��6ޢ,��Eh����2��N�#���e��ub�2��[�k�ׯMf@
9�k_��b_�wp����������"O ���<��R�t�@�U�ԁٔfvf��x����%iۙ8/�+�څ�M��#+{/�n&&��&��ؓ!�%O���&#x˥{���(�$���6���0ޛ�9>��4=ɥ2��[�Y��z)�N!�`{�ؗ�.�O]dU��|j�'�@��.���9c�c�k�V�����2ĭ�O1��7FK�D��\��5Ԑ����`�G#��xhf/��4�0��G}�j<rO�9f0�j3k����o�Ш�IQ��a��-X<�?�o�m�7�?�,z�����v�b	���`2u�oڿ+������3p��7~:��ő�L���9*� Y%��sXR@�<z=��Ю0�Z��0_��l̏���=$(��(��KW.wv<�3�6�j%$�r/�L��\��ח����!�N����`.EC�RƠ �@`r��A|.J7�s���ppd�rgz��"ހ�3MW9��?�l,� ��yM9�#��H���"�*�L��]֩��Db���rG���u&?x��&'�s`��������C�h��a5ڰn�H�FD��ҳ�a�8�06�Zk���+��A�Nx�W�������bL�MhQ ���*#Ev2r��9�N�f���Ԯ�Z?���4�
ڑ�)ܽÈ� TBu���o;�/�y0t	�|ǮkH�����K�t�wƺ�i�M�%\�`��H�U��E�з �+�+�y���[k�㮺�M��=;{��)��}���&HՐ @W���ّ��R��:�� v@G�~��M�U(EqmJ���d� pGJ���bAh_�kogU�	�`8�3�e����`�۹$���C�-�����}��Ux���x�͟v�U;��uA&m�|�e ����x>�-i҃s���7��^%$�?�O�$J�<+K�f]!��Y��x��(I�%wT6�7��8mܹ;�y�� �8�;��6c����
��,9�E��!��n��jǎ̏B�j&iE����ξ��K��(@�E�f�-Q"BYxҜ/����F��=
���_>�Nڲ0����s�蜷�Qb�@4�s��y�ƋM����rNq4S�H	��ျ��@��F�׿�+�('d� �E�L��A�E�'�	��Ǜ�$o�D� �{'��������ֻ�4�dc8ư��� �w�� o�@Vg����i�> ϸ�,7"zw�x-,�CtӶ�"L+��/*�M"	Ҷ��[�㜗7�d�o����p�-b���>R=�*�t����k��K"��pR���cnGRmנ��a���/!:D�ah���f���S\�uZ�!��qM>����-�3\�/z����	��դ����kzQY���I��-�w�2��$���Bq3�Ho��/�=���e��%��zt�W�Wq��NӸ# ��u���|\f8��[Ց�fdέ��EugX|�o��=�_\H>��j��4��cI��,�]�$�~�2�����@M���HȮ��5~��Bj�Cm$�M���f�Z�s�K��f��I/�*��]ք,p�q���$�Zg��:��'b:�&���l>W�-�q���ļU���q��xjKw�2{v����ɱ�Pٻ	*��Ff'1T�4Q$n�DnU�s���z���s��������C!�S��׳����=���(���U�Q�M+HG�U9�2<�s/�]�������u���x �!�K=��h�֟��UG�\c^��;����/덕M/4�\��ek�s|�WR���1�?,,�YsU�w���Ju�&�Gy�i���!���m��hgb�~�.}-ނe͈���ۨ���=n�KNT���%��ċ*w?O>)�A��`':E��_Y/�?�y���&��=�Y;��:��uJH��Z&���W/�l���j৽y;j�}vNl���w@R=� L>j.�[ϧ���BP�M�(���bS����DN�����Q>#�6�����i�6���.u��6�gX�R�y�KL_Q�O?�L�V.a� �&����48���*�����c<A�;�[B��gJ�)�'���<b��2{�rY~9�W'�YU3��)�2�F��d����mT���"��-j:��	_ �7��#�΅�%����8h�ڥ��R���P��X/�m��Rf+�X�|��O�s��<�?��dp0�
�WėV_�
�.F���6X]´�bi�º��I���p����A�H�Ļk]����J!�谒��[c��Ͽ+��#ƵBu�2[�n�̔'��D/���,�e�:��\��/�����wi�cmWV�X�������n��:_��ɉ�/�^����A��q{�\���^D}Z��D�8�G�����RY!Z�!	t���:���9�N��t�2;���������(%���"�����qu�zn/�[�3�ݡ��: �d�ؗYP}��B>I7�fSz
�G+m��I��`I�OQ�pS�Nq	m!1����P�����I�Z�n����"*�fL��z,ں)��c�
/,��rDΕ��<XA�Ք6�6FZA��2_[S���c�@��~5��f����j�˹	R�K!�ڜ�D����D�e�8�Mz0���=���.���
#��2P0�l� �	��E	>��Ώ���~P=O�J1��̸!zK`^��֖����
�mrd8eF�eD�.��47�#���+�)o�r����{�D>w�I��8�����X�p�V���&W#yF;�A	Nڈ�������L��Q�L�_5��Qx��דW�Í7���P��4��գ�^���uT����K�Z�=*T��\L�ۤUE���:���o�\��ҩB3>��Ipp��D�a���:]p$���KO? 6�[��A�u���ϫ��7T6)92SMű��&�u`����Ǐ�*�[�D�PH���_|M���<��ԏ��g�E9�S��u��A������|mP��f��qƅb�s֘p`��l8��}�%�A�]_�}��0$�w66�˫���n�s d+"�BP��^�_j}���lyM[@<��&%�
B��	g�pa,8��F�+O�`VN��d�k(�=��`F������b�N�*�0�ۇ�\Uu"�j4���ʋA�[�����Xgd��[�ȿ�����4����>��5-;�_����0�� ����Mњ6�y
��!
�d,[�H�V��Qi�ȩ񊠎��A�ddu�	e���o��F�uz=eP�ͻ�Y�����{ŉ8��w�U"�Ҵ�PW=D{�O�&��4�.=@v&*��Q�]�<��!�\�e�O��#MXD�p0�q<�ω{�d0���Kzg076�H?~�e$pw�q���3�Q\��%y|�h�OC�6�*��ܟpt�J��K��J���\�L���׎e�~�����L'u�!B���k�="��zSG+�fY��@�b���j����Cv��̿_�gS��I;^&� u��}��D@��a�����;���"!�b"QA���	)�G��$�����^:Nׯ��ϣ�:7x1Dl/}�#�ffx��Í~������$�{' ��'/������3���b'E<Gy���ʏ��qڥbV�M��y��ӝ��Gz���̫̿��{���)�{^nc H���.��愬l觐E��O��Z+ce]���P�h���p8��H��Q�#|�RX� ���^��nKN�4q����k���K�n����(E�ޖ�l�[��D$A�����
��gH�����neJ�96d���v��2�ߕ�%�-a`�`7��T`<h�Ĉ�N��h��9(�Ya�&t0��2@D4@��d�����5*�����!�8�����B K���q�9'���25�
j���{�@��eJ�[۩\ P~��@�}�����:^���T�Nи���4H��?������/����F�q�ɂ��J���Z�e�Vt��;�J�I����Y!��#�}�0��@��x�ƈ��2 ���3��I�Vkt�(Ȁ���n��XB�֒��@W�5z�%j��ii� �LMdӗnU# F(�	 �K��U �׵=��wa]�Qf$��)E�Z�����p\���X��R��0���$+���T'���F��uTG˞���|?�L"�K9�N=8��y@U?�b��H3PJE�|�@�'���3պ�Qu�Gׄ���]e�u�5[dtG��Kr <D�c��~������>���H���MdG(Y9��-�T����}<5�<#���`�PL�G�v�#�oj������u���(��oG"D��5*��2AR���eE�0���gΑZ�Ud5����Y(R�mo��p�c�<h��x��30��d�x�U���J�DDiX
7l;a뛻����h��3h/$�V$1�\�[�E��5GOi���]! �eO�O���~�����㘁��+'x�o|����g-�4�ӋB8��K������^)5&���[�������c��>�4l�Tk�F�������N]!ϣ�[��!!ea���8p�y��lfZX�a���0��>�|�M`�9�z`옖Ri��|��'�D�2Ǳ�ߺm���4�<���� ��,�=����\�Ɓ�����	��"W��3�`�vz��ijo�~-_��`�wUE��i ����j?<�A(X�%|Կ1���+t�K�Il63�����g������f]��G�����Sיִ5�vܟ���?!YՕ�q���,J*A/xX��b�X�lVr�} -8��Su<f/"���v;�g?�*������4�6�\��ڝeED��Vl����e��Q��m�Y3��LI=۲/74�!���-tv_E��䇤'a�d�Z*�Q2�j�0��\��R��k�� b����'��yK�E-�k���|9��?�F��/+�Y������u��$rk����Q�,��5,�*�Oǧ/����R���T�4_�9,u\�V<�����}������0	P��Q��-��J��pyJa4N���;ۏ�������$����Pg����ȳ��0����C�r\��;�H詙�|���Qt��k����X{��<�H����k�+�Qp'��˼����.�f4�� �:��~��:�n=�un� h�*��2�k$	�h�z����x��e�I#����|�j������dkMh�˘?��>"�)��@���T&�D�����#Q`��5���E�@Y��x�r�R�����{��l5��nVJ��<1���w(��|�ʌ
�O3wGn�i{�И���Q� -��� /?ӾҪ��?���y&x}�Tq���&xH�;�4�4B�p��ujt�����?B��;0K�ť$'�0��jE~�S?���d �)}�P�<��с�Hh��4�mt�5W=�)*�t�z�HJZ��ă	]�>Ζ#��r�����u[g��.�AB�O�gz&ثz��A�D�g0�r��0�5�+��~����p�zI1=y���yK#Ȋ�.�)�9��
H���:޳?��!A.��C��9J���<������-��RH"�N��s�*��FߐA��kO�ؓ'���F�����q�5}{�v�/�$��t��H���L�OM=M����'%?�$ӄ�66���,����bJ�*F?J�aF�ޣ�BP�h/�
B�O�\ځ]��=�]�ء���a��H�7����0�u�4�]����ٝ�H��s%&C�_����ݹK�7����]�����qG>�9�]	թK�'kM��s�wCZ�����_�tG�7h��W�IQ�0�1ٶnP0���h����1�o��6*��d���v�lP��H�;#�w��L��j��,m���B���AK�N�C�4Y��n/�Z��2��y��Ig9�K2A�^�ѕ����g"ʮm�%|��S����G�C�;��+�X��.�j�0�S��67�ʴNFD��asW��y!OxM�I�j���l��lഡC�qxq��g}.8ֈj�\��D�idv��V�w^�������E��~����7��r�.2kvY��v�<�$���w��N�XB�x-��^F~��Ԩ���tJ�+�m�o!+�&��o�]Ə�0��a�6Ȳ����sǧ[��ٷY�+^� }h�]Y��E��;�����7:�� �m��6��ùࢷ̨�����I*����*g� Ť�@>���������U��g�Aޭ�}��T�(�j��2�T�uc�l�:�Vg�"Лe�h֢��X�o/�k�b�{s�=9Ġ �x-���22��x�f[B>�N��o��;9�۷���݋L>v���p�6�/;;�2�� �'�}Zj�]��N��k�������~8�Y���K�Q���s%�1aj�����d�����2�K��w����8?�ɓA{r�&����^�D�I�kֲlx���9��ohsR���yE�Д�����i]`�g|#y���~c�T�g�0�IǪ-)Mi)#͚��v�v���9�i�'��L۞R��mqSh�h�v9�¨�����!�Wi�k�����ʎ�!��^MH�-�W�B�$V������eೊƼ}y5O���:xi�����!|��~�B1�v��|�����\;ܘ�+�`�2-v��ss
�y4
~��jc(W.�\3ط��櫫���lV���eA��F-��f�D�NK�k�7�>�T�F�ۘ��ƻ��1�,a��fo���_Z����~��3Q��	+�F�;,��c:��H$�17�S�H�ڙ�$�t��4} ���jy*� k�ޫVie��z��j��$���"�*����x_�@k�s=V��2il�k#� GZ�w	ˈ�m���6\Q
t#���v�0Y¥f��s��Ƙ�����i��.�X�$߾L��#��s8�^�S��
1��)#2;ed��"L:y�����{Rc[]�Á������U��L��z�k,�ꮷ���
�|l�����Ow{a�-��5�*&�L/	��V��6"�ED��.�kk�f����T6�CV\>Q�k�����!Ԓ���DiU��g�`-T���SH�iC1�6g983W�VL�X03$\�l �/���XΩ5���U�� c�+RDm i�װ����LO�Ni@T�t�.<���Xo�m�b1��sh�͞�{��[�7=&)�|�W�4��\���H3�	eK,��5�c'(�E���%D��~i���Bl�y���N����`H��.(�b�DL�g��M�
��� �h7$��1�$q���6��]��R����3Q��J��kV_`2
IZ1�v�a7�������r�وW1��c�G�:=��Ϳ��Q���R����(D���g%Q�S��7� *,��0e<�P0-38��>P��Ml�w�Qηh�Hx�����(d1I[f�&g��={����$�(Z��/Лs��i]��~p����&G+�,!~��@'u�ClGj1��.�^ ��Ѻ%��ѵǺ��!r:&�E�}�Z��+��"��B�r���ra�l��py��x?b'i.j��Pp��e�\�a�7�	*ztk����.}�v���k���%{q�sN_E�t�J*��nh2b��;<b�s͠��[�q��������;@!MB�I�O:�a �w�~Jc(�q�oA?�O����M���a%<��C�1�*�^�Y�}��� >��7�  �����To+���f~*WT�N2@5�5����u���M���V4M�
�SJɩ�;$�8՟{qJ[D�N�Y
7[k�k[�h��ɥ
��8���n2����z��Ib��?�5Ϫї��t�F
�Z�F}3+��uل����f�Pm�91-�(�M���O��0 �.��[�	(J`b�a�7~c<��g`���Nt+Z���x���ܘ��|�@�i����
U� �k Kvb�����s@S,eCDGf�,;��c=Ns��N����݋#��IX.��:�>����<D:%H:S5f�d�A�C����:5e&l8XC�cPJ�*���4�PZM��8��Z+l~����q��?��	*��
_T�o?<�Z=�����5G��rm���|��3�A����|�2љ�3�8n��|q��n�M<*���'�ZF[�׺Pg��1J�R�T$x�$�I�� ��	t�
q����D�\ě��e�x(n�o�2�FP;@FU?x�<|��9�W,5^�U!�,�2�;��2N���^A�����}�����ӁZ��'����+�;[���F�P����i��i#�ʚ��à}eI����#_�ǫ�utc�0uj�k�8q��쁇��#0��|F�QC�-�Vd�"��j<\�fl�^6+�s���>�&X�}5�m#!�rs���׌x�+3�K�3
LH�	��A���p��<$�%�_��.P�����>Ɲ��9�XJ�'��M(�Xpem;�0�Z�����f��T"ǋ ��Dz�g�W.1�O����;2��ܤ�_d��UB��yi���B�&�$�5@�Gg5aM�n��C�
G�$�)ח��;@,�/L���|��s�"R�k�^�0�¨U��_�ؐ]s������6)�(+���y�s�(9X��fF7��cJ�xn`U) �B���k�)`��b�-M/�/�PQt�����8B��jLX���,c�pPɨ��1���	��8�Ñ��\	E����B�̄��)�(��c�gqg�k� ?�4w��#�(pk�k�����,�����hCt�릲j��H��<��٧͆������i�/�����M<��3Q-KbN�
���sۈ����y%�����͹�^$�_�c&�_�f� N��Jpu���o�]�2􃣅���d�5f>� ���z$��>�>�&8��Z���\��H
��x�S��?�(P�H��S�H�t�v(q�R�r���5���@X:���&ڄ�����?�~M�i�p�P
�"	��.R��4��HX@��C�>�~�ȶm5����/qi}h��yG�@��?�k��43��%��;���X�����ζy��H~����g�f貅L�ˁ�`�	������>����Vi�4�����M����)Ҙ3O<Uq�|�s
4�r�J�M8�*z�P�V���&9g�v�P�q��������z/�L>����)vR�H�;E�����钃���4X�	 Pѿ��8k�������#�"�G�Y�9x�Wk)@�m�1��1H6�b�*9���"�"�"b7`����W�5_��A��3��ݦ����h���:!0��X���$��Q˪�j:��Qs���ɜYA�{a[K���� �� �(^�z���:��\X��W�]�Tw�N����}�8�T<��7ߢ|E���{�ޠjF�}P����j�"v��U_C#�	�?������-�������hX���>�U)6��S�sh@?����fA�/F�� 	8�B��\5d�t���No���dM�������=�S@u+��P��OCU�#���y���s�C��H��ʲ�3���wG)��7e������I=���ޯ#!38L}ރ
ަepfw�毡{�edV���иEkHTû�W�9���mA�jS_O�����,z���[�w�5s�����l�9ZxT39����@5gd�RL������d�p���65�˻Q��y�f:Qݠ�6�"��y�@+��Xi�Pr
j`��Vܷɹ�ɲ��m�'��!�=�f��\TVXV�aw��N�i���-�\L}���n}kq���Zo�>���g�zָ;g��--|��V�몋��o��*J4xq���x�s�O�������:�fv���+�B����X�R�6�F@�K����V���nq$ƟV�o���T���P�	��Ě���H���<�>��if6�ƅ1|2��:�LV�r���'��?2"��UiԪG�$��ۀ#;��X#��M9�à�uB��䣾�u�Z��ʤ��4[o���ENU�_������������3������^�+w�����}�Min�1Q2�� �#��H0G�L�LlV �5����gb^<r�P�x��Gl���Q���N��p��[R6|
��/����=F�C�G_���9�+X-���4^�=��I�n�F��;$�M���%�)C�5@���>K���J���x~��$_���s� �c��=�G���Е�L ���ft��bR��D��\_�T�H�A��2���cY��P��k�1�}&��/r׸#�]��,�"yT�'A��y�,���~@�۲T��/�b?^�s��
�.�c���H���pM��e���f��ic&`rT��a!��q����CTi�t�F(W�!^���ti���}�W2��~�9���U7|�3|�*�ґ���?��r��?.*���)�(�1�������k1��
��&�a��mh�����eNL�(��p�A	o�$;�=��B�¹���4�%GI} �$ռ�R�xaZ�\̽�����c�S��8&�@LI@���&����(�|�+�����dvw	(Y�Yx���e1Ba y
��!��6e�V2������Ε4?-��yYe5��ݐ)V�+�2�G�XH|���A:F���00�������kM�ű2�Wͱ'W�\#�>���:u1e-u��
Ӭ�����b�.�]�0�ܞP��2?]�P�j��"js,Z�F=�\E�"r�Z&�Yb�x�QV3�l��嚫8��V���c�UQGK� Ed2�Ö>S�ru �?g���'3�7:��rUï������ȗ_0���!9p���ܡ�YS�2^���)���? +t�ﻎ��i�Rȶ�r����Y<g�����`R?5!S�q��+�L���,����-0�G���DO���7W~�0YoFJ�:
R�;�r6T�h��h���{]��~ r��K������ͶR�z�_�O��|��Lg��98P����׃�]��+�����06�6����X����.S�BXX:�j�;E;^�e�M�9���UX�@�8�^zoh�<����Kru�p��
�&��]{&o�I�`X���e�iY��J���Ա�и�S`z��� �����p���<R�q	��ի{���������R��i�5����g���)��5\3K����?�"M��0�+\�8����i�+Kw�~�����x�e#T��;�j�d/7�fZ�U>�2n�S��h��'����r����=��̭���BgYb���#>4Z�\���S��V�Y�����O6$g7��&��)�`o*�}G"�	>	,ݦW�D}Z\��GF��#e���~���/���O) ?��( ���V�a�X��W�t*:N�VU�p�����;=�kv.�Y�fg��>K�V�Fbm}�e�]�TN���SptNn!�g�x����L/FL@]�f���ͷ� =֠�?-n���=!�ېg���o��2�V'R��w>s �B�����`�د�5-�-5s�"B�'&��灙
e�琧����230q����ֆw5}t��D55oĂ$�����̲�o�W���&6���[��_y�F9,���Doe|��A���?`ty� zq��C2����Lf�����i%��@3�l��[�F2f����\�/)L1��%�0Ls[�a^��;S��h���9�k�,�A�o��t�K]a��y���L&��,�wi�i,_9[�E�%z!5$�L*l�o?���|D���M�c���h�8�~�E���wN�eE2U�}):��)2j~����4��m����ti��g_6�=�V��?�]KyK�E�^aR�Q3���X��'��?X��B:�.ۺp1bepP��Rq(ۑ��l��i �\�]PŇ"V�7Nܙ̒P�E�2����Nީ�x�JY�������/�~��j-6�w��&l1:�� u��G[�I ����)��Ur���`����s�߭��W�ۣOQ7�a�M)�+������ߴ-�K���&ö�'� ^����#��/���56�nJ�\.A_k#�2Og����P��.�q���=)��;H�p=x��T"m�Ga�[��!Q�&Wvg&;i����u�D�]9(������h�v��N񎣄�:�b��XOW<�S<�����}(���ҳ������`�\3| [i�ǧ	���&��J&�A$�8�a�n��۷x�i�A�:r�V�;H����Pc(9�P�ntֻ�ź�+V��]��](�GD,T�x�����SvX?����+����*z	FVI�l`7��TA_��%��y�:R�F�����5�b�	s���;�&i�{K���'k���,2������J�)�!����V[�3y�F5s�9�u`wr]d}��4�rC,���<�b�~�Zy;���^�e)�ғ�0={��(�����{=f;JSu�t�O$}�9��i�o����U �D	�qΡQ4w)��:��4.��N����m�*�/�SKn����U[S���/�,���m�[
w���"��̆`|ϥDe˴_������y�5������(ǹ��Y����1Và+��A��?�)�\��R*���t�[��1 ��~m�h -�.i'ǭ�W���*��I;��f�F]<Sm\����&�P�Ř�+ކ���&��^m*�C�A�Sɧ��
�K����I�u�_a������7�s�{B��J�� �Zf��6nea���ie@���^gX �u91xϖ43�Օ}��C�bv%�����ń��z�6��ڸfɘ$��t3Z7OSsd�fQ<t`ɟ����K=mP|�ɤ��\S�1���L�������]{�[#Lj�K�7����I����{����~�O�m�c��氢�>��)��%�$d�i�� )p�+��b�|������\�䇔��k+���0?)�2/=�R���4'�M���]l&'}�����e�1��=�үc�԰>,G,ʹh���f��a���8����xk�{��KjL�k�A�y���&�wPʵ
�T5#;��̝�g�����F�SH�����-��ո�s?�a{*��{6�@k4�;��X���W-C���1�����{�_G>�q�A<
�;;��V��L+#�Q���m�D�3�SY�3lٱ�����4�ݯ�`	gS�Ʈ��g�+��^�s[\�!��q�2z.Ŀ"���t��RS�;N��:2���j�b!��_W)K�$�$~ԡZ�}69���}�Z�c	5}���T�N�'�V���
S�l��ǉ��B�҃,p��߁թ��i��JA��g�dȠ�.�p�y��H���y�=�o����Ě[hܡ0�s���x��&�������N�q̉d*,V�^H=J]�)����5��{�.��M����W�;4��(�	�N�@r�*�������l� .�\�O�����4���N�� =��{���>�?�K��Z�s���.��΂"|4(�rǟ��=D,�"����K>���v	''d�d��e}>��Y�p����M=6��0*�(��/���g}�Um4`���.��P��5<(���.�E:��� ���)ëv-j�.�U~$�P6D���V��Gx+t�n���z-h����i�|�,���E���L��߀�5�c�r����������T���W�pٚ�/��ȘFӓR'��%:ݦ����� I�Tw�`ئ;`Ǒt��W>�C�s�¿=0t8D������x#������S�]/�Ҳ៬5_<֠���N؜PޑS�@�M��q<�h�?ڐ��F�D:�ٛ�ɵ��7�?�\26;2�Dq䛺��=b��"�j����?�@�^��֣6�j�d�*I�0�N��w,��Y�f{8�"��w���?,�����)��
�y��\��h�^jk{�����
���?�T�b���n�h*Y�DҌ�j�zU����! ׄ�� Na���������������'h�L�a��ڄ���L�¹9�>f�\�KW���>�]V���eq��eGlӼn���\J�Ҝ=�%�;�b#$gm``z���:���=�z�x	���%N/��
��Sa(`D��~$��B۲�.%�VWہ���p&>�7����-��=D�i	F�Q�Ɨ�=�@( ����W'�k��TVy��Ci���;��z43չ�E��;.��vq�o�<Gy��f���h'��QO4:l:ح���4�n�l��@s���S�d!.�8m���aMQ�u%�c��m�%��xGz�C��F�{y�M�d�;)�8:A���ͯ��DԉZS��EeU���7�,���8��@���WJJ+Ê ��3��oQ�Q6�R<Ѓ
I=��P^)�^wh���t���~��if��I��[m�w���1y��b�I�B� V��.Ȝ'*�����%��[�hM�@:N��-p��,١S�c�h ss��kUpw��hٍv7A�$�:qd�6[�m��u�i�ѹ�	)Ӻ��$Oy:*</D�$��nv�D�,e�nrm��Iw ��J����{� #:���t�<�x2gᘰ��ލs&l�;�S��G��J1�����i�-!w�`UĜ�''ZB$�9��D��ϡ��a�(�@�E��ځr��f��":��,W�Ԏ�(,��#���>�lH����ߧxn���A�c�¢n**Y�֒.�����E�+�oX��k�(�zD��%x��m|�+�<16�<,����x����9���� ��wyK�5�-K�~8����h�G�=�s��Z���ċ����D��n��k�"%N�r��&2|�u^�#]�KqH?�E
�+�1�q�1�n^A[D���RF���K<���[D�/Hq9�#��2����ښ~ڧd�&lX�]Th݉FԳǆ�J��BG�G̃��cMqk�޼�-���$˘gF��[��p3�Z�̌�ݎ?"���D?�.Ѫ���S*�)��_=�E۫�X�pe��l*|IH�?VSB��3�Z�����\? .�a���Z�I��3��"(��ph�n�����R����y�Y�Чo��G}�����h��hnN<��&�,�q�S��o������ǆm|`�C�O$�d���(Ϥ�)�g<�$:��v�Z^���K��b�M����U�N�fv����X��H��{$�Y�6��O�ɤ#��k�]��l�m~�@PNnc*H)�2p졔+�Xa�kjO��T�I�b��A��N�'�RL����q"���RV9�H�z����2�����[T+���W�2�Q�(+x�h������|���|Y�E���7"����]�|F2$>+��_��E�4����y(��si�9ͮFVy��s2ۤK��b�f<�XU�?@������.1]E����i�ܶ�6�
��	��]�*����;+^vaj�;�օ�kՇKs?���UNd9���U1}5 Wz[*`��c}`?["�0I`w�"�|��Bp�H�ȏ_tD���Ow����Q��N��
��[s�h�Fs�S��/y�z���щ���}:�d낙[��ao�L�#�M"�/w����	FO�B��������ꧯ�ԴuթJx��������fK����?����H� <�H$��d�m��ȵv79�A/����g��g�IB�!
�M��}��9����1��1��|U@�rzX<�c��펿 �)��s��!6P*FZ�T��3Nz���U�!���o�{�D��`?����m�DK0|[��ԥRWO����`�u�W���
;Z��޵zj�*�9i5Õ��[0�� �֡��ә�+��~�.��v�t/d��NF;kI�i���q�>6z�ܛ���~�Y�%�dӱP�[����
�����C$`�Υ
�|��#��a�:F+� $_�xP�O� ��{���^U��I)������]#E�-n��$~Y�хOVM�b��g��$����w��!u�6�V��NI��!�#���kQ���.���1��� +_w=WsZst�s,X������%s{�I�At�����z�����IM�����8�*>����J*kq0�qEk�j��ƨ��/)��?��r���ey�Ic\4�����W3�js!�	{ǧ!���Ru��|&�!+��7a<�O)w/� 3|z����Z�^�_?Ǣ
P*�Vwʙ��_���@D18��^p�*D� }�
�g^l�Y���xS�m��Hi ;lHf�P\Q��oQӨ�v<�	+	��T��+��qI���/����L��07�#z@]|�sԄ������!��3��<�	���������|�&ϻ8}�O2�%7�&�ީ��M��Т]f�I�
�n���Q�v�7��;\��EQ�%�J+�/er�z.��������-n��y�~���e���T��~x~��z����2\����G'� JG��}��>���6N1vs)$_C�e�
��6�����պ9~4~�*n���DP��ƍO�-���	͘K�:3-�wj�E�&��y�i�w�枏_�4`�b�CX�V�{�H��n�����Y�����y��Ke]Q�B�-������<�v���� � Qˈ��E�j'}�Z�z�o.�j����ʹ��9��hY����ʣ�=��12R�uf��vJ�Ar���VOh�9[J+������6r��+�q={3n N���J}[}/�s�7��1EɈ��>�[e��#��Ǯ��5]C�;�]]�s�)gO�cJ�k�e�7|�:�Y��u��~pm!�tw��/�t�1���̾ȡܕY%�V�Xum�gI,�}zU�'
��y�>uI���0V�N�Ъfj�%|�ʖ �C�T�Hĕ(�1��w(�:�̲W��Zq]�m+(8�4t�.��{�7���f0B�^A,�2���?[pQ��n�g����8���9���5�;�D��ý��y![��i�DK�y��X���*�`��r��S#�(<������"=H��q5wsu%~�B;¾�;��ABz3��^5�?��*8x��bHК\��vP��`+S�-j�'<�-)Cɯ�>Ͳ���+r|H���'[%�д//1����a�����9��`݊����s9��}��P<�.pm�	y�y�Dײ�#��q�?�O����*�\��Q���6ew�	�-��'�t��7���ú�t��ҫ�HoK:�LǇ�t̔2w�����	����?c�j��Ǜ�ڹ q�=�:-���}ũ"���I㨺qܕt��h���/?M�K����r�Z���1O
V�_Z�pn{eS�ע��Z���ݴ}&���s�BS�oOSt��y�	�e�DF�%V@F�(�>���^ˣ�S�ش���V�tá�!9��[YD����.M���)� �Q�ͳ3��� %�q��d	b:���qck�Lvf��b)l��� O;]���1""	?�;�٤����@r��vݳ���8?�$����_58�]Bҧ�,C
a���7��s3��S1��Fm�/��OC�>YH���@R|^���ڼ�F�A�_��T`�49X����!�d�/�|�r�2�Ӭ$%���^!2���d�R�(���Ǹ�|/�  W��'�����^�����2cDYn/�j��.��gf�������#k}�PyrWZ����k5�Ǐ�b:����Dd�w��|P�uX�1���(��ͼ��XMK;󻓤��(X�y�r" ��DD? ,��?�L�?m���KM��{
�_W�x�3�` �����q>��B���p�eE^W�53u���7�Vs���	��b�`{3$"t����8�o��y�m��O�NᝢFB�(�9���`^�������k4&��AUJ��!�a�Bp"���&G\-�/��x�>�\*D���׹�{�ң��4��.��X���~yLUGYtӐp)~V)�V���+d��: �����,YZ5':���Az��	�bٌ������^��3b˿�x�ʅ�A4,ǉS�� �s��� =���a8\�B,�Ot�71
+Mߓ�@�ON:�f���Va�E�U���!���+�r ����[�����R|�ȿ�{��������J3:b�#�·=��A#�[d$��{����7�"�r��G���Fg�i�D��9@f3L��w�+��C���z�$C����?�Prs�'e�۰~&�8�|(3�h�j���_���}l�F_1y��YhK�~6?�"
�B��[��Y�i����'G�M�ݓ��n�f?kK�o�yΨ�o�зto�������M��<��h��w��X嗯��P��џ=�ӉKO)8A�R,��2!3�R��_�mq�PX-h��&TnJ�č�g9��	����X\X�a>�_%����H�����=t�j6�y�g��[��c�gVV�l3��}�, �b���n�j��c�{�����gdROF}�fU�;V��&�^��Ӓ���$ �-~R��T��*�j�e��|�:j�A}�h�����*�٫H~�x�����*�����X��k[#��� vx�W��^$jǽ���4�?W*dõDiA�B��U���@���P�־�`5].��c�~qI�'�]�Z#c�P�%�박�i
�ﹼ��v��^}!ZW�ϴ[mj�귌o�����^|�_��)�hE	�G
К�4B��I/�k�����D�DT�T������u�[l7F�J+���g�T;Hl�P���<`�K��p+)A�T{-�-�-Eé�F2<!��>�%�P����'/���yl"mE��%�R�bg�^��7Y��nC
ҝ/v�p'^}<�|�
o�L����O�t3�T׿JK9z��Q�^���-+��zU�N�!�2gs�����FcG;2l���X\�i�o}��XY658���˝m}Q|�r���ܚ:1��$������F8KH�؍�7���u�P�2�_�V��u��[ �������k�@��'�X�O�����US r&�c� ��Tm��!x�Z�u�ߕ�,㻧��S��0�"�E�K��AI	������W��P�
ߖ8G�N5-�s�se��I	�C��.��4&x�V���D�f����h�h���:��V�Ȕd���9�$b�'
�(YiL:�۬&hh����?���Æ�ļV�##1{+�������m�����H*7�Bn����9���Ћ��^X͐�n!�=�T�.�kib��k)�Lq�O���.v/�d2Ļ}(�0��u����,��C2a�O�D�=;'��[�R���.��5a��_�B�H£Զ���Y�(������'53�\�(��CMc�.�Q�,�~J���^Gc��>LZ#Q���WB�`�C�z(�f�m�AZ��ImT�n.�ȁ�P��U�݅�I=[N�;d3�2��M5�P�
A<�͑�X%P��	�U{̄y:E���K��A訛gyÃ�1^��t3]OjZ^�Z�"��"��*,k��'#�����a�T�ahũ����zE�����,�:�u>DMo�O6Ϩ�Af��U����,;�a�K ��z�5X�#G{��-��Af�Kם�n��jC�=��G;����kZ	ؐ@IM��I�Z2ߝ!E	�x9X+p�*Z5�٦�o�\m"�
��
Q{��[�N]Z�H�\`w<���~�=��*���{Z��I&o
�[�-��p��{�8����#�->�gva��T
g�-kK���UH�R��hc�����(�a��aovd���y��(%�{��c�Oe�]s�A;k�N��{�Pm6�
�p�XsT[�@�fc�I�#��_C
"��0�_�|� .����O��(���E�k�f�iv�U�+`���5�2� �����7�fP��i���c��Ƨː�e�Q�tbi�{S��&�j{Z��MX��&Q& ��mA�p�/�=��%r[����L�\&eZ2-l���j��9h��s<ت@�snlG���{Dh�:n�jŕ�X�4\Jx4@2��_y�A�̑<z��a�B"*�]�H��ڦ�R
��H
�(����&���ŝ��E.�K7p�^4%XV���cE�%��qo�w�H܃;v����9�kk���h;��V��Vŉ�`��߸1�<���$#���<�[��,J��Oc�����?����ȂY���^I��UO؎$�:PsR���q��2�>�Yyd�\`Cw9Eo Ɇ>S�V�jEpH�G�\��9K���)_�˛��X��{�GI��(ww������/*K6k����DԒ���z����%�첆�9��=GI���Axe��G쯎6<���G�"���t�XA��[�)���J�r+��4��ј�a">�w3�V�eL�zS�I��U���I8�5�gu9�����d��RCIDG[W��)+<���1I�E
.h��	_2����5���Z]���`�����B�n�j��qt�OB�-y����9��e�')Ho�R��!���s�'�9B��� �`3�5&������ې�azB;�/����E�i�y���ŧ�x=��H�|�6�#�7��B�J����!����g���MNB #��:�VwT�B���n��ʺ�3�Y2E�2gָ��L7eӥIBc����"�
���1��7�Z�
7����=wߑ�H����DuQ��T��	R����׆��Q�1��;%���}�M��֡�OZ��ᴒ?��&�^�~TdW�P̗5����%�2g���%5Y�kx~g��� ���p���� �п �f�㛬��.�����n������t��@���{���O*8��+#;~!~^È�&lY�OA�����a�.��%���zS�sB:�F�```����bF�$�M�P?\�o����Åp����*opuD�u�4��n��ӻ��	_�!j��#7]t�&�[�a
��u5���Ͻ�B:�V�VעlxFİ�7��_��g-���z1�,ھ@d�T��J��R��@��E�-f�v�*�.p��#��PI�k�n{����n%��m��4�҆oI������#o��-	�t�� ��Zj�����֩��8�v�`������}/�����Dizo6�D
����������w���rg�J�����?�}P9#~S"P����-|��<�W�������3�Rو>ߒ������&�="-�*�mSs�C�����:�5 �_~b�V���0�)�+"[R��,f��k�vЉJ��<7�)��L�QR�@��;�!3��lSI�!@�n?u��MjVE�[�e���`�b� U���qV�t��I����<��QY z�0	�w�ʪov�ˇ�4K�Gg��<Q�ՏOﲬ���VP_����_�R�N�L�����כ�=�TC8�:�%�I�e�NG�l���(-ٖl���}�-��M���1�'�1 ��!4��G�%���izo<�v~c��:%960�f��/[	�he��B��p��Q��
l�T�H���A��x�)��	ڹN��D$PV{��
�r�IB�@S]%�Hf���bҖ4�ո�߼Ub�!�s���8����1�P������֊~�')��l�C�3�[�RE�1[�p���ꬺ���xFi�t+e�9H0�]��O�����?�3[ʻF{Q �3�.6n��� �E�
C��Sq��-�h����G�;��\CQ�yF��)�@�|���'��&�]���e�K���A`DQ�d�]c~*�⽿��r
����[aSKfea��4޼���F����RZ2{�= ��:B�,_�=�m��ւ�N	���wK��&�.��Pz��wJ5��_RE~�h$��&%X֛� sO:2%8a~Y�!g���E�Qr���;�v��N�A\螮� V�ф����ȱ:avI��7k�Ÿ�|M߅*_/82�M ��+FTǰIl!�1h���M4���,LqvM�X�����B�E��hshB��Mf���P��%���kB(n=��[ "���p/��H4�C�'.U�n�m�$�R8��d� ��(��u��KT�}�$e]8J �؛>���Y��]�T#7)8�ů"�ꏗHu1k�
U�Z)f�CA�s�>]U����U~7�#x�	 K�!�����üsc�p��Ө^���7ř|�b��{F
�C��ZE�Zz3��M�8���[�ŗ����щ�E������Dt}3��Ρ�?�n�C�E��ﴄ���b��pʋe���O�	(�<�>�w�{��:�^��?|�>/�02��x2Y�����;�k��S�Ƃv��M���V���&���\ �q謀�7��ۨ~A�&c��J�!O�H�;��YT5���t)�>�PA0:�q�~��_����*���̾l�4l) rD>.��Ǿ��m�!�	��ā(�i.�A]d�!-�����)��p<!�N>�~5�-|�<�v�!�.���@y@-�L`xP@(�h|��@H
[�������.����f�v�ꉍ���/:X�A`}��ίKM�Y�I�(��&:�~�D�ńR�����a�g�}P�����p�x��	�L�l��7���;t+_��[�� r�)j�L��{؏���xU��y�Y���{+���86�ǡ��4�;*�D���:(�&�WӺ��w��O"��-���С�x;��_/�%߲j
85l+�	!�}�Ǖ�E�8���Iޭ�C�$dJ��>�w&g�3�%
���;�6�Tf8�?�(;+2��@ |�nD�%}���p�,��i���;��g����U�L���A�>T��S�V���ފF��h)D�!�l=���,9gb��$`��F�`�s�iV��y_)����7X
���l�=���_՝p5���wI���xU!��e'=#%_�	���'>V#��_u����c>萱'
��/�^��{���H���h�p�]xN�P&V�@�NOؤ�2
��'ew$�\���X��]&nP�/$�y���>�c�8��}���R�����]�k��������"��_^��[��fۉ�9!�ϋa���	OF�x����l=8|��ّa̰^qN�c�Qi�	�v��جF�e�<��)���Tv���"�+�yY�k���oK���!�Ǿ�~��5�s��_�"���E��#��󨲉�)i��[3�������-��(�}M���qJ�����S�����`G����&Iø͛#Gb\Q���8(��jwU��:$�?}�%"r�Ds}�9�p���	"�dM���H��l�ZO�����D�g�V�o�x)�|�}�#�Cb{�
�Ų��ʐ������fӁ0�j�$ޙCY,���
h}���¾�����]�(����訌o>P��,���S�X�``���dsϱ)�p i�by#nE�b/Q�+k�ʵ=�RYA#��Ws�򳒾�v����D��6�)s�6g �o�8q� �a�l�x�� q�蝝 ���M�b��q�t.�I|�Юe�=����/�B�l�xQ����g�߆T�Mp��ŝ�Ʊ����צ�`A��RH�h�h���F�g3�%+:.�@3O��i�DI�a��E�<zRZFj�a�K�9{�ǁ���e=u=�V�Hr�ںŋa�(b�gD�?�
~'�T�li�Yy�&ul�CG_��X�2�2Nr;�yH��rF�.��<?�|ل�qSCs�#l�+�����m�-��
�^E��	�dX_D|(&����_q)�,�/B7�(S��#����������)�8n��@Y �r?��"�̮��ܞ�m�-M�L�w�ْ�u��xD�'���6IP�m����T#p[��X�`dbw�J]0 ,J�ē`�=|#R109�E)Ҥ8�,�r�XOfh��="SQ�
��׆8a[�/��oG��규b�֚Zc����O`�t�N�A�\��+$�3��ԢQ�ͶR�˞�[���m9a��Q,�<��3Qti�Ѵ&g��H��#��f������	�a�E����^1~e�p,k�=��$�q�~Z���¶ u�o�9�Kȭ����x-j����,�J\��.�dsC��|�I;c����$��~��R��2�Z+�Bg7�����3��5���(c%�~�4 �Y�8�vuLX)���G���Kغ���|�H���.�Ο��1�X�~�������I0*אuaDv����gUȼ��=i����߲�:4i}�@���H�H��^�@h�nq��p!v��8���M���̧i++�F����f�l��k|�0�0�^t�l/�
�U�=������4���,�,�M8�:˵�,k�f�xVۜz���k���3��]�V��L{.���K�Я	�[Ϭ���36�y�;��+�3����A��*��Z>�t�m�j�^-nq&:�J��u�ɣ��2����]5qa�4������+[�X]� ��$�|Zz����#�5�Gl:º�fc��i��[z���d��%�EHbN��l.�ປ����u5�X�*�����6Ĺ�k�sZ�]dZY0K�zK�x���u�LD�..70��@�Յ�̸��|�� �PkI�՘c��� f�!\�ۣQ]��3R��Y�,��LK�\:$k���C�k��P�-�yS5n+�Au��&aTTS)�c���D3�yB�(e���<��|��X|!w�R
2e���rd��,ඣ�m'� W:7�]'������h�L��u_$�iM��6��K�?j��4�M��'f��ep�<�H=Y����bF��Cx�WO�E�ebN�����=���?����m�	o`�,��ɀ�A@G�¯����~~���xX��f�y>�:x���b��o���S*�D�	����5��V����R\��`��9@�-VP�=Zg%��ޮӪU��G"{]*/�#c����F<Z8CNZ�;ٲa��רkd	���Չ��b�S����<*>)rĻⓞ?��k"��v���m�a�V���9��-27�Nu$�Wc�yh?��J�iKM���.f.L-�e�F����,jsq�2��N�E���/�`>K�y_b8��I?;}�Z�%��ixCz�C�/g^".5�~i�6���$O����.h8���DҖ����ŭ�"��G��G�e]��{Hy.s�X][�հkV������������푑�/�9(�
� ���h7^lIe<0�M�N����O��:�5�llç��H��L��fo���l3�A
�/���䐞\o�HV�����e�I�r��Er�߭%%��E�R�5.���̟uՆˀ�7�����_S���|�˓-��$�~v��6��i�I���_�������u�|���1�ڦ/�����q�4�ꧼO��A��t.����X35��ȅ�Y�2$L�I�i3��݄&��"1�abd��F��ѳY�Ǥӭُ��� U�ٴ��2�UaR+?�V*���˺���r��T�"��� ��7��E�&o��8f��:���Ww��y�%:i|%�7���ʒ���Yڽ� �N��{U�o��;޶�J�+�����מ'gv��Qw����`��f��}�����P���R�Y�����c��=ؿl7J�ʞ'��2M����	�k!��@��7����{��aJ� ʇ4��b����м�R��^�r;N@z�P���R���y���r�[��X���3B��ڏ0�}a?M�b/Z�.���;��i�d���:�Y
_���	�9E� z)�����Y�}�*�R���	9஝�6t7h`���Q+������=��� ���ne�\�b�Ƀ���=f�A}?s��0�u������q\�"��aK�C�E	_fy/��ߗ�fWӑ���h��[�Zzq��Z7���@�M�֥̉�/��^11���4�!V�,�p����|;U0�'���3ÛNw�c�)xb�z�=P�#�T��:X%����Z���1T����f̽6��egY��hn�= �m�o�1̬J�õ pDz��h9$m�<Y��u��݈���n�</�U�2nd6�bKslu�6��_I�,(�ިx��*�ܬ(U8;��p8߫�z!'N����^�+=H�s�#�i^��Vpp���7��̏��	c���r��נ�[Xۜ?�X��Č�ne�+��@lP�07�il�T��\*�y4�Ef�>\W�l(��_k�G6h�����i#����W*�]��#?JSN�۪[��wM��p���B��U0�G_��x�- H}0Ii%7�~}c�_{�����d��A}#���x��V�bQ��O|_D�ڦ�r�:����a�2ܒ�"3�!�_����n��M�\x~\������Ag�%��L�����7�_u}��� f�nQ�&{�/�AJ��Y��-��j%��r����
ƸdMw������K
%;�促#��	����%�0��l�r��=xU(le�^�-R}k����5��5>�w���w0�~��_f��jG�� ��Ƥi��%-t�\���[��	��^bC�������2�a9@�����Ě?�����������sY3b��#��>�J_�P9�:ڹUQ�J�����d�v�cf"=6|�Ԙ3���Fc#��`�, �"Bt��u��5�8x�B\}�O�Pk^�F^�F�I�I��b*�����R�.� ��zr����m;�a��������m��O�g��Pf�^{��i=c_�|._G��_��6������.��ݽ��p��]&5�5�L{�I��J�.������%��� WY�jGm�`(�LbB�	쾷�6w>�����>J�g������-g�	�(�G��ȧxZ��k�b<��S� �9�y��	�'�[/�jCf��)���V@���5�(Ld��d���0�5�ңwj�Q�VUG�j�N�I\F������JǼ�w�1�v����U�]G'��y����r�� ���as�*���Y�o
C�(m�������dEY�˔$��8ܫgPF\���Z@<F�0>�`0�ޢ�g3��+���+��h�Հ�h���Le6+7c�["���!��B��3k4F�SU�F*�ǐ��h��>?a5m=\0�C�y:�/9ծ���R?�:�C=�Jѭ�l�!s哎�_�����ܴF��^��ЖA��M�|�/n�<ˎ�s
�k�t�����9�bc�,'��m��z�s�Ȯn��9����ȫ�dm7;�}*j�xt��9l0�vZ(����3����{���y[����Ȼ�ؘ�2�Jy��&���D�'�xФ�֕͟��x@'�8��қ����E���_-Fа b�=����j���mӭY�Ҹ� Y�x�����r��!!*$�}/ �W�S]��6�b���o|���S����)���.�/���'V�������5�2�dS�.ga"w|����d�	�K���ZdQ�P�(C[�{�!�8�&Z�qIM��kf��^�ě�p�_Ze�rܙ��;�<�����*��3�k6V)�F���,�`��]��<�Vv��(��ش �F�oȗ7U�_�c��U��[cr�a_g���'�&����S�pe�Q�W88g��J�sYD.~�R����gۊ�Ve�Ȣs�!�<�d�7�Of(F���)�E*��"޲3KGI����,A{Kש�1�G#)yi��l��2�H�YM6�1�a7��W�0x����?�E�c3r|?���{VV�.ˬ���p�������N��/�[�B�`d&��&s%@4��|*xgz*ɜ,/�hn�h�V���|F��z�C1�U�8�=����De�O��ꄍ.���1�+$���֫�ck���aY���l�?9�����Iv��>�z)�\�sKvd��Y��q��d:[!��z�BJ�4��YB�n��OlX�g$�5>���]9E�p�I�J�	Nf�y�J�J���$Ly���Zv\�B��F��D
�Az���cS�PP�|�a�e#�/j����F&-"����t�!y߷68<�p~��f�bf��c<�}�f��y9��C-oQ�Q�'zj��]@J`\�\�����M~4w���ԍ&�7'��M�:���TP�����u/P �A�,o�y�������{Sj������o���m��L��r�o�nޢ��w��gt�Q��H�����B��(GF{��RYa��|�^�BS��u7�.!�j��9�%UcU�h,�v)���u��hp���R���t�`&��ǻ=k�������6}�����V���?������>�v�r�4�+�&.
˧ʖo0�b���ywƗ;V���V4K~}d]��A=*�H��0{��F�P�$�5x5���h�Z�/y�hE�wwϸ��Y�Z�����Mw\�r�"t��EnU�� ł���'N���פ�޹ ���F�	�t��F���)��2����
�,�!�)v�%>��m����X%)���*�~B�8W'��_*�f��KH��O$�S-�D�4m���4����q�0n��9q�(�@���߇��8KU>l�ݥ���U6,5���Y�,|�H?�s���LG�*�L9�q���MN���qE�T�=O�6�=p�>*�N�>��ی����y�31"`����+���AS� pK��@H���#���QzE�j*���~����S�5�P�}�F�y��R������tq��X���ۏ�EE��j�/����kW� 6b4���?6����5Jʄի��I_-��˔�R��WtXEJ<-*r�OU6y�2߻�7��{���`�HuEH���VV~��׬�C^���k��1��˭��IN�(ʮw�u}����8��*�2�L���ro�	A>��\&.[$�Wn���Yn};�{��l�:+��h��j�	�]����N�y����K������~$#^\� ��3�:R��9�6����[GH�9�ܲ�ܹ��cϳ����=*7�&}����]�k�)__a�= �XM�yvZ�}�Y_��N#����������\I���1��\ۊ�?$k��@ڑ"�&�������{Dd�T��!�s�z���T� +�s2xosL@bM�X�6�� /���N؛�F��#o�=�aJw���l�ʓ�DN^s�0w弧�����M���a�r��� �	Æ|PrEJ��JB�_�+�����Q�'n[,�ȉ_Q#�9H �rs
I�|=� �=hl�)ᮨ꾡s`��=�&��%��>���
?Q��3���w�1�ձ)?L�������w���YC�l����,S��25(ԡ/���2qu��Ds|��t�a��N��Ę, �(y-�L|�!�b�o\�x��Z_;ԹkW�×{��*/I�d��1 �.�m�[��w����[��o-��r�@�!0N��,fh/,��/�����Q�|༎�p�w׳hp�ܓj�e27P�O���v�š:�|0�1>H�fb��[L��&#I��}K>a��L1A��i���~�m�#����+�]�W���C�x7�9-uc��i��z�oeU�5����8�Y_��{��Um%�^�i�=;��ڧ����]W��rl��+��&���k��(�YG��9��%��p��y
�%��&�B�j1����H�{��!d>و�b���6�~�a#ǹ������Ǥ�%ۉ�"��Gw�w͛n��.��͡~c^@�8��NY{Y&�l>a/�"	�7e�
�{])����M֛�������3��t��\�.�����\*N�����5�c8���Ԁ��f��߼���[c��\�[�b%���[Z�{,	fz����e<�Xϫ�Q�n2� �3
d�i�)=���Y�kg�F����QP$�b��U�o2ࢉ����.���������>��}�R�w��@*u�n��D�_[�9r:�͆-t�{v�ܦ��������!�7P�6lݶ�;��Ta9���ڊy��;f�U�Y�&�*�e��;Mz�5 9�-k��	�b����ͦ-�
���/������L��rE�T��+�VC�G��'���`��~N|��g;5A �
��j�LD��9�Ab�v>Y�+ϡ+����ޘ�^q?�����NF˾.��)Ҧ��#��&��45~�B\�E�k�l/Nϰ����9�31ߺ5K�R�"��1�r��|#M�{���6�y��k.�紤T�6�jY#�̥aFu��BK�ZFҥȁ��I�I�l-W�?�ٵOg�8D+�E�G��Hl�E���� E���vk��+V�ΆD����>�u�K�cQ� T��M���e�=����[^�.��H��J�ܷ�\�G �+0�o)�SB���fǁ�`�ժ�gt��>�	-�G�$cqW�z�T���ߑ�"A)r8�4NE�L,A���9XKzrMʻym�5���O�nx>%(��(m�c�4x݇�ǽX���m�!)LL����#r#��'�	������T�%5�fY�o-~?��l�xl,�Cz&��p�e��Y��� P���Z�!�t��i�φ����93k�tǣg�s�}aw��o��C�zem�����g4�Q�rN�$[�����#tt	��`��x�i�ף�L"Mh� ��-�}�|��,��[���%����ŋ2Kh���� �ϣ�;19���0�s�t����:��$c(^0�a�{Xѧ�C����N�``R�R��.W����YA`�_A~t�s<�U͞�ɯs��2��.�����x���,ʬ]yL�J�G,�߾����̚&ɮ<�ɘ2{�m��;�v�"F�EA}mľA��l"
rׅC��Jk�35����#�v�&Z�e)�����-�/iQ��''?^�rl��}���3�e���W�J�MK��u�:L�#Z�I:�t�Jꨈ��D���g�*q��9�_@�9����朲IϮ�" 0�m���Ъ�L�{���Q��--��Vp����`Qn�aG�݃��_��'>�T��;�'�c�wډ�!Ҭ�9���W#?f�i�-:K�����l?C���ԡja}���"s�#ȡ��;}ؓ�Q<�T���eĞ�J$�W&��&�;N_��F�n�~�4�e��~�bxw�����xsh�G�ݡ ?MG;�W��N�ă1@���'��	�؟Y7k���et��(`H��V`ȿ��bc]R2�8gJؼȶ�|2"�»B�]�S���<�J~ʬ�.]}��˄R%�bձ��Q�A��d�)��O�V0/�����!`�a����oQ/�t�T��$r��d�p'��)��X\����ŲG��Kv/�m��W!:��f�����j�$�� {�bϢnzv�^����H[g��6�Ni�!�Q����y�N�����i���ʈ���<J���M��od㶎����=��Q�kv~�l=K�n*�}�;�(���<�ۇ��ڮUu��I޲�Y��KB�:�\v��)'#���[� >��N;l���/��X?���6z�Mf�I���g]��������B#T^���f�%��4[d��]�X�zK�,,�4>��]O�զ���MQH^;�)���UZ�����|�P�G ���uI� �MΥtO'�[��\���}:ǋ%$��	��څ�Ѱ����k�^l�zv��g���^(9`"��[ꂋ��1�qK
��P�9_'Y�z\o�b�Ü���G	L�E1�TV�*O�8]��^I`�4�X7�O����M{Е�t�zT��?����C㑓������g�V���ޥ����_��\��9�P}���T�C��&��o�c��{��/��:K#u!��(��Q?�I�� �!lKx\Z{���%��l��x���
���KRW(�<�C<�6��w�ٜKRF1���0��ĝ�9��蘡�G��}���*��˒�"8ܷsP�)ӫqZif��j�����!*���1�S�&T�­��ʃ;�&ן�y�^^�Oz��i�^I�=�h���+eB @�`m�X ���A�}�(@�co�.�i�\hU��o����
���ΐ��}J��S�% H7&Z��Ϋ�_����n����t�{�5ȥ�=���N�od�!�)� !�>бߦsv3�R���GFm,�b.<T?���ma�n���k�5梁��q�Y��t�{/���Kٴ�ApM21�z���v���C�9��C�%��<�C�M�OƛS`,B����+����=��eu��WO7zɂo���O�]�.��:1_M��>3��KU�cꑟ���%>�勩�ʫ^�t���	�+���b*��9���JdN�����F��ϥ�x�5BL��^F+�(AK{%��zD������V�tL]�N?b����#�0]^�s�����L�k�e��s��> ���5ˮ�`f��
�z�N�H�Ӈ��dTV;iM�gXnm[cTc�<oR�wmb$�|˖wx�s�
�Fe�|��ٽ��ѿog��	z��7�?�<J��6�0�X�jخS�l_�c v0st��2z]:��{46l�Nx{��� E�9�qor�=�p��,Tp{��F?�+�F�$\;5U��y�h+v#_��qJ�1�#"�~rئ3xNA����Ԟ���qHإ7�N�վ�¿�]��1�o5H���shtF1�B"�[��ν�Old�`�5�9k�|W�����v}�#�D����}�V���ѧ�����I�`+��U$/KT�>��h?x�ZC�e=�kIKL�PBj��)�o)���ٷ=rgFN@�y������Y��)g􁮛����+N���zd�1������.0	(�h ��2�Ȋ����)M��V���}o�h��$a�ʭ)ϱ@�n3Kټ�a�凎�fZnj�����j~_����5{KHXHg���U��G�S�i���Hg�Y,��D/��v��Χ�?j����C���R����j5��7 ��0�u� W-q�p�[�\��ʖ[�ύ�V�&�(��̽uN߾잭4/�$i>��֡��`�g�L��9�Ԣw9���g�\�������������\5��w��H>�_Rf2��Y�/����	��]�U<� ��*��o�N��\k&�O�c��իt?�z93��s�k�6���M-�WD��Ƌo��4TYq�0r�r�	�,���v� ��%�ڊ��?��\�3��zx@xx�T���j��(gC?n�7�fIK�,%ㄨ8�C��]
q0qF4h� j6lĞ+CP��o�І���)(��T��i7��"kgx�����"�2}�U�UT�7P9�_���@�e!�X沊(��ou�g�jWj$eU,K֎X*7�|z�s�����)��}E�����U,�.�G����^��/sAz��4�0V��jT���;K��a���'�7�9�d�˽]A��U%�'9�_�e�x����l,28�Y�)M�qI�2u��(hWM���9���m7&ONN�Ez��j�3�Sm-���견S��'���v�I��;!-*�l���f�W�Z�������	��qn"�O�V��|4�:�����ɳ�,�w����n���m�'��=:���Hl�Y�`U��ɛH�f���?#/�=�4� ���F�`���$v L3+ ��}�8��L�W*n��C�G�˷,��ݩt<�.����F?Fђ���S4�x���h���B%��n�>�b�C�:#�x�eάY��E/�&���8>�A6� ��T�̈�w�^Y�y��`��H>r�#�t8���[P���׳��[�#�q�hp�Dz��N_��� ?Ҳ���e���L�^ֈ+#����+�)~��泪�j�:U�-���x?��h����S�j/��ػ@9����H�&
��3׮,�Bd�Ʌ�Z��{�����
�;��h2<�bn@T��_f���Ҽ]#z�9|ܰ��N
���ň����NfM������eQX�=���(up&��M)�g����ki�??M�T*�j�j�����Ԫl'����q#���^����T�np����A��uD�o���`̸�!�UN���IA8 /Yg�֐��Q�)4��-��>J,�M�Ow�2�k��#0eu����!;U�v�OAV�JH�ܶ�Jil�!v����ٸ� �Q<uf�^����?�&�Ɖ@�C�)=L.�x���v�2�t��K�G�@~h.~���<�B�O�a}hN��v����)�Ǫ��������jC����*ͫ��a���X�����28��Ŋτ/��id�&�"1?��[�h9X:{B?���6�rn��by�td�hգg�W`�~(�Q�'�C���� O�;x���B���2���/�$Q5�@�:��{ˆG��Ǩ�1�5��N�R\8���B�����wd8��S~߂qR1ځ�f5��)�Z������"E/\,�C���,<E��ƝqR��î �I�\^hp��"N> ��~���g�"^�|��������~85g�LZ�Q;�����#���t:�n�n�Ko�^b���/}����������+�߀ 0��*�S9��e�6jv���Y�n�6S�ˍ�W��}�d����	�ǌ}%BH���	�$�F/��_�!�e=K�����8p<�����ZTX�;�nXQ�5����B���E �Y+�9l@vn��/�ږ*5p�f��\�7��f���'����_�+	S���DO�� b,�f[ (D��-D�p��:ĩ�!�͙#��K-.����?�H�v.��Q�i��r�K�Μ�ք��(*�r�_���K��{�k��5H��G)-h�� Uö�x���6�������?XI�3 ��#��)X�u����ޭZWi���l��v����j�ʯnޝ�?��i�#eW�Їz����E�->���}�Ka���q�����j��K�f9�Xo����1��O��y�����=�<p0I{t�R/�*�������w.��aA1�ؼ"Ҹ䢧�q�IH��SV.fKj[�!27E��$����[� z���Ƕ��W�Ml�����B�����tdo��pg/��Yt�$9&�B�:��vT� b�X��n#���fpgt(���0���.�S�ZlJ
͓��0̔
�x�ػ��#�f�d���{ܜD�h��#�ܥ��	+ޟ��_<�f���T�\wfeQ(z'�� c/��^�ћw�(j��E�$��ӎmq8�m�}���m��9=d�Z��yX�\�1��ѓ���/0��"ۊ~Y��X����6vQ6)&��}y�5�l�\&Τ}1L�ؕ������W]�0/'���Ʒhg�x񾦿9��/��۶�C�\f�F:0����C�2����Q)�����2�CE��.�)�V�,��f�b�h����+�G�j�7��ܘ@�TbF"���}C��g~4�Ԉ���V� ��ew��$��g�w�k��M�� =w���A/3/j#Ϣ���o�}."���ң�3��岰X�J�4�ú+�:�i/�!j[VT���о��&`"b��	�4y�o�Ix�4�����JTÌ��_n��g�*m#�PTo�9D��=���◢0'��Q[���xu��:b"N�%\|Z���S�	r��m{o[m��sː�iǅe�_(s���Ԑ�{ڵ���s���W4,S�⦛��ASC��^F+^cSs��.f�D\�C���1��vو���o]�����D��m��6��ķ��!=�䑳1ϹO���TDE%Ճ���-��S*���t�74:5��N0w�&!�l4���iǜHg._I!�� ����/��Vx-���&,[!�c9�u�a��͘����1b�ne�n�@1�E�.���Ȟ�����
m��b�o�f��h9�lv�{2����S/�}�s"�E�}ݘ,��Ģ���
�"���ڽ]�c?	�Q'䡉w]Po� ��
�yQ�lY%?�_*�`p�&�� ��@V����a��v�Vy����@�/=��c| ��H�p�2Wq��x�6L��C�ʟ�ֺ�|,k���f5h&1yE���a�@M�Њ�.R�m�VK=Z�VQ�"P�b�F��-CH�����X�~2����Ta�:Ο�&�i����- <^�3��a镍�+��D�<v�S����􈿪�wL��P�����?����������`ηT��B3�^<%�2�r�P�D���F_E�v(�c�I	W�zfN�¹63��#���=�U5Qo�1A�"����[��&@@0TJݵ�	��C� �����SR2K7��-��y�uy��%9���a�E[!��'��n�R�l���H☘-5s��.�����\��7d0S�=��BO�1 I��GY2��y.Խ�bl��
��h��:[�7fU.��P����n���'H��P� �b��0���nK�����\��7k�"LV(pv2�S"��z���(�ʒ����oȁd���Ƴ�0ekf m�!�r�}+I�ŏ�k� lu���h����5�ij��']�E�.�wEe���%ZR�q���z���"|/ZI�B�i��Ec�)�b?�!��{�Oߎ����M�65Cr�A~�O�rx#�����������$�����/�F��)�o�9'��1���</�g����=��?��~�գ�WW���eq���M���|&������!/����=���E��8��;��cNգ��{�u
��V��w�\��Q�ՈT_��� �M��U�������M:����O����<0��������W/[#��B�e��7</�'���v�S�	���|<f�@�jRN���3F�����J��e���+S�o�"����t�A>�l2��L�r�?�V��P��U��P�	�>�%����S����P}x�.ט�f�R(�.Q]:�v47��;ށ$Hq�V&��.�j[������G~�T^8��zXj�cH����ړ�d6���9�|���p�1Yɮf�*�f��S��D� 4}'��l~�0�)J����B/����1\�pO�mGBkS/e��׮�$
aU]1ȭE^o�.=�0�����$v�^�V��B�z���b�E�DN1��@v%	���{&s\3^���I��Y�Ȏ�1�4�4�3'�1%@��,b�ʕ�!a�L}�U���<�p}�Z��<��l4uk�8 �7���Mp�xy{�'P��G��{����X�sI���	�r}��Xt]k���.&�mM�eW\Y���c��o��U�Fg[�����Fk��qq#"Ҍ�{@��/�oCaA�Ƚn��������l�AN}��B��ϛ.����\��!
ȢEm�y�A�m:�t��(�ͤUI`=��p�F*����[Rd�×n�1�A/�뭺e7u7u��W��Ꜣy>&���\bm�A'�ъ���{��ϻ��@w��6�	����3��s���6g���X��,��g��_#nS#�+�\"����߈&&t$�^�e-��Xq��w�S{�.{<Z0)�� ��u�+>�vZ U�G����_"� ��Ӓ`M���B�꼶�/���QS�F�f�ׁ�`"L��Bb$��l�I*o�,����}�.#��;����D��ۧD
�Sk�������B�p��gYt����F��9-=X�) �n�6���(>B���Q2���Cn���<��ƪ�+�m7;�r0o�d��\�����9k�Tl��0}��c���I���{sM�R�!���Q	�c_�0���t�C,��۩�����)��������/a����p�*�5��En�HQK��^��)}�%�-i��[��@�w[�/���:Ur K}y�$FSsפ
��~�ͽHNO[���5k.��c"�UEr��ہH�>�i�4��,|O{-�p��""}�9�?���@σ�h�&����AK�<�O��i7�A.�%9��Gx�@wT8mܵ#�C�6H���h�b1&_��`x��
I� O��p�r����K%���5�Cb��\��n��g����^��`�+K2l	��&��j�d�#x�4�PSIj��iO뺥u�����ݿ$�����lÿ$�w���>f�Ld[)op߯3~��9Z�/?�b.Ὑ2�f!��f`�|��>�$�:6X���Q�Y+}�\%����jc|��M�o�X�� �[� ��S�C�T�s��k�H!�+���t5�¯~������&��9/�Ȍ�MNx<(��V���2�ͼ�2x*M�P��.3�S�R8lڱ �V�+3e~-^�	i�n�tT��0�����t#��[�Vh*`T4X�����HC�-�!p�ܜ��>�/��O�{����Y�+��!��-W�h���Hm�B���������w�.��P�	�z�y�'��-d���Mh��=�0A���w�β�G5�o�&S�`c%5g�]�د�z���(5R�b0y񨤁b�Bw�l�c~��l?�س��8�E��lЯ%�(��)J������|��]�ʳ�����_�:�P ����F�F��B���h�\x���V�^�θ����7��PE�h��D�2.��c���J$�մx���Dm�סp/��].�N�cr��O�3��MM;c��{�� ���@��p|哷h� �;U*�.����g��.���f�����(s��R�B�w�h�����s��������(F�ԃz��`2���53Y��qA5{��m����`IG����)3|�e��"7G�~z��l�w~��� �!"Jt��kGvp�����wVb��4�<�IXh�S���G[Ta��$���P�����K�*� �tݓSc#���T�*t�s�Y�*�Umd���ta��T��(�O�W��dU������Ԁ��f}]�!_n�i>W�{�	!$C�O�� �Ʌ�[,�å(�Zu+
�#獵�܇4�l6�����g�-�A�xe�;�Z���0��֯M{�J�_;S=�O6�L筜@�������3<��E5=��&D��'�:-�M\��+����a��aG�s0�$�~�$�����j�2�w�'� 0Mfȉǳ�ې�-z�:��L��󫢉���s,��F�G\�WW�a�7Y�YD����!h�Uz��]yn�Rݭ���"+8 ApU[����~Zk�.�3r�(�8�s
���>\d�׀(���{�|��R37�
��ÝXj+y��2�{>M�ҪWy<�������e�S�_��P�+�?�1�@���3[z?G}��dVb���%� [�y�m1Ř��k���an�ںh Bٶ%�@ر[΃���9�3���Ù�VN�������ݓQ;o ���.���K�
;pwX¼Q���dΊ!8I�`���.��(�(��WIKX�D�0PQ�l6���b��G,���sI���qmLX�ג�����(�N���=S�)ψ@�9�.���oP�ot
i�}����JK7�]��][s�I?��X�űK��0j��Ⳮ���8�݀г&�#b�Vn�.Mn3��߾J�����X]��!�GI�L��,z��pi�	v���$��#ܹSh�d�����YM\��I�{I0P��uu��.ٻL�݌�O\bj�J|���K�VM�F�q�t�)���$��q�`���@�8qq�]���?��1G/+�{��c�4c��,�Bwdgk�<	����d�����]�w��V�ܳJev��4$����39����pZo�t5����.vkN�+;2�S;ը�$������ ]�)F�y7k�����*	0'&h��n_I�b��@`��Om�?4S:��$�{iF����6��[�R�FM{7��;�bPjN1��{�]���h�A��D�kE~=����a��y�g��`��%|�6��nC燗� av",�mӯ��%�k��{̈́}h����RV���<�*�z��ӗ=�6�^�
���jW���u�������](�І�V�4U�h=JT�<�n�@޺#��"���ӢV�§�16�(���Qk�9?E5�\N�] Cs8�9��:4'��|�U1|��{�p�a��X&�iց\ƞ/u���� �7��dҝF���W�sUV弅�,��cL��r�����k��b�w���昿�M����0a�DOT#ۇ������P)���$Hm��C����W]�"5����?h%�0����D��LlEd'@Pv�P�*a�-U�jt���a���S����q�ƒ���]Êv�6 �*��dʹ#�r�8Z��k�nO��IH..��ٻ�g�E����߀i��y�������x��P\/�ƾ����:O@�'��<� ���K,����С�UϨ� ��}�,z~��C�E���aON����dĞ��n�>�m�tAhd>v�C�p��[�4�?��0�oo�2�H����\��!t�oo.2D��C#@�|�#\�y�/�A�!�̖m!	��	�eiS�%�2u��f��xP'0��@���?TdSG���-�����7Z�"��[�vY)�&��쌸�"?~iP���R� U>�l�=�����B�7����PM��Ӓ@�`�^�|�	�'�Ϊ���7X��B%v"�1j��L�b�Z8?��ji�	;�
J[�o�����G���^m�%ʀ�}��E�5��$SO�x��㕄Pq�_a9��@�e����!Q�v������P��aw�������<�e��K��$�pj{���:�Ր���»����7�z��[<(��)�<�1�g�3�t����򅂵��>�2�6"�(�x��CY��P��߈�|������|X�|5�A��6)
����"T�E�����!���]���$��{,����Rb`�iI�Mv� ��� �{\:�)%�JR��b����ݾ�ab�V�\W�M�}�`���gӸ
�2*苅��ה��#�ZlJ��"��R����qt�K�Oh*OS��^C@6�HI,nM��-�J�8�����%a"�=.��!�>T�����A�؂=LC�	T����SΎ�r��0�ۨ��o�u��j��#G`�`AƑ��V~I��Y\��!8C����H=�5���c=�p'P�Y���!r�����{���4�I�R����R*ݏsC�3�-�����6��n/���T�^
Z�4��U�o�:��b�'E �S���B/7Bo���¬��^;�E���<�83����)�p�/����wKt��i1$��>�	�2�β&�_����	�u�mr������)sTH.��*�i,�=��-��D�����P�������(L�񛥦r�����VM�Y(��:�d=�)=�7"u�m+Ԓ٘�U$A1�O}ݴ�rrQ�,v�Y9���#/��bC���V2���
)�2W������f��2y���.�#��	25<t��ey;�ORJ�ԇ�5`N�#l���8�2�.�:�T��eKd�c������ô)¿����]������r=1���ڽ�aڴDp�rv���8����զ�p$!���Az���T3��Qp�_���b�����IM
�Eג;d,C��ѯ%��.����ͻ-�H��$������wM��9ˋ�@���S���v�q A�J��L�$�M���]��`��qT��7+�q0�}��{�{+󎢶������mw9����?f�#��O��0Y��ЕQ|���(gò�'ѝ!�XC`'�G�&0�"��}�pM�}���D� ��f��6d0Nq<d��s�,�#�gU}6�Ϗn��s�)��B���qJ6k��a)3~�]��'�����M=�.<�F�ҝh��^���X�1�18�U�	I�gD��ke��T���7��;Y���`�K�K`���Vx\�}�J]ɖd���_헻��R@���|�X6�ҴG� �sm��m �n&��y�m+^
�^���Ec���B��sv�~~q5>!U�8yW��B��
^.1u�*��1����I��qA�_��M�MD6=�C �)fr�U���8��'�쿨�AC�A2I �U"�(���Y����E.1S���(���`����o!��!�U�wԉ��Y�tZ�^Ը�;�1e0;-��,��@#SXؤLD��JW6Jש>�>}I��O�u�Nh_i������4��B��B��i�hoG�g�f\�WxfA�R����ڥB�Ӣ1tۻ�"-�� �7���80��=F.�q 2єV1}WK�u��.2�,�m:ԷZ\ qx-"]�h�L��M�������8{I�'�B�P���.�7�v$Lgd�:
&
Ľ<sE�a��X@bm*�9_��r���<��Z�̊wE�&*P#�|�zr��$��l?ȞƉ�l���J>4�5d�ڔ]�Htaw�(��/b�0ɬZ_jݝI��F#��E��b@���T��I0�E�h�YjKԠk0�J�R����=AVc�Y�c%vglN��[�\(��*�VD�����3���I?��BDoyj.?Io��� �ڡ��D�*T
N��w2%+x��ֈ��+#��Vk���^k�7�_ "/���O�w��M�m7�����G~�*J��L����o^�)��P�d]|�	|4$��It���0��$X����&�o��VU$v�z,�JT���� Ɠ��d�	�k�r���:!��#hU��IlB�2{x�'�������ДTga�j!Н�t�7�H;���D}���C{˾컪>鍱$���m��h�=Tg9 �nΠ��ޔP�xe"�a����ӂ�#���:�"LwK��Y�y����:�>����9�˲@j7�n+�n:$�$- ��@9��Z���0����h��	3tm:G��j�y��)�����T2��&� |���7m�$T�_�9 �Ӓ�%��*ۅԏUXn$��~������-�� n��;��D�V�:�DX9~$�\��U
x�(WW�-A�!��ɧ����V������(�3!_%�Q���u)��y踁��筧�8}MP�6��Kf>�������hU�y-iH@_GS�N���\����h�bngiPa�������m���VyF�������=��#@�q%�8�����(|��zϨ�4���~�����Z��Pc�v���΄�&ٔ
@-uM�g���!ww������Q�5��Fi,i���?~讚��B���9P��w�:��p�`�	�f���|p�#�\0s;Bv���^&M�7����Y��vi���@۲ȯ`}�l��Y����F!:��\;AY}���r����D��Vx�H�#�m�������M��G�̂2A:�f�1f<��˧�ɕ$�FR�.Q%������f��[r�,3�L�Q��	0���u	1&z]s�b�����ۣ��J
ů�\ډ�=���ZEiP�O1�r]_~a[E+������U��5��Ud�M������w����JNi�Xk	������2�P�J��Q8x�C��c'q�;�l����/q�VpK=���z�j��3�[��-�, ]}�h�FT)rۨ�!~��Ø�;z�0M����	\�[D����n�$�ΟIӡ��g�;3��˖��z�kŌ�����������c�;�TE�I	�}�A��3&����MX��D�Y�GOf!g�Y5�Zm�@��x�3��|��ج,;�8_ �r���r�t�
ܮJ���h�iD��6�8��&_g&��tb����W枿�����'�J���h=	,�Ny�+7��@nE1��T*��x�����/B��
��Zb���;qn�8{��n.�k�� s���hf��POԇA�)��z�?�׹��9yr������VG3�	h&�6�:_֫�T���ߊ�C6<���P{�j���)��
��9��� ��� w3c��j���n�6L���ۃ�:�ia�R����(�==�j�kd�H]��Q�?�ռk�#�d� �٥Z�������Y�j��=�!�(��i���+ w�U��7�3�^B��_�I�{h8;�c�;�"��z"�/��`o�=!�/2�\z'J�1	\�f��]B���Rx�g*�D#&1C,��mB�巄���@������N����9V�^�%��a���Ff�wUQ^�Z�Gn�ˑ
oN�h���uN�"������������0�ۤ��Ę���RyS0��/�Z����$�����LR?KD"�������HPv�d���1�7��(6�M�O-��![y�����h��>V-�:4�"usY���^��@�S�� ���3��C���<���&�l�3����\�/Ŋ�?�5,�o����Π"s{�Ӝ���l��L��
 A��l��g���vU#%�=��E�C��r;?��L�+ �lqk���>�*�i�)��2U�� �m��̽W|o���`�������+uywe�>:o&�d#��3�I�fK��ޟ��"�p�w=�2�'�� ���ҍ��1���t��3�xѻ���)�M��Evsc��ب���F6Thws�2���N�|��;�i�?f�$��~���؂ﰱ�l���x�4�A
�J�ӏ�R;&����3% |�S�8u}F���H��t�|V��Lg�&V
$�
K��J�OesEfQ�����u��1*o[ �� <�(�����)�9�����{詌�u����2��hx'\
xu�d�0�N�y�"�����-n��`���@h�@!���y���=z����j�I�Q�x��Cg˷�jrΆ�R^5ݚ,��]l{�=�89�Z�
�*�G�Ԇ��Q脉 ��S�Ԉ�j���V�'l��B�-��T�`�2�v�ܣ��WA�`�:Y���*�02��L��."�#�z��'+s�K��JD��+[���7h�q���d����D9X¼s�d�렮6�~�%)��X���a�O@TQ6�$�!L3E��R�R^�����~�1�?�߼v��"]��/O�-X��A�ߩ�j�V�~�e�z�$�o��C�JR�E������p�6�h���#%����(!xt���ov�y��rn&������X/�	��"�N�B�[XQ���v.��yM�#~A��@��W�C�L�)<�u�< t� ��g��M�^��}�e[�����78�iV��4���:7�I�����������b��y�B�>��MR{�,�zs��z��v8:�,?�k�S)�6ҏ�6i'	�;@K�Ȉ|.�B�=���Ġ:��5�3�ǆ�c���PAc՟��WA���/J�A3[M���@g�V�5���݁����ڹL�_&��
��^�Cj-������5���)W���6m�v��T-_��;�Qa�q����w	���Fk���^�?�]�M���I��3�s���� i���M���2��}���A�w�X��]�'�
��KA�E���	t��`Cu[>�`«4TP�9Z��1l,,���v�\�}]�RXl�R�h����J�s�uy3�[���+�ҍ*���h%.)�ӉA�U^��WX��I��e��	܈��;��#��Yϰ�JE�d)n�MDpf*;���9�Y�KbM9�થ���W�G3�r�� �ص5���M%Ӿz(Wg~p�To����u>�hԠr���8���r�����`�����]O���Ҝ��T"��ѩ>��^G��'���g6�����n�L��6�[�IX&w  �K䴒�=��cXQb$��ц�X��y���D���$���ya8A�e�>Nz䕛�+���k}F"���0�2hEp�.|8$m3\ZM�NM ��f�Ë/yMh+�A��a)y}�&:t#�wl���f�$��[�v�K/���l%
�����l@����>R���'jd��Ȁ��_���rX���
¦/˩5��n��f�?^+[�1Yr(������׉1�>����7��X�^sE�kз=��~�3�9d�l薨�ر�(7!�2�(�I�})�n!qi�W����iư�7����$3`���6��l#_�iQ�Ow�K�$��F>�o��k�jm{�ʱRI�_|޷��X ~�����㿳'��p�H��JOl=f�Q�4~qFd�F���E�EIY�߅�b
�Ϡ��
�:ƲR��_��Q�.��a?���$I낚��A�������XT�9n��up�t��u��W��o
�����e�iB�l��	]E3���6��{6=��ho {��>/�{�UY3?�G���~%�O֨u�=\��Ŗ��nR�ޥc�u��x�����d��2����'��	0�}�n�i��H��b����#-X�\�ه�s�ʒ����Ć�L�?�KǛ�4}m�ǋ����l�h�%(��aA�|�s�&=N��T�I�י�錴�l�c�bƣ�� �#����l�B_oњ���${���(4��ηG���%_��5�.[&����i̞��P0�<�'�?0'&|�?(G�F=k�{_�G�\�C����N;���u����R���ˑ��=
�眴 �#�U���\^F"\S^$/��	_H�$)��������)�X���'-R�������ĩ8_��?Co�T
]���_�R���)
�&�'�Wɡ����oK����!�gd�P�pܙzX������������h�A�!�������e�,-��'�u��bq\0�8�^�]o<��%��i����.�����g�+o����;��o� ('�_�:Y�+9s.A(���$�d�M?��]պQ��p�	���h��}�8m�,�3㧤�n���]~K莢%����l)����h���s��z���y�Wb���b&�p?��EƏ����-��'�7D�!6�p�`��[ya�s�	�c�M�᫊SDEl�.�YS�rG�_�cZ�u���$��G	�s��)UZF�Oi�$p�Z�|F'(V��f����	�w��to�.P�T �������"r#6�@�n�`��FĮ��W���*aK/�^'p������-�β6ңq9�R4�L��$:r����1���TXi���|;���� �C��л`l�~WYQ��Z4�X"��F"��^���.��Y۞W[���<�r�0B��~vr{<&{�J����Ź��n*��r�F��r}ۘ9��X�  ����r�"t��o�{ ���]����Z�լ�|�|B�?���wo9��k=K�.G��'�!�1v}�j���V݇��Ԛr�{+V���Š�{*�9�B�-�ϻ5�p���=��9��]�$!b����JK�IDLj� i��)�V����� ��&�y_:��̶�bHRz�H��@&m��V&\xZF�X�m�[�F�n$���<�%�
�O�]��u�vN��i\R�v8�_k�JJ�1ȋ2�Q��ݢF�v��+ߎ�"�F]rמ���<G�CL;@�8I^�S��m���Բo(���97Z�U��^5 6S�����%�AҠ�z��;Ԍb���bs�Q��z3�	'î�R�>�$��8�cI�.A�Ik����������,���eX8����/f"�&hvGȸ�:h��!+��CO>J����q��F�UO����׺QO/ۙ�DԠ�πjڠ,����t��ʿ�7{/6t�-�-KF)�x�н�k�O
גL��ʲ8DyQ���u�d���'�$����'8����s� f���>�}���p#]�OۻfZ��Fz�f��@��ԋ�(�i���� ��g��ϳ���t?�(C�HX��ҏp4��A[�7L/��R~@����/%�:��q�Lr��mI����W㟬�U��G�������Z�mob�.�ݧ뇔�"�����,�>�b#��Q�un<K�F$G�!Ղ@G�<&7�����cu�_������Y6�X:������Q��=B�:	�K�(@2�?G}7��C'J������b*��̖�йo�Z3�zJ҆��ժ���n�-?y��g��~������s��v����u���h�����T����ч)�)��J�fY�l�c+��u�@�|3O�{����� ���F3�`�
�xC9]<�+�H��Z]�Y](:d�H��TEO�z�T�@`����"�7>8�ؼ&|�~�� �
I��Cmh1�;3��и�V7��D�F6�jZ������8@��'R"��K�oK[�.�(헕��m>����-��'���9�'�Us$��(����8�t��?Y`yb��))p1�iP� $|�����%�x[B�fj
zV>���-��I|MU����OP�ٞw&
ȋ.M�����N�e�F؅0������8.�á���huRNV{1��_R��C佲��p���K%l�S���e��wCbh�V��-p4����!�=t�����v�M����4�0�����c�[{3�����ՙ�_���4�~9Ç�<����w���Z��z}K%����_|�Z�o����:s>��a�0U�܏����t���C%�h�IbKʧ��lI	V7�m�2���b�*0})~Ya ��1�j</.�X�|>�:+����
kA��Hx��2l��s���8�F)J�< Ɛ�'S��Wi8�P��yFq�Sj�����9q���K 8�3�9>�){�A jH������=�d�6f���������ܮB�:�1o�=�oU�����h�_E<����3L����J������$�N���Oe��}̿-忀�� e�;���I��$�Wt�`1�Z���BG �Jٖ��[)��2�=�݉��	J����|�U���HD4�aA���"[EZ��A���OD��t~�}��.tNj���%	/����(Hh��g��DF�8\��*)*�h�n�e�7�����5���!�mv�n;�
�].*_gh�׮#s0(���7�	x�i��߻[e:q���K���t!j���M҈<��#K�̯�/(�N��Z���nɈ,�*X�6V�[��X4����]r��u��8#2�FC/]�^ܸ����
D#�c�^sj�p�Z��f�q��Z�M ܻ�ڒ����$ �d�t4SVF`Ӡ��~�0_���~l�]�n̉7df��֎{L�\����%�C׾��%
4W耓<�B��gB�:�!�*[�������R�P)�[�p�.4�xߣ�g�;�ح𝳺e������[�1�̘��D5W��L�<��w#V��-n��v�CYg�O����T�P����_Ӻ="#Y(\����s7�{�Y���'��ki'��t����5�q���	���[��U�\���$�Ϗ�����7� Ξ���39L����[�>X?�?���������F����cne��-խ�H ��C��hT��'�J�_�_;qY
����-ne���!���)�����j p�w�q�>���as�R$�K����Np�s���Lh��駌�M�l��|L��I�d��_�W��PbZ��r Smt6	�fTS78��~���w1��"���x AeW��d'K�f 
 NO83=s�ⱓ����T�(��5�X�ў�(Z���^dd���'��J	��{�W'~��g�B�0��Y��n(/�V� ��P#���gv���~6[�1���yO�m��y�|�V?���H���Y=S���8\�f~���C�>�t��7�E?�����PG�i�r�����:�tK�������!1��S{G�
��~1E��O�d�b�G���ku�5� 6�U�Pwj�3&Y��d;�KWn*��2i�YYZ����h�e�T ��.��FJL�k3u��+Pξ�<JC�F�w^�(���7Ϫ�';�S����1O�)��P2��BYh8��鰪Y�pq������U�}�6k��x�8�iU=\lf�����E�4k�a�����J\pYF~�������%b!�M����GYF���Z=z�#�G4�]L�{?}� ��_`������O�.�\ՕA���#��~�S%���I��b?�k���Q�0�s�V<���{�͜���y̷ވ��Ӣ�����t������p+�=I�!2V������M��ɵ�^\�%�-���t�?t�S���1j8��l�szq�M���gOy�+>6�ȹ2	��&iH�5���>]\N�{�E�r�x����P�3b ���M�ִ�S%��B	@�/C^�}�h��l�.8��67�������',16ot�+�(�>���C�թ�(1~�ƥ���-�l���$s�y���0��fi�y��Z�Bn�]h�5w��+qY3�>��KH�ۻo3˭e&3X�j,�P��#e��u��E!�oFG�Ct��<�Q��ńUb�ѐ�|�l�Zؑ*|ʔ���� 2yVuڃ��B�ߖ�3jnJ�{�J���m�Υ߫�zje���5�P|��&����@̶�鋄���b`�ׄ	,:��zq&_�Ò� |8�9��ēN:}h0*TuD��Au����1dD��(�����W8_��}�P�@	�W���x�L�+�
�+Պ��`Ӱ�C��2t7r�H�)I�h�r�)=�F4�u�K�b Ξ�.�^�X~��1!���X���>d+�UP-����4�e�1���u��"�o���}��#8���/��F�D
���+%�J�7G�cA��|�ɚ�	�Uj������
0���2��f���͢k;�v0�9�ɰ�n���l�2p��$��?�Vm��pub��@�-�!���@a��p���L����4c0�Oo!�i��j�3vŝ�]"��#�����#�)�8X���]UP�� �x�0~��t��7ܸ&�b�1���;V&�6l�k�Feu�5�D�q.�����:>��ΰ����}y{e�^�~�V��7�����m%��9�~Ә��9>\y�7i2��Q�	eِ����fC��J�͓�Cri�.��f�,�K�jg�	xv]��x/
��Q!d�!=����BZ�K��7��7��% SL���#���� �mʍ��i���gZ��ku� O
��CrZV����c��:IU�O�%�*s�i�cW��#�O�\�>߯��5uq���'!�
04[�-�'�u��;��b׌y��g���9>U�����p���q��%��#�'@��ʉ�����w��"����DiA��=���f�L��-A��,�����?�G
d==���g�J(�'f� ����>��[�Q������] f.|CH 릍�D�A����d�$��=p�'���)6�}���g�Λ7���Q2�x;	p-��ٵ~?h�JЧH��
K$s%�^��Ѻ�����M�.�3&�O��3n� ~�O:�̪T^��D� �z��kw��07�^�3H�=���1�o5��tn۟�%>.���d�cM��%��&Q.�3' ���t�3$B�D�4��<��LV��p�'RD>���*�H�76���[�-����1�ɔ8-�ȵ��x�ۘR�����Z-#���:q�I?>-��h���]�Ok�F�}���Ф�BZ���9\*?Ӳ�j[L�f2Am]�e��p��Fۑ�i��Lzr��j���L��=N�&酡FL�����YP^��@S��/r�
�yTZq"�� /�MĢbX�uM�M�]��F��*N�SEi������JQ��1��M5Uv��\P�ߞB'��q�dU9_�� jq!�d"3��M�)8GO�pv�,�_��N��,p�b"ͤk!�G"�]�ţ�%؉O�&\����ln-~C�-qUۿ?������-J�x�&�	�K�����6t�ûDMA��B�ؙ�4r�C�Rt�w�J��$�M9��식�-"���r�#�=�ֿ��������2��p�S���J"+(�][��88�8��gd�@j��z��+�`��s�@�w(� �p��E0d������6�(a�Mɪk~��b*�� 6���,�xjo34n���#��)'?�����Z�� pťXJ�)(�a�:����D�_6ZQg�s6�n���s9��m	���<�ҒD	k<�/�20��Q<�:W�.Я�tJd�q��2E�[���zX���d���ai��&�[�&�[��so#������M�2[[X��Xx�H��/���]�}B���� z넝,��{,f��B�Ytp���z��ϕ5���́V�U��2L��h�}��.!Mi����2ا�ܢ�nalIp@����x ���qYk��2X4�5��3�����<����������SeH���t����=�����nz=Z�?��F�UJg[t�h�� �d\dd�vB�X	{U.;���V�T�u�C
��?��,Al��\����J�V����1�!a{{�r��CJ|�y�֎-nTZ��mo#�<�>�n����^�S|d�:b��=$���'�5��9��W�����F�#*�����^�|�3ZE�L_N|�njK���Az�֨*��G��ڧ[�*>����o�E4O�Bz��a�-�V2%#/��mJ�X���c0kkT�Z�I�(m Z��?SלXlunײZt�@k���_���H�7��KC�����==�}�U����jY5����lC�V>ٮ����:-r�Vez��[@�1��}h �i�)�����o_���5n����k�����^��vfP�OA���t&��c�?�ڭ��lޡ�T���;x\�^f��*�T�K�<��k�!y
T�����gH�a��&���15�E��q���Z�����j�8�s�B��/���v)�<�/f��T��������KZ��1�*��7�W�� �9S�T76$��9��u�y
���r2U�\݇��^��4 |Qe�װ=\��_�][X4F'?\�a��7T7St����x�Q:,v�Z�94�6 ��?L3����R!�,\���6�d8�۾iox�����\C�J�ܲHvEt����hi�5y���f	`l)�'�Doa�G1��h8�.�DWi��n�	ٱ���QjH��]�����hZ0E��qN�T���u"�f�e&�߾��I/�1p+�S�Rpf���h>ާ�'!���j.��R$�kXq��n:����,> $������P^Pbw�G��Tݔ�92�1�R+q�������/�ܰ���fS+�\��u2'^�8�A�����}(��K)23;�_`���][JK�<���J�M(�_�I��֑�^�=��21�$���^�KTݔ�y�M�*ڏ��NIm)X���K�3~S7'SYv��c?1𺀷dK��&�f8'�c�����4�u��D��s�@��z�����ʪ�V�R d(�À���%���7�h�3tw1�����en�8���d�w�B����/bb��x�QΔ�g�[����t�Z��EA�g�k��L��a.�g�=�m�l�m�m39�����ۃ3��8���G���=���yU��thƠF�tȹc�Y�p�?g^'k��G�k�ܟ� �y�)��Z6L}�d[��e2:3N�(����Kx.kޕ���UV��`ɥ$�3���?jx�+f��W�5>�&�\⻆�W��j�4 �R���ɿ��@��֮m�/O�Z*y��xp�uk�I5�l��M�_(��2�kU��;
䎼4���?�˷*�"��2Ce�5
ƨ\~�"�w��WU�@W��#p#�!��@ƈ�9���/ M��7;t$J[��:C��ut�,Ϲ�oט�g������C�z�C����	T
{\䅚�b�`�U��I���:B���S�6I���~|�ү�>��I��k��G�V���[<�X?�3W�P�L���@-��0҃Ы ��:ύ�*7m�1�y�,�d3�mn8�pz�e��B�����<�-�F�;1�,�v����Z�"m����s5�������X�_B"M	eÜ���OsT�p�R�	d[�=6]�H��Q��� �/̡��fhA��dҥ�۰�o���z�����>4�/���:�N�;8����5z�[�'ܚ�&ώ�m���v�j'b��AU�Qgopi�#X���~
����'4:6���N�ҡP�D,=��[��U�R�O�[��j�SAE�e�;p��>J��A�Zԡ����yp�ľ���.�]z������M�+S�hkPL�n`~|9>�G/فt�)�]�33�����X�h�fl�'�B�;�I���<()���l>/*�[Th�����;c���f�%��x��Mv�1��0�+vU0��ia��_���~w�
�o�]�LY�ѡun��dܒ"뵗�0��ݳ�
<[݅�s+��[���0�VU����wT�o�߬=A+��*��g��X�C/��S�dW��+�a��Z0�eq)�z��r�ڧ>��\�00w-�a���?��r.mg� ZD0����	�C9�,���e� RH�i�\���\=CHS��AJ6qB){���D:jL�9��Ӡ5���h\��H=C��9��z�/�f��w���٪m����s"���2����s,^�/�O��(�?���d�Ed�aXN�	D�X��-����[A�Q{��EH�,h�B�����@��:��z=�`h�&�����A�,�ov$T�|�2N��B�P6Xo�!�p�W�&5���{�+�V%}���˃lt��\j�HiVK[ic8޹Z�V{6R� �s5'�oi{���HN�V5����蹞�Y�֌˷+s���*4��/u��ǧ�Ό�˙���+�E�������Q�Sɏk=_��E��g�#���9Ic�h�#��� 儵�s�!-��#6���!�h�7��]ef�u6v�[��L :�]6�S$��g>��$��"( 6���n�jn� ��0u���Z�V��Ӻ'F&��xdI��m��]��V`')������gZ���E�7�Xݾ�%T��[�Sj����ͫ�H�u2�h�bC��<��|7�ƵA/��z,���$P��_�!dvxnv��sU��v�-�-���M}�p�w�8���`����r�.�V�A�*�.���3ۻH4M[P��۸�e�Ҫ�t�1D�w�l0'��_��v�읪��(��!c��dZ>�eVcM�4��\]N�C�݆<g�j��Bd1�r���	2����P,�˟O����5ԑ�h�����t��8��
�<�:��3-=����՘�E�a�5��/҆b�u:V��"4n�
��'J�y}���"h�!o6�  >X��KY��S����/3ߛ�������|��a`Gsu���̟�=�V�0q�-�*T�5��o��[?�%�������C �<S�f;g�	wU�ɽ����l��:�zD���F-4l�ј��5�M6�\��J:��=�4_�!,+�Q�a7�n�\�L��á��7�����Ӯ@�8>ȗ�1��:aLҩ�4T;AF���wf��8��\���s�W'uy�<��g��6X2������n�YS��&�'��o�pS$��嫖z/��%��4���K����2]���*�V�ؙ���9"�7� �UC�^��K�D�h�*I�*��u��"�X0��qRC�X��=�>��B��k�ՄL��^��/<�������amԘO� �`�iK��Wvңϐ� 0c-����@Zz���,R�$Ko��	�/=�[��N��9��w����q,w|�ԀN�5�/�Uz��(;����M�~�����b���t�C�ǀ�.�]l�f�O�y��"���@p`|dD�������$�P#����W�;: 
V�g�!���u�~�ڽ���pP�Ȩ�0��p��L�gGx��FD���!��ET{61L+ʂh�t�]\����w�2�b���1�;eTZ�)�{k��2��
��U�$���T�(�~�r^ 	 �O8��1ɩǏ۾�	_��B����Ӌ�i� �����Џ=�;��`��ǳZD��\E�}
p�R��6��1�����od�nL�B5Ou��g�2)z�Y;��k�����epSXs`kYר`�"$Y�%C�s����տ-}[�yQȩ�����@���<&���2���W�E�!B �;Z�Lά�j�]ް��Us�y �O�C�/�-�4{���:�Խ��4�;O`��;�/4SM�>t$}�a��$�j���+�8%��e�z@��U��2l�DA��ս&AE����m;��/Ē�~I
�a�>�ʳP�����֌�����ളv���K\8��&%5��X_��µ���tA{�}�^K��6RҢ���q����y֠�xSǭ5�'�U�oJ&���/��[�����5�CT� �057��x�z{�tz ͞I�c�Hp*	���AN�Ki�;y�S�SVQ�v�A�����%/�Y;Z���E�k����]YR7�嚖�j_�T��ڠ��Ծ	��ٵu}�o�Nu���.og�23'M�I��p�q��tr!�H����̫/�cK���B6�GV�M9� �� #�C_z�-x_�ac�(W�u_�4a���^3�ǡb8p<R�H͜����C}�ol�����yԀ��t��Д��7]>F���Y�B�D��"j_!�e~l�������
�,UEJrBi9ycE��[BY��̑�w����ב����s��JaF�~���+�^Ə6r��YE|�+,Ĥ�G>��u��e�2愪bp��5s�����U��`z�\�|��e�c��3�����a<�}���N٢/���ʿBg��3�GmL'�As$'��q"� ���T��#'��BȞ���5&�L�_�YS�9O %]��l�����;�50� 7Esr*�L�Әp�/��k������q��]���GR��HL+��u�Na%cU����:�f��*he|��3Z���-pȶJE�_���(��B��?�"�����r�\%1�*��z�BW�h�X�"�ő���TvP�i�m-y���L��F��h! ����Ao/}���*u�i¸��Ҥ�ӿ {��RQt�N�I���w	��Xl(�l�xqR}���;Ld��lY~�!,�}�Q&No�]��D��	��z�2������Q3��mD���M<*�9�T��|�uo1��,��N=/+���-L�q����x���b�$��r@�˹�	������u��#��]��$^��_f������]�͕�P��=��<�5�D��紟x֟�b����m�6 �=gv��9`��g�'P���O7U�'A%�A�ܘ��9/�4&��f�1�Ҧ��p�_b=�Dș�K�ǝ��`��ۖO���Kpb�9���c�3ݗZ�u�R;��SKW��v�,�>��vWV����&� �E�m#<���̯�?.��O0HIl쬵���ן�)�uF7�CE��sM֐�,dBҩ�#:�C�=&�&G���7�q[5"�ܒ$�)��u
���MD�,'}���2L�e�a&N����H��n�-�GV=���� 8��Q� j�����Y�����'����� c���E	H�Ǎ$;`���[� ��2�:=%t�l����%ʛ���BӇ�̈.@���P������M�g���C�����T�zˇ���(n�
P��r����[��L��&}2���q	����d}6k'瘿�^.���Yh�r���ᓿ�lx�+j����"�)��l��16�:�0�� .���~	jPOv�0�'J�7����
�_��8n�jv!0R�鲕�#�34��衯<-��E�C���I�Hت����;�NSuV8�������.��B$ׅLΏ�yh�pP��~��$n�3�\Dq�|,t#�d s���)qiIn�����
Y�}U
�J�|D`j�ѐ�N�4��W'%'y=��8�=��] ]W:�~tv��6zvkq ��4�Ț�^���� OK�־v_�h����t.��Q��~v13�b��w���T5ǫ���v�v�T�����G�t��Z;�]�\%F���i4 �S�i_��c��P b��Y��-��|E ,��z³�Y��̋ɷ�^����K{G)���Y&�0�� 
i>���S��2���]�h�\59��|/s�7�W)�4�?؛U�6�K	t����L�E��R\���æ��=dcl�Br�`d�ӫ���D��b)u�3�q���E�b=qʧ��.��bc�i�����#r}�b�{�h؍��!�� m�j� �-������~ �dS����yf Yp�_A�5�R��yQ)�j;E�8�
����I/�d��J�ʗI\��r��h��}4�B�5a{�� 3�����V�z^�o '��h�4KF�kA�*h��Q9��ܓ���ש�ş��2����P����(�3?i��l�IS,R�x�vӞ�0B�G�apd;���h�]����� �-Sdyïz��B\�����K��H������S��Qe'��N�$��C�(HR튾�����ǲl3 k1�|"?�N��I��L�� �}�
��ҵ�T����b-Z��x�?�[���zq  ��c<<��T>t'��6�`@��z�&� ��F�lP<Z٨�M�.ڱS���'2�Uڨ�q�r�޸d�"]G��8s��3F/HR���,�Rb�vT,�̇}H�W��J��._9�G�Gj��bm��0 �"�Y|s�1ưޖ�ld��ߌ����jg���5��	����h$2&�!��=E��啺�y
&�	+��R/�qL�A��D(�W�Ѹo�P��.X�,v���7vb�%5��v�Ɇ71䋱�d��������qlW��OF8�j����$�!X1X5�7A'H��宫B�WmDg~v�D�z��H�	��gǩ�'���JUJK/(�wy]�ެ\@c'K ���N�����+/d�]e�	ȋ�va]�����zd�x���\�v5n��ߎGe,!��Ik��/�Y���8��f�w�B�{�q��ܡ2�K�n�t/���:��68eQݝeWq	O{����jO�s�㡡��I5��m�Ƴ�히�9Ża��
i���3M�����«mc^8dڵ�z��/����n���c�$��_�/�����ۖ>UU�K��/�H;��m���
;s�D��n��n紽���dBg̝���ٿ�{�N�����HvB�����!�C�<� E0��/��g������w���3zo������~�#m��R o�
?�(�a���c�����Ra[�S�R�/�  ����pd�xKR��N D$�ow�A�����sA�'n���6�"��@�y�-��)u5�Y��)�0 >e	����C4�˜�"m����z��8nc@1{���v{�EC���Y��+uD�X���'�F�p�7��H3��K4��Fu��ّ�K�g*hH�]��;��#m���H�g
y'\��_��LkszS?�eq�>������QQ�����n'v��P�K!�M�3��Ck��B4Ȩ�l�Y>5a�g��&���F�,����� =�7],���f���+��w
��Ņ-�9��,�18GO;�u:�ڑx�!�;��0���Ҩ��:St���P���ne�0	��L/���j��ٓ+t+�}V5����,!�9�vX�,��/j�}8�Bz��9�2[;�Đ��{_6�]!�V��[�S��y>�vG|ݖ3����6���w�jw�z�e�%`@����P��q�>i�f�0�$�QT�Ų�x��(���	y:R�ݺ�*nuZ��y��VyT�!1���S�>�(}�T!z�>ўhƃ���.՟Rn?~�FC��~�Q+x[3�r�+[���j�$l�/&����i�S �2�����pa*�Z�W��-����"0y�����y�\�t����5���^9>"�c
��_.��� '��F�ܝ}m���]������E�j�n���Pf�B�7q�ϥ�z�rW1�h¬_�A�g�U��u^�9ھ�닉|�w[�Dd\����,oO��5qKL�4�9O�g�Z)�1���-�eCM��~��o�_��R@#IA����n�	��6�l�����Mn�`�� c��p�R��l'�8m�1l� WT�e���5x��9�����	��o�����y3���L �;�'�S����'�ؖ�v��rZ��B��l����8�O1}!0����vY��c��B�9;�c�|�K1v@r�WHپr��وܠ��*�^��F���P��<���.�ǲ��y��]mfi]� 5�R�'�d��x��U��g�·�����3[�-��'0/��ό>���l_�����.��.�����x>E��	B������b�ۧ8�Ys(��ʱ�`����9tn�����p�)e�O��4�oz��r`�*yfF�>���P���N_Y;��e���C�k�Ә"�q?�f.�b���ߓ����y��I����V�;,# =���<Y~᫿vA$���g�h3�Hњ^���jH\�Gr���q5΋LN5×���Š���)�H�Lm��B'�_��vT�X8�5��T����令v���@v�A	�<����+������ �t8�ZC���+�C�Aϡ�.�HH�Dx����,��S��[�����x~�������C�S�;4���I�Lh��	�z��~u������1P�Q|��Xo�t�-n&� �jb���-���T'O�DHf�'�?�}��U{aA�RRei{0[�G�d0 ��yy��������/�]��>��(cM�e��luN|�k�^?�O?�'�ńZ�Ap�W^8@�嫦8瑩#Bt^��LU�_����n���%��@p�p,�gL�a��l]�����cu�9qP���8��yEB�Ꮅ���az���w�(KͶ��h>�<��M|�=����RC�V��,�� ��Q����Uk�`���T�Lz7BP�֔�.��#��Ss��2,8w��w,�%=Փ�T���e����'��^(	0,��x�
l�}��E8�xg�=�Ƞy�q�dЊ6<���
	��}SF]+��.ks7y�E:ݣ�
��ìXO�BA3^��%�BS2I��
�$�.ĝ�v���u��G_���.���8�ѧ�91���H��y�<��+	�N��8V�M�1��Mr�X ����o� �Y����E�Rp��9�Ac�P���{~���h�:�݆iF�K��O��8u��[��M�	��K)�[ؽW拰��l�{����q��>���c��K°	�VڠM��#�x䍯݋[�'��8	jf�:� �WCݱ�q\�g�p#�R�y~d�M��R#�tV��ac�����yL&��]��n����o�3m�٫6�������Q�ˑ'�~��M#������L� ��'*�V��Bt�qƚZ[�E����e�~�`�k(�=9E�(�8���9]�	t�B�1K#���%?�kla�}v-�e�-ab[L��|�~�3��G�ͅ;��[��l�K�
�zJćA�&���aHy��s�P�O��-X�q�L���;�q�^���Á����v���
�	"��^�'���8Q6�6_ 4#������)1���'j6�c� �z׭���Щ݆�i<�
���D߿�o1ܺӉ'y��b7�AW�G��_�3z>�sՍ���� �%{��!��j�N3�n�k�W+l�>�&DL���U�:�iI�$����?i�[�oKJ�91uk(U�ߡ�k�-�iCgn&b��	� A�r��ñ��%�����<�v0�����.=�W6�c����e�A-�vX-+8�CF*��=�W,I��O�Q�s�h�C-8����"G��Қ���n\1�^�(:gU�9�g��b$���O�bw�
}��y��16�J~`.�Zg�"� t/]}*�3j�s eW�Yr��uXӍ�vф�_l���n]Ձ
P������:�C�/�{�%�6G���T�.�$�^?����k݊AA��w�/`���T>|O��^
v6�qA����e&h��.Pz�<�c�ǉ��z(��j�!��Y�?�W���J��=�\�1�,�-L�~�e���a�������X��i^��U��w�iw0e4r|�]�f��%ͪ��#!K��$7����J����	���}�I/Ͼf:ԬU��q�Žm��v�]�Ze�MQ�c�負��}��bA;X�E�D�VW�y��������R'`�2�lT��㗆����G��1>��Ԁ�����]�
�\�>��sʥ9���>���'"��P'w.��3Q������M�d�:Q�k�5_��������K�u��a�3-��7N���+$���%�ڸ3>��VL�(Kr����CSG���&���XU�"a�`��\nD�\ra�$����<�F�Pf�о9y|́�����\�ͯ����:�z�ob��zݐ��{���7o��0�h@y��a����w[��v��ɴr����^����߁o}ʑ��#\�N�Z7�ϡYE"�@�j���^�51��EҌ�+US: .�r񮐵�?ފ�)�2rĠM�qH��SdI�l�f�����I��P]��ȃi����$+i���D���mZs/k2(�`G�Xt�	8�~tP���"JՏ���_���<�yDr�/Y�C��p:���"H�x��z���>�A���twL�B�h�E����rFG�_�$h���0�����b�U�4�Z�q�� ��"���c:I���ۿi5��,"����F��8:���z��!���T���צ� ,9��׸qsTP/1��;ZϺ�-���W��Ƃ���|@F�^J��|�4�y:��<���\;�ު�:�(����bC��ڧ������Ój!Z|���8�/y�MF'!^a�f2�@�ˢ*��|���!e��|�V�Z"���Lv���T����J��+O�i��:)��C�٢ӿ*V{0Կm{�y"������c0�f& ��u^x��Go	���E�$R��� 
�9�!��w-
2��w"�oߺ�a�|!����*ۑ���TB�>�la�����?�O?k���}C[p�"��顇Mp�	��bc�6[�w-ՆIWߵe�}��(VL˙� vj_c���o�����T�ڇ���)���A<�Q1LV>`�q��������`�J����j3p��������Ӽ�Uj
������.�����:��[-q��_9��A��D̂o��Iw5���q���¿��[
@#��8LSiu
������t�0���lE�e�̰!�v�?�1*
�I��#��c��e�)f�1�<CH��:O����L!a^�tGƂ�P�C�Z����L��~��-������]1&f��Ă^97���*`T�(�.i� �cw���q�^x�a	A�{�@bR,����,�����_���������R�>���W�:ѩMmj��$��^<�\����8�w��tw�ǳ>�⬸i��`H�T��v	@�-���r���\;J����w�ũ/xY<^���t�:�]1����ɞ��;���w��4�N�Hu�-�A��+�|p��Q��'u�n�ˁ֍��Хi���S���`V��<���, T����Z��~��ϳ��v�����������s,
p]�\�Mh��L�YV�R����~qU94�����[�[r����`A���?��)����_�#��@�:T�����������]�o�J��4do& �.�N G+�)���o��䨽Ojrp��?�L<$�i�F��e�����c��1**W�/��CD�Mb(.H��̕��"�$��w�`��qD��{�R��~i�9l���bo%N�Y��ϖY k�̾��`#�fV��h�����h�mn���7��	��9��N������G�q�����jo*y���ݚ3���Xd]z�	_��(�5wG��"$�uL.�M���ЊF�>"q[���%�Ne���z3���]A��:<%��e���g<����j�E�EZy0�6Ñ3�h݌�i;�{�����0�4��e��R���b��96a4u^Mp�c2�n$��N+�¹8�E-��͂aW��[…6ө`��KCJ��'bQeAG����<���{�7s�f����6Q'�P���Φ�Wg�M���+l�3�S�
���V���Xҋ�'F³�Z�`�3�5-�磴W�J�����>���x��Ħ8�����ʚ��?�lªz�$�ʙ��&޺��@@�.n?�tǴ
$&"{'W���.��7��{�s:w���ؤUȈF"e�-��J{J�F�]��hϞ�B���5`�:���9k�A�ۭ�t��]��:d�=��o�T���,zRb�A�����e��G�dpX|N�fG�B	��	�+F��{�Zx����\J2/Xn������o�Э�eI%A�TwsG��v$AW�
���3cY�D9u��k��1����^]���3�F����{��׿֜�޵7Aꢈ�79���fF|	������ O�n�Jr�lEX{���c�E�$�f;�,����^�1;��Z3��r��!��K�����')`�F��tvF�����g�!��)�BE��IO~�h����n|X�j R��h�RQC������Z���;AH�B�dp�7��x��U��t���x$��*���7�̿JQ�Z�EYI�$�T��UN�&uK֑uTI����:9�f|cD�Z!�a�<t땘�I�D;y]v(��Sj8��{U���4!��N�Ƈ�o�K�n2¹�<�f'N�O�?�2cO�����k��W	���EM���T�a(�-94��u�݅^�a�e?�C������!��t�}�E���aR?�(�"ߢb.Q^悵��8]�N����7���ژz�8j��w����S��8;-m���d���i��k}���X/����M#'W���B]�T&�J6�_�S��3��"�2��A���S��tY<r�#g8�̠��*azwg�	K�[�n�Ľ��nӤ���H���Vc���x6l%�cb+,j����d�`������F-�6!c�['����;6Q��wY�����WPm/��4�V���f�	6y���) ��?��.�^J��/��w��W��f茬r%-��B��"4��r����5!�q��Hz׋>�G���~B�y�C�
��+v�9�!�M+�9Chb1�IFF�	rU���41
���7/����	Y1ѓ���3�;Y%w̄�	�I=�fWXB9�<����\lx���Нr�zS�+�)�٩o�m��{]�~�M�æBz ���x�]�O)���Ck�aD2%Q�����?�w���V`չm�ڶ�~k���ѓ�^�����>X�y����|>(��k�׸�Y��(m�����!�ֶ!`�Dˢ�p� �/���Y��|	�i�n�=��A !��}�4��u.����wHȡN9J��6$�O(�c�<n��l��W�,e*-����=ҙ��ъ7�+ch�%��>��'��B2��?<��FE��D�dFp=�G:�Lp�ƈ3�(���p�Y)�x/����d}��a�-VJ���m5�7^��7r�c"���!F��t|1ɉ�G7[(�B�hHٵ3v��e��?x8�N`	��O`�rێ͈Q�i�$N_i���T#Fi*p ���A�"�i�"���P��6 GA�7IǦ�Q���M7�w�I�KW�
^XV�5�|�acK�V�eM�eh$�)v���f?�&�OGn*hq(1���C���q]�ud�
e�݉�j�B-		��-z����>\�3v!xG���3ĺ�msw*�6W����[�N�2�iU���	��Q�9*&Wg��s�N3}蚙��h����V��Qf\�60GFXN��s|`ӵ�
�-����t�q�O<T�6�G��ΈD��,�h�E����4��B	�ի"-��q��%|3�(IX�}ƪ^�}��ǩ|����N:�mk8n!:a\?��s�|?E��� N�.B��δz�ifmbC�qx��PCc�w���ɸWv���QT��V�V�w��qD���B,���˨�9�93.n�/���_µh[��+����Cj/�Ǎ�}
{��5�?«Rc�6�\Wk���y8�Ԩ��A���g�K�اI���v�jG'�	���Y��xTb"i�e��}�� ���/P�gӔ��@��[�����t��D���AG�E���!d�"�d��Z��W�%��_�]7l�b�b�g.��1Q��+��r~>�O����Տ{A&Q�����A�J�`X�]�.�p�:k��Z�D����_��O!t9�1�
�2;tk�k�f��6� S������y�,7L�p6"���y��[��9އ�E	pP�f��$f�^�^2{n}����!sa'Xja�҆���ë�c$a�S/��;�	����rz�!ui�V|D�T����(?J��s��܎0���c����3�=�
���|�(	R�C�~	�q�*��M��w��b�I�$�k���WC�&=q̡� '�e��%!���A��������|�H���K���`f�Z���w�iG'zIJt~*.H�T=���Һ�`�.��Pk�ŠVA'	��ІYM�XIɽ��&�aGWD�moQ���=�Zh7�w���8����K���A`vh����7qU�&��W��6���6γ���.���Z�Q���*&�P��]�2�Y b\�}q�h��>����{��9��WL�8���nF�o��Q� >��#B��9�h�'m㊚����G��S�C��g"�^􁠕�0� ����&C�p�<���E�\T��F�C(�*W@R�s�eԜ�MAcѥ ���� M}s,@	�	�K��z+^�)S���;��������эG��X���wF֠N�%h��%��(p�O�_��R����':[qL��z�<f�����E�*̶ȭ�pi���0t�5�Yv00�z�[�=Z	z�n���L���&@+Wòy��Y��n$�N��S\0ۥ9�W)X�p�QN&�F�}4�2ж�{7k��+��4��<=郂1 ������YL
@"wT��6RdF��,��I6��r�_y;1�=�W��J�<�թ3 A�=��Ꮟ��(��a�!@<���Jm�y���l����x�������b�KR�ą[���'GL�f�$�x�l@���v�r��Y_E���u����v�"��Ei���Q�x��1/��c@31��c�EP������$( Ϊ�'��2)A���q�$$=� QM5����^o��7�(*d�,�t��W�0 z�/Q*M¶�����or�o��J�*'����̏��FS�MI&%�@���u��݂��]�źA]xQMw���/�mmht�ڊR��h[h���� ?In/:�����رl��]�ʦ^�8v��>N�Ll�]���4�|�B�5�M�Ft������`�R��/}}�`=���.z�-��IOeh����i�\�f��?	۷��*���)
�vת�f �s+�sQ�" %̂��I�^��h�/��|CA�U�^�n��:��rx4��)�O�u��]��������?7��F���K7+�I�@��/�ES�� ҽZZ�/D�D��Qؤn�#1��аk���U�@�#�~�x
- � �� �������&��MY�A�X��l�}x��3�T�r+AH����b̐1�B!wObа��=�9%^������1�dͭ��KT�*s�s{�mo�͕�D�]���]��g4A9����2R���U��o�DyG�b��ע^�F_��a��Y�y�`zbZ͍��N�N��wH�_������$� ��㞋�K}C���/�)4DD�j�n��V��!ݏ=� �V���;�PMr�C`=T(
���[_p�:̿|�� ��$���^+>P��D/f4�Q�Ǆ�0���H�Ugb���I!�B3d�����!d0 |Q�Du��J��k[B��F�^D���T'�&�Q�����3�9_��Y6m�V�]�ʖ���������N��<�.�n�a��i�~!����Zxa��l�nۓ�Q�^)!��:�E �"!̿^��BwzL�EΩx��t�i��	7#�@������'a�!V鑗�.1a�����+G�r7��E�{�9œY���'�P�6_d�u���z�Nbt�g��P�y�]U���?q��"�� �>͔?[���Q�ޡ�"�w�;i����n�s x���&֙y��ae\a�	N��:6Q�㩻&4�4���2g���}^��X-|n��1ŧ�Vٕ\�Pը
_�9,r��!gU�M9��Jq�)�����{�8crbN�d�J��'AoN08jk����{Va��R � ���ҍP�5 ������O�5����^N�@Ǌ#L�K�vX@8�Z�#Gs1�7�L���O0P�)B?�f��n}2��J{r��R<�Lr�ɸ��n��n��*U�m����4�ݼa*��7��.���*�ߛ)(���}�s:\�is��Y�+��e��ɠ��L�q>[��%�c�[8�.�P�~���pal9��x���Ž��%4\=����,簉	j��e���,���b ���L���%xt��}x9�ʅW��dk%DB�C�AY�j+�|�'����vϤ��	�pJ")�}�V�*��g�;�d�8�y��P/��~�����ݽl�:Y�1��䅎Ǖa�!t�\W�>�x��,˃�[�o�i���2�G�oF/�:�t�؍��6�C[-� >��<T0�V!����'Ղ��v�B�qQ�A/���f���䑻#�59����j2;Ϳ.�M~u��&3�KC���4�Џ�B�� :�m���yZұz�v��/<Vr��;�9l�t�)�]��{�j�t?I�(�e1�7������zn��� ��6�ç�и5�$�+ٜ=X���h�++j�Ȩsh�����N�E,{L��@x�jԷ'���HEs`��8��Xp�']�t�?q	i�v�Ƣ@��U�AG����u�Wg���p�,��i�[A�0�sws�"�O�zk2~����9=��0
�TW�Omzl�v!I��*�q%7�G���5�.�jiX&�"�⿅Xh�.�?�����|R6;��d�����I�H\3h�Ç2t(� \Ƽ⟝��?'�Ԝ���m}�� '����Y�P�2�p6����Y@�}j��{3�����x<P�|g@��?ͬ��j9��O'V&��[I�á|��P���w��/4�u���-D!Q���m1��Ul�N� g�/��\Fx�L�3�Y;������h�i�5��_<�k���ƈn��(k�m��<}-"i\�n�=��~\м���9�B�p�N�R�3(�7 �5�!��*�� ���Uς^�Uޟbp��~��+b:�C�h�܋�!�iK�� c��A���T����L{�e�е;�j�5����fk�죮e�P���_�3Pp�^S�y�@�m�*C�������j�!��L_�=��e���:�ww|`+�u���r	`1����TU�񟐗߬Lp����/˭����SO �q�rb�F|\-�^қ�hAS�&N86P�6���E��[�.	��rY�g��Z>;E]6^C���ݤ\�T��N�sIoC��}���w��@����h7S���\f`J�q�LM��Qr%8=��E�j��/�p�OO�i Kf\���G�9+� ��HWMDBR����!�����"��~DS�c��L��������T�fvd�D��kv�h����WTp��{�Zk;�����<�`5Հ�ت��&b懻'��C@�Y�`���Ey~*��ǣ��"҆�`�?̓�@�i�c�I(���!d���D�C�d��&	+V�77�d����Ā�>֌���̙]�f��agJ��;��]��.�Ř.�[Eby�u�f���2Oc@�KK5�h���Ϭ��"������s�P<���B�JX�)��UC�p�a�8��o�q0T�Q�I�$5�fM:��y�7Ǯ�s����֢�vosr��J7X���Ǧ��"�Z�`F�|+�7%Hg(�h�8������6+2|�w�:Z�t��?XY��yk�)�^b��r�dRk$GC'YH�	z�hW'Es���\�!�Пm����j7���6�F�CRP�`�w���P�t�@{�0/tK*�*A�Z���9��
�K��\��99�����7Q��#��|)b,X�������G��m��F�M��P��(�c	p�N5D�L*8��h�f�RZ'c� �(�Z ���Cѥ0V!�_����F��D��ĞY��r����b˰8%l;����)u��# ������/^�g}Z�l�7l���(�ۄ��;EWx��~�Z~��s�H4ޭ��qQ���9�kD���D�?����$޿O�a�B�g8�M+��,ɫ�{��o�z��T��W��ni��Ns�ֻ�eܗ{�|�҂S�[1/X�N'�� �-ş��K�[�fnk�Eӧ
�f��n�A}����[w�ά��`��������DCuM+�D�����Kla� ���Z���R��K���9"��Hh����<F�:`�m�F2%Rփ=$fwZ�O���_�O)�ʒ�WL��T�/�r�o�bL4�>'w����c1�1l���[��1$G����6�s�UW�T�5�9�`,Nc<���~��ġ��ic�)�f\4Ǡ�neu�]���?Z�Z��� ��;܋�n�)� 1H"��႐�^�r1��[�TBE}�(��t2�T隹�>��2F8�"�R{�/q���P���8��SA��$J�F��4�y���@�z��_���-��0��/%@�L���q#��8���ϻ��G�33'��v�8���˸��3C�q ����w���U�2
{����S��J��z^�(�~��)�9kk�cG�V��W�#`c�au�s�(���E�7�' t4�����96���c�����d�J,��GȝNs��?���$L�o|+����a#�&��c��b�p��nɻ�����ץK�T�Tɽ�2f��/z�$�I�|F�Nn+�f��@7��h9)!���T:���P8����A%�|��.�9��iR��V��&
w|�&��-�w|B�h�t#v�=ZG͐Y�͛Gq�����+J㋾�
�sr���u�+B"���0)?�����<�n�a�e�����Wx>b����icY7<�����$R����<�� �?��;���?5���$�Ŋ@lA�!��^��|⬊`A^��9|Gp����c�7����R�T_?���"�k����Z���xiI���Ce�J^�{�$� @�t�{��[��b�A)hA .*y��%�:�U�V���U(<��X҉����o�B��u�}@�$�:�z���B��E ��_#�af�����q����*S�6'��]�`��ʙmO��񡊗�oR!��k 3��3">���{�i�Zu����e�G�FϜ�����M\縆�r7����,[9"6ո25$�A��X��I�c@!<�(�쇋�2!����2�3�3w^<P0"�9`�?de��N��<L��Oy1�n��d���� ܘ8�
��2Q�TeJ��8J����dE���jӵ� ����i��y|V/��QJ���E�c"��?�g&���E����1Eֶ{���%,��H⨞=�#�E�{*d���Ah��S8v*�=�X��������R�;l�_ɤ)�O��&|8�`��rbě��.Gi���˝8������d�� B�-0�fB
9^Ζ���)E�D�w�]�;,������j�/���P+ɜ�l9o�1������14`f�q�~��r�V����$�$8��N���Wm�a`�J��)0EAS��5y�6QS<��*]/�ꎵ�$1�h�>`֟P�_��lX�� ����̃��s/}�k �~���l���ޜU�t2O��m���J�w�0|1J���WL�Z?=k䅫��%�?���B�ה���$����L��(�K1���v�Z�X��["?��+������>�C��s#b��;�z����XWW�6p$���ʱ8�������4ƚH��ls�}_i�O�[��l%L�95LY[uIlm>!�¾��|�f2~z��Xo8��a��T����h��D�v>��{N3K2�k�S߹H��k�>��O���?�)O��֯*��|��Jj�7.x+=u�9C�U�4�A��՛��1Oc����|d"�n )��)���O2r�=�m&'3� Iy#N�7P�V[��2���_�,~���G�+vf)륉�4K;��v/����8���S\4��b�Q�WL����)����^�W��~���k4��`��&5���$�l�IH�8�b��?�&5�?z����+���ɓQ���6N�o�������o�e�� Yp*K�j��Y���M�����֚]���C�xw�FM����7�[���K�������^7��Ӌv��u�Qfh*��Sۙt�^~+��P��\��9 '0��J5ѬH	� ��XC�%�*���d-
���w<$� ��H߱)� 9��9C^��sV�UK�`9!1!�v�bƕ���A5�8�ZBZ�n�uܵ�#��3~��s5��N<#�z.���z^s9�ID9�����f>�S�i��(F �ܭ��x�"P&�=�Zi1����)O��n�G;��Xq\�bH�r��{.������F�ioь�n|�"ni�,�T
����^�@�)�3� ?�@�� �C!_�$�F��l�,������|FSkn�-�ǵ�h��}��)�Ny~W����Q���8Rc;���� κGܧ����(��XS�и�-	�.T�����%�+�OKotQrT���'�[��܉i�x�@H�4���>�H��V�Q���c���a��"��T*���Ahh�>��I��h�i�7:>^��n6���5��[�#گq�_��	�U�em�a��άQ���'Vd��!q)�sWCy�<�|rW�{P�9-$,����6�?��^�n^�N�u��&��X2���~���U+u�Nk��@Mf��Z,.���B|��=���m�k`E.A��T��/���(��<�L�Μ��QN�����"ַ�٭�v;�����/��¶�k���c9 h@�JZ��!V�I��f�C+��d5}y��a6D�4.e�#H��_[/d��'�>	�NH[T��	�8�Z���]� ������k�%��D;b�ޕ�����g�pnF�K�; �Яa�IwFiCM�S�VK�����[5{|d�����H Q ����+ܴ؀�`I�u�햰��������u��}����%�����ln1���x��?!�(��О9��{D,5��K�7���"dm��$��p;^�Ǳ%�����0jv_1�'+�&�I[z���=�l'QՇ��C3Ɔ�߂'�j�-}C;[`L���dK#�"L��z�	tݏ�`'F7����֙�I*��Y�h@�/�Ҕ7��P�8�V�Τ��d�9�iAz��2�}V%�LfE!�Sy�Z����X}ʼ,�U�ұU-R�i�hu{f:��^.��~3�{uU��z����q�;I�z:;>�WdI�ߘ�v�/���ZB=��9�,"��9ͻ �?�.���{��s�5q����`l���8�8$f��F��9엮��a��8��C*O�>v
jh� ;ꑚ�K_T�U���rw��P�j1������e����N�0"�1ǛC��~@�]=��6I|U�=�]��M8��큥��?��-���ϾmW��	Aa=m��}��ҧ�ƚr��`w��=�u������_I��v}�L�R��#=�Xk��`z�zm�{��;l��O���D1�{;��ϒ3ֺ��D��n|�&ΝO�r4C}��>��%9��s����d��N��N�����Z1@���1�ko+tck�ّI�!�4=	����{����@!�H��Z�>���Jyÿx�ؚ���L$?8ߦ��+���#���N��zH�!k��ҋz�|�B�hG3'�=y�[D�N`Γ���T@xv@�Ѝ�:��a/�H�u�|^$	���!~$,C�䣡��4�ql�l��@�(��@f3!�G{4}=�<��s����|E�BCr�vJ.2p���N<%�������O�:�z,�&z���Q�N�r�U���߾J�F��Ě��d!�u�+���x��aڽq�H�Io��sR�&��x�LT#�"w�Yƻoo���t����z=&w�o��	*�G�;������^TϏj6OFI�n�]��m]��I0�x=BWW��6�g�qp_��!ڿ/���'���K��y3$��C*ʠv@]��H{�K�~d��t��j���P�*�k���-��WS���"˶�9����-g=�T�qM��;�.)))b����Y2cؙ����^��n�f'�܈�Ϡ���e5��
n�<�T����IaX�������W����`�\M��~�U�(���e��頯(B�K��$�<�ހm������v�x���$2ȫ���s!@��r�]�����ozp0��B�??��I�T�y�-���q�UGhЀL��S�x�PhVcL�Wg��,�U�[�8�}���wj����u#�y�ŵ	NM��̯;g�D�+��������?L`��~�i>ݟ��d��[�]PH�YV�h�
�5�B�%�&������M���� lŤ$��Q����3wq��V�)��nlƀ+�7��Ulϗ�cJKCX2���4�6������=tkr�RGP�$���v��7Z�����f�SQ��
���y�$���z���d)�����JQ���9= ���w�<]@�ܙ��^."��JbD�#i�P|�hn�R�[�Z�	#��
��Z ��,��R.Z��1o���e�B6��ےv3�㣓	lB~	��()�=&=��A5�v�~�k2J�����?KQVU= ����4��SS�)Jvd���O��bY�$@��J��f��Ҧw(��$}bEM��r8b^���{�[��X�����jsQ���Gx�Ɓ�|���,<�3z�G�<��K��ib� ��Е4c�b���m��}�j�X�Vzz,!�"��+��#)F{�T�!B��07�[��%�3�k�w�靈j��>+�4�����%�H�&�_�Du�.g4r��-뎣�Y��4�*�Y$����I�	�m�$Ԝ�� ��Ҏ��cd��i~��B�}�8;3���T�����,�Ó��IP�s��uC��
�^w�m���0������=@_~��~���vO"���h ?�"m����$�A���'L��c�+&{b������srh��ऍs�S��轢��^�Ӣ���@��d��Aك8��G��U\Un�'ISk#�\T�|&B8�������������$_p7��BBRf�V���!������A����%SM�(��]/���Q��+�|�Le�O��G�V�f͈��a��OE�9��yO�2�?A]����ފ�XS/�8���7�C[rC����]�%ěwe+��Z��)!Z��Ey�Ra�����x��=ɭ:������P�{�MF��笔+���̎-��	���KhɈ����vT�4us��?r� �%�RT�r�51'�uW`ˋ"c��B�G����c��"���t�%�7��r������wo���b�@qd�,]��c��i�]��Ҡ؍��ԝO+���Չ5G�"��̬QZ!�@��:����Yt�q#���r�'���τ�7"�c�ò˰�.q�Ԧ"_N8�Y�����J���b�םT���ٯ-�@ۡ2z.�P�'�� aĎxE�as�\(��ƾ��;r�|����SU��k�	��~{F�jr�wF�s��#�m�x��+�z���%j���<�v=X��J�i�4�],U�A@�kL�N�0O^?-��W����̐�z]�vmڪ�NIh��U�Ť4��;��%q�s�#R1�ړ��B#�yrB4Q���ǃ�:>�����Ǝ5�k�_�&Ug&�v-ñ�OHKe:���\� Ci�����ʲ�Br�K��TE0�<kp�g�+bF�5�;�}h~O��]uT�W����|�<|�Ѷ�SH�\��5P�t�)�niUI��w���`�9kۦ�D\}�93�j�,�w�-�j���f�z�!ޱ(� ��u"��}�'�f��c5���׾���'bř]�tVh�����[PC�ߜ��Y�!��ِkZ��H �Fgˑ
�8��U���l��d��gk؝C��gJ��������A�4����%9�T�4����M��if���߆@~���z�2R��P0�*5P(�͋l�*��oe��h�S��jx�=��j�L(|):�Kһ_��/���W�s���	A�a��a% ���N�h�6:cd��Y�)�: 3]S��`����N����r�;YS�с��3MD��V36�֛?y���r��@�t��6.N}��@ʋ����=%��V����QϤ9��A��04��[�~i(��[��13���ʋZ���No�9#�7���Ċ*{N�!��q�_�Lƣ0�� �4܃�����]3>�*�i���S¥Ə7y �2D�]�ZK��� LM��"�ăٱ�� �dʭ��Mi���۳	I" ��ꕻ���W���D�l��{X����A6e��8��a?v�>'�Up�~��Q��Y�ֺ�p��ȇM���tᎻ�z�|�jz�d�9����.*�Ȋ}�PP�_إ}����J������E�!�9�B��O��bo6A�s�o��*�f��q�#��~:V9Ow�ɨX���Op�r	�dr,ߪ�q�Z�gp�9�o�|`��n�~���Ԣ�v������3�y�:��O��Ƕ�#����-���)�mS���~ �ټ8���s7���-��?C5���GtT����I�L�]�^֧ѳ�zY'0���d�`Q��d�5P�$��� iD�U-R{<zxfhͤ����4��'��?��"dC�x(ZqWM9G�nV\�H"2M�Ҩ�)hCQ�_ԣV����K�.���-��skƢ�=j�����rZ��iߓP�4D$���3�R����JW0�E�i�/tv�h����v�&��JZ�=�m�"G7?��Y�K�ȍ܎���PE�e�0h3��`����%����#���5#6�bԯ� �E�z����:~����N#�<ҫ����5�Du�y T�럏���Y�DTM�~�J�,���{\V�&��e<��:����A���q'B��D��E�Kjv&J��髟W�΀��E��������sf�hE��ju����.���y���	T?�8���A��A]_�F�쵳<MG�C�Z2FBG��"����?�C�Wp��K@�@��<ud��!?��n�w6��5R�&[���넜���6��q� �� ��`�5�K��^#��b>���/���h� �;{S��'>�!�9\k13�.�(uY�RM.��=o>�of��������*�{�5��Ƨj,��Fq�¸�BL>�Ry� }A5� ������6h�� ��0��Ȁ�ד���NPyM�c&�K�9a�)��;���3�Z�ls��������mh�z:S�ajNUA��_(*V'�g�U\e�3~(Q7;�'f�����fF��3tH��D1��M�3n�:�4�<�Jl����g�K�@��=�WUK4���v��OՃs'@F~w�t��!s�P�6k]m�����|�Ȱ�r��.���,"ג��T�ޜ}@�B(�V��K��t�&�����,�4D�k�/2�j��2;ES�9��@	P�"J婵@�≎��M���S��J�w�.��̎|����1�x�Ѿ	h!��
��Wŀo��D
棎���ΜSV���4妈]9�Y���*�M���U�2~5���o�{�?S�Aw��7��x�����/P�a��]�����ay	@lЮᅏ-,P�9��J�-^s1�~��bu�((\�r�tbo[�����r�k��.ِ*�#��cW�{L19��7��G���O/lW�2���p���b�W���H�Q-X��NVL��K�7���8�k���k�{����l�i�?�=�9��y���j�Zօ
��H��P����ң�a�
UB�t�k�i�4\��T\M$�ڟWH:��-k�7�D�
�������S�XIW��:7>��;Z�u�-��?�Z��O�0Vm��������gl�zGXWS�J���ZCW�:q,�e0��m*���s��ݣ;+�c+܌4��W�>�����v�8�Yg�H�}��<
@yݵD$tF᜷9B2s�@�eF��1�M��|�/H"%�B�^QOv��e5����W5,lA}�3=�o�@2b��
!k�
�[1�z &�u}���_�1>�C������� pI.���B���|��.19�b�;tKy��Wf�'�G�PoU���\ċ�i=K0�b������˗	sm���H{S�y8Ls�v+X6�A�Y��3"� W������:����{}0��#ky���NJ���ʌ�Y�ձ7�Z)�?-Jy�(����P����>����7	CE����2J���"��Bc6�@�^�;;N5q��4V�݁���`J	q[�����
��؉}��X�>�;=�mc4�a唊�q�aTͻձ	��Dr��� �����嚊��B0>���4�`����92��`q���M#'$1�m]�ǚߛ��,$Ę�񌡈�4�=�cY��NN��Ё�9!�D�K����nV�K� �@�1�0����`��P�3��q�4Ĕ����Щ�X��srT�">������b�	�ϋJ �xV��t+#�a�թ:�$��?O!��A�� �r�lJ_<γ��a��n�f���K�,��2S�3C1�$�?t�M�"��q�!}HZʹ�]ܢ� B
����d�È�c��j��p�mfO�DƊ��$N]�V�w~ގ�+�̦s�\���B�)�2{nW�:�g�	�SN�@�*�&�k���N����10yv�7[&&z�׀�}CS���e­]�u���|��P�Z�֋��C�� ��^��rw2�:��Ϲ?�C�:�3�K�h�}y�*�67�*��-���#JD�u�?1a�}r�#z�RV�`~��&�lȑ���D��I��O8���!��c��� Z�nN�9���'��TA��є����q ]�ʡ��P���b�*J0E4J���²�B��^��?~��u��U�ru	.  ���	��Y�*����.���];��8!XoA�Uqw�_�-����#�!>W:+���=F/���Ĕ��(܀(�4�.PR�F*�;T�]�T��,�lV�	� �м�J�t�� (�5��{�g)Q5D~G�#!�RW�j�Я��������]�Z�-����'L?;�\�ne��c�> %�³�7W��&��|� �?��0�=�h�:+��?;��R��6�q$-���u(!7���eB���Tij[���������hU���ψ�1k�*��@,-�ol���=[��v�ȸ���.XF�/8m�r��n^X�����>��峹r�!s�I�����c��ӅW��}��ﴃ9Z�~��/�<��ڱ�(�y��7����]Y�t�v�䩁AM�m��aV�="��xGW��'A�)
�Ӡ��U��c?�X��;I��"�ՔD0�}�W+͔v0y����.��\噔� ��5x��6���m��IL�k�{�I!�Fh����Z���������D]b��<�(� b�=�F����c*���%�M4�y=��FT��C�iCb<�j<��)�������s���ė��΁��`��8�ʱa��
"�J��*=�[\�/�w0n���ς!���v@��p��S��^bs�!k@��x;9#��A��k�97��5�����	p�����EC5FpDhC�7�+KM�;<��s�?q	���:;�Κ8�m�n�ض��X��{u��)e0+
��%�eO)w�X�����Hд�=��X쯋�%pb7o2�r2JLr���[��! q����/M�ZZ��g�_^'��01�Θ���p�����2>F�e����Sf�6�B���p@Z�i8F�4��=y������O6D��j:�~?*ɗ���d��ؿ �HN��3��aL�S��5ݗ���7ビ��>��	I�������A�3]�.����~SE6�O?T��}��("���;-�C��q�h��g?<�Vx���yq��{m�J&/���%3W����)z�%�	�\,���<`+�T|����/p�WA������/*��5��iS�֗����ڡc�TX��c���dj�&�rj0�cV��K����/
)��r$���;���R�#��ͩ�$[���gխ�����U�2:�v3��a�ݏe�>TC!m�n%�,]�����{>F���xokl�y���e��zJ�H��1�d�Q�%*���pی_�%��8��$&:c�e]��"���*8�6��1��|�sk8���7�1���r!g��CoC���Z6�O�����:��f��M�?ԆX�`���d	�w��E��jP9�B^�~���p.)��J��8la�]��g(}T���;���F�s�V�G�=��r�{%t�S~SL��ί*1*^@g���l��bq2�mPqP�Z(�6 KFS$]�
�ny�>�%��B�xk���?���?�����}�Y�7�����X�瞨D+�|>�toU~:��>��:�f�qΉRAܟ��L!U~�`
�h��h@� Ca}�#��
�=LQRx;=�~�Q-Se�9w���/���a9��Ֆ��8��6���޴$�V�*���K�Xty���b�^�K�u���"���oR�#�����#9Eu�1�ʗ@q	�c�I���%_���6��z������7���[ۗiK�
��͟��sv-�7��i��>j����Ju�-{�z��V�D��(��7����pa�ۂ�K�D�{,5 ��a���;�n~�W�����Bu�]�K��"��l����<�mǱv�)�G��R[rt�c�A!��5�j�c���S��s�[*JNT���C� �e�'��T�&R�Q.Y�����B�@�S�uy�=2�>��û��Y����`�~�-r�y�J�x��7�dGu�8E��tr����2� f�kN{��[{����m��#��4?Ǻ`Yg��]%!��)(�܉q�Q;�DM.�< �y���K�FZɃ�0hB�H��.���Q�d���x�H�P�$C�^f���L��$>;�pТ|���y��@�,A�G:V�rt L�ru��@u�e�NXɡq'>Ü�;�ډ>��'F��o�<xck"­Q������]uc{��TFQ	�c��	�om�f4c�QՀ�� ��������<ql�/���£8lbӓ#�DN�J<��ߝj0��SX>�C��R�X�Os����\ޔ�C(�Ȏ���A #e�Yn�Ȑ`�4F�fw~��%Qx��+�7K ��J�Eos}�Xu��R9R3=�F�����T��0����
'��#�C�������I�Ǘμ"�)����g�D�D8�e)A2y�ףrE�'}�~��h�k��)� �Q_#����Ա&?�k��q�P�WH$�����/�o�T�����%��|����yՇh�o�����&lgǠ��L�s����0c�|@Ⱦ�6�� �bE�	�������Ķ&/�J�R]n��hJ��E�ݼQ[V
$Vp�����ew�9GN��S��w<dJ�F�o@��3 Wc�<��<�̷����J-�IJX޾ڒH����8DH�ۤ^3��IZĔc��L�~��td���Ӊ�]'�f(�
1�p&�����p�4�/���+�����~��zw��)��5i(����� �kj�F����۴��à�Et��{ɉqK�PG00'��lӯ��F���̠���f"��ּ�s�_� *����K��.���G����(��LB1���[���I��U�}�hBAߙ[���H�m�-uȗ爜Y����n�lK��.��ӻ$���i�fV
����w
�L�Qti���A��n8Mw�������K�vfT���)�$c�zw��Vd5-#�����N$ܞb�=s�ˡ/O\����?�p��t���/�R���䔦��TD�AԟkC=�>{n�f8��ہ� �$UG��{�SVp) ��
y�����L��7��{m�_#7\�n�f�-��Û�6�	5ր��Z�}B����1S�-l �)����}Qp�gh��4���.�����>��3�595�0j�O�ߴ�����W:qfU~���d�:-��=����~�Ho���buyy���X0���\MB�>���z驏��Z�ek��Q���|��٪B,�4��{Gp֬���Sa�Cd�v�#��7���ބNS��'���y�,���< �b������a�]4�۰Ѷ�GH��G�U��jVn���+�v�ϴ�	��@Gt�r`��#���ߠ=`��1E�����ӽ_(Ê?}��!��-�}�����:���h��N��\!���#��Re�:��Ա�]�
v�'��ͥ9�ͮ�� ���K������
��}��Q[��*4Mܭ%ŔD�i�U+�)���'e3�/����>�!5X��,�jH`��"���9[�]��x��)P����gO�/�Y��OU�|�gL�A�����%e���T/{���>�����ʒ���4���%���{y��i����,����}[U�>���z���*[da/e�y��n�n\*ǝr��[�m'��n��Kz�&H��DB��=k^����,��.�"�n��F��]�y��M�S�����;o�~w�O�iϚgN�/:Vj�L�Z:y>.Lh��U��L�N�H��;,n�m�KJ���,�x MR���&n��pC���Ľw0k�������Sg+�`�*d���k#o��P�03lɄQ[�$�2�7����;�j�m�a�JL�_�I�N�[� >%�*.�	��$�"Fުm.�!��kV��1
�G��fJ��Sb�,�i�3��]�%�I��M����6eS�n��#F��
<���=�k��M9�"����V|L��#����K$��;]��S�rF�� �ޡt�������(�{<z�1�U��;Q� �*����yp����ю}��ו�]0����� $ ���Xo�d�@ �	���ō�o����Yq��u=�4�ˍ:���3��&�Hi�Y�����a�(#}�>Y��"��un.�z9�ӑ6���5e�����GC*7	��CXSG%>ɞ�Z�WbL�u��ϋآ�����?��F�A�����7��S��=(�ڱ,Q\����I�����?c#�m��H-�%�yx̚����+��#��~�fm�|͵+�%�D��*�V�J�5>����Lj���P�&<k�Q���ZS����l���j�#|�WCq*ؒ�랞�0�\!U�O���f�A0�������t��%��r�kW�|ߜnOʉ�Jp���2ŉF��mc�U����ɤ�:qrhˬr�]җ�a,d�ۃ�B���'�u�<4���%��2��Y�n[��T��e'<�������#h�,���h�~���a�btU����t���������"�R�I��_Z2nr���W���3B�<z�����	yY��_��N)O_Rf��m��Y����iD��e��H���F	}R�����Cph�u\�"�V���[��}�q��ͶN��](y�"�r4������d��hD-��l�VE��	A�t��H{���PhB}X��Y�r- !�E������r����R�����A�7��%뜞�p� Z&$��_CA��s���l$���Բ�D�oc�37���w429u��vk�uUb����Ծ��gގ��F�>9��&���]�#fv0K�8}��SMs|!�����1�㄂u�C�^����>�����"I�*����zAƚaB%�<j0
�4o]�id<���H}� �,��/�����`��G�'#��!6�0��Y樘3���i�65<�|�4��`����Ѩ�R�t>�� �D%��co6B�&��s�4����ZC��oqzf7��U�C�%�䀆����bD��R\�[uv[̍1��UZ��AU�������JI�b���6fV����lkhw�����pΛKl3)������R�ogv��B��ggaX��Uq$Ϟ�`�&�K���-x�]@$����!�����
�ֱ��]���o���羔����80�y�
�&�TW�#Wa;uX'ni�??�SL�:���H��:��}Y�{�%����0�a��ħh�p'=��F��D�2V����.t�T*Ȗ� �P��d�n_A#n͎	_ JK](L{���S �Ү?/%�$Zt�_� ?���/��{z?R=��Ry�>����ͨ�IZZfi���F��,��F%�h���Oŕ��;�+!�q�sH��M.�b]���Uj��2�N��#|���1^$���!g������Ke�?LW��:c�����p��a��N�����yG����&@Towѭn��V'&%���f$�=�+~33�vO�A�os�o21W��p �.�m���&.���O�c���eYŵ�̏�n��mD�[D\�Z�[��L����6�: z_]��Z�ߖ��*��<�"?/����wA��������c��z�gU�ͧ��+Jl���S���-�rc�}�"4�r����Y�|��h*R�-�v�	.���?J�`̣4�|`�<�]!5��#O!T/*3Mr���o�ʊ���N|�%v�~�  驨)��*վxG�&�=&�ԗ���μ56 ��&bS�v�۔'џ��נ�K��׳�Z|�*`�X�d�j� ~�V܅Wh�M������:��xR~y'h��U�w��s>��Ï��N����*��Iii��EW���E�=�B{n�ܵ�c�����0S�@���Q�H�Y���$f�YWL��Q����>�^����L����\�!/zKH��y��ŝo������w��=�7d埤O@
�;CZ#����x��j�'���:@���+)�%�vzAt�Mܴ7� ��[�_�o@2j��b�U��MXL�x�y:�A'�����XQ�yK�Y�}�w�+�+��_�Km�a�ƣ�#��7]턟%�^�M�bD�v�`3��{�\���z��m�Ᏼd�]�(l(�~���/���rd�l��1:��mas	HYC(�Ŝ��/-�������xK`ӈq�ӕlb�o�~e�O�,�q|��g���,���v����$| ?�d𕉲c��f-m��� !F�`��6 f���O�*���Sf!x�/� �� PMѸ'� �j�r�K1�"�5���>-b������Ұ��hƿ�tȘڀϷ@,"���Q�}wDk�#f�z����V	Rm����h���	y���p1��"a�tC����&��)#[gZq�(�:���"l�3=�&�n<���T��Ni�V��ݣD,���Q�LJF��� �CD3e���h��mT,y3�m����`��g�o��YO+�Q�6ٷ�׏Ζiox�����y��u�GZ����*�}���G#��}
�\a�\,�+^_	յ�ƹX�3ԥL������qUq/�ʦ�u�GR��~$�,�O]87�l�o��*[����>�:�OeUzL�ѐ��E������X���q2jI
òl_ׄ��L	e'�|Fa=3�Z�����b�J\�*��-��P7r�z��&̼�6�[���O�!�S�pc��_eh�ͪXbTH��2yK�#Ex�?]��+=�w�;4?P��a�R���/[r��Fl�k�#�H~"v{P���d��������2^���V�o"�A���O����(���X�X�,�>/��
i�N�c&ӊ��S�)��k�3�k�9P/��ĺ�$ʍ�h
̋5�r�v��Qζ��}�V��� ��=߮t�sߎ���9��ս �e'j\��T+J3��J_�;e��ڳ��Q�JH���f��PI0Ҵ|�y#��F��M1骭]d7=���&wc��Ӂۂ��&��a�爓�i�nC�u������&���w����"g/���쐌���o��Ԍ��8!&�+4!�vH�\�f��v��'pJɧ�f���-�$x�������\�4#��XG(��BN	l�N7۶AI�&[)QiGuqK��W�(:�_�������
�g����:���f�����?��Y��+>�ݤ(O�th��?X~V/���p"��*|�Ⱦ\��Ч��4ohޏ]u����b��GA�����u)K�ٸ����5�$G3�ƥw���}k��I�?rп/Yּp�X>*a`/�Gbe�=~R3��k��s-��}�S�k�&��ֵ"�N�Ak��.�U���zw�jL#��5`�� ��lcAiG���~�s���8~^�v�bf=}Sɡ�����d�����t�!�2PDґ}�Hec��(�,&���+�m��$�o�!�Nmɿ)���,Bi/�_�4��ʍ29�x�1��=ʘ23�[��v�F�� ^�Ζ�z�C�T7j���_;���s��a��$T��R�ma�儔а�=Kz�X��	�'xq^�,e:UU���Y��d��4~G���¾��>٤\�5��nH+MJiA0{�@UkvVJ��w��u�D�2,<�����;G�U��:73�"�𿎢��S�b��R�~?'�@�X8w��]�n_�{�2�.u����*,�� �Ǣ��h[�S3�+�
��.�b�W�ԛ���j�	0?jB��V�׳J�Z2�Q���K	�w�<��s�p�&�6e>6X3-,��oG��wIp���`��z����	�,��?[��<�-,���GϹ��^,��v~��@D��)XL�	�������,I{��ы������*�P��(�F�H�Z$��D�s�%9�$��|= ��6���9�!32���CA��Q��
�m��s�|@�tD|j��K�O|���3F��֧H�(e�@�5*��8�N�f}x�������[N�=?f���f�q�ב:
a~�1
c59;�d2�Jd�	="I-�N=3~�%�D��w��/����&�M���[�w���B�&��
Ԍ�d�"�Ux�A�������|	���UYA0�4#�K91��O�d���^�7��w��P�]���&V�C]'�����u�k���|��o��2��N'R1bE��fH�ȀUK�m.�y�3`��Yj'�L�f���d�mB8�j���?��l�K5��l���Ȳ��85J�>60)��h��O�_��ݔ��IV�j�u���}���%�H$�;Z*_đ��Qv��R<��|�9r�=NOD��ڽw3#F���I&sx���Vj�'C^g��fPG��6��z:
���qRQT����cCaDK Җ�7�AO��J�ձfa�,!�����K�z;�i��K�ᱮ�E�D/�S�pȿ��=�I����~��w;bo1*A�.�/�ʋ��İ���CDGC��+���9��O�fo��S^)�S^��	�	���Vc�?:ˇ�M�S5��v��(�O�b[���'T��(%�PpGg(oc��SMԄ5��;}?(]j�z���x��ٙ�c��c�$��jG�ī7�H�Hwɔԅ�$!�Qd��vtԆv؁� QWA�$�z�{/Xl̕`u�˚����a�GTg��oH۰$AeSv�k�{���~l��m7�A2�0W�m�]��E�Z;�a�W�8�� \>����5a���h*��$(�� |w�%ә��/Sւ��tڹ%;
���+[6;=��?	��{�����K�ܬ!��q�ZQ�f�e�롞5��I=�˘�p��r������ﺽ�S������`u%(�%�뮚�Q�ߛVВ�s��8[��HP�FL���7�j�$-��H�!:���b>�XE8���-W5��r��	f�(�~c߻��"{���$�"�2�h�c��\'B���_��P�g�׬A-M������/����t�!Żv�ؿ���Oo4!;J��������m�'�uF�ㆭ%)_ى��L�!�r4����M��a$�"y���q31��'�p�-k�w��G��z���;��=n�[j|\��b�4d�:�h�݉�^���ҟ��Z�)Oł8��mѐ!B�=W���E=d5�3Ӿ�v�@`l�t��=�X�^�;'�(��u�Mu����v^���:+s]��<!s	���uq����4��ך�Y�7d��Sf˖��9�:��~B��ؠy�����)�E��]�<�+�J ���w����0N�v�l���͡���G6]�p��9�j��NX���<�W�����$�
dD�s'Vy�P�g�p"@�u�H�~eܕ6,�y<���$r(�QE��>��k�RS�A��\K6�t0+鿛B�S<7�j����%�Ms.��+פVz�TҠ$����s��S�����ȩ�x1��
��=�L��݆���<,B��)f��f2���8��ת��]VU׽���91^+0����7v�k��R���l��b��W���p��V��v=�f� ��р����ɢHM�ʫ�*Ͱ��Y�8���2���}�f�,�?^�r��bPT���Sj7��u�ə70ձ���ya�N\�?�텹CI�d���U��
��`���:,�>�u�"6࢟<S�r/�l�ω3��k��?o)��{i��l��>���Yf,�����:2Lt]�����i͙�~v��z��>�T� ��/L�$T`f�%��r@�R��W�i�����ڬ�M��l~�.�WIA#�����"��4�d�2[��ɫ��u�7�S��MY�b�7�.�V$�=Jy�F��n|�����k���&mN�Ѡz�~[�4���K�����j��}>��K�O �t����A���%T_n�l��ja���0 G�"�4_'�\�8���:PR4��[������ST�a��@%���оd1���n7Dj3�Ei�'K���O&�?l"�(9�V�neDL������J�6O4������?07��2�O�kRQM��u��o�������;�j/��O!�*�א�I����o��"�JPo����m�Dm9 ���]�6KG�ぞ{�氄ot;t�4�y����y���OG�%�")���S���k넃�� Zӱ�o2�)��a��L��xZ8�M+�����w[��hr�/08��ٶ��`u7af��k����A�.3��.��"�E�rvY��{���c-ZbPB�w��Tb�t��^�f�b��}f���i̓��$3�C&�|�-��C�� ac�5> �����u51��.�O�@�4��Ei*�h  ")��q%pvP�na��1���!��l�B��t8ë\ƺ��\��esЭJ��Zp��I����v�'s�ͭ��FS^oqpR����uh��2_�=��u�W?��rT���[��[���.F�e2�vA���!��Mhly�J��TB�;����I9Ed��0�ϟ�����X�޷��|��~N'XM�7�Tds�I�$}����,͚��Q�$ձlXYm��� �g�T稚�X��wy���Z_$��Dٶ��!v�O�
����M�׈�@_��2�J�o_fk�F��PM �6��.ieԍ�M2o�z$���N�,z��Ey������D-w�`m9L�3ض�_��&eT���|�
�H�Dv8�ʊ���r^���Z%ek���b��p�Vߌ�9a�e6j��m} ��� zbn3Y�BG-� ���\@DU�?0
�1x��_v���R8d��tew�}4�r���ц��2!D4yh�޹a�(���Z��pP�3^��º�O��m|��DF���-߫�<rA��my8X���� � 0�em�5�N�/���0�Z0�4�W�=C����q�
9 �&A����,(��=�V},�j�Qk����W�6/Zއ���7p��{O��Z6�|�+�}a�O�O;�Dಽ
��|�r��Wi�bƭ��P���ҵ=:���b4�Y����vHˏ�_�� ���~�:�d�2dp�e�²:���'�;��xG�/�5w}ɕ�^D?I���}r��zPu}5!p�\�zcz6���
�=�Ȝ��Qp���Gls��^��*<2��n��Y�Ex�JPF�-A�$��c�0��A�2
��+lMŌ �)��H�Υ�����h7��b��^��BɎN��=|�-Pi�|*�$�p�>(��Ma!F�ѕ����|8u��`����ڣa�FCA�m�[Lz:.���U��������>��nSj��x���A�x3Xup��d�͝mUɠm�Mՠ�?�뱫�M�������~x6���p72
�f�/���jXQ��9g�+���p��+x�^����Hw��W9�^p��J��B")��]/�N��l���ZbY����}�2T�^�֘��򓳻^^\� +kfK,8hJ��b���>Gc�~�/�W�
m�n�K���*y�p�l�$2���(1.ܦ"�8˭���N�gc���&�{X��m���)Q� ���Br�,WCʿ/��(�6��{�:�.Q�:?�2śl_d�<9!�)���'I��7·h\�ܤ@�бa�+�d^(6�4EZ��� &�ܢ�P���z��/��Y�~�~�)�[��Ss�mu����A���Z�qSn�Ȯ��?L���|�ή7� mRu2��u)?C��ѣ��D��+{�*��"z�)�΅Pon���*�&��]���7�*}�"1��8PZ�{X��˃Wϋ���6�A��?��C����W;��y�Q�DUl�o���׆�J8�ǽȐw�!��e )���)�v +x��-_)|ѡ���Vh�G�V\���'�=hX�F�"�j����-���kփ���;@>kL��
�G�"�q2�#���([8����+�꯬!O�rx�1$�.i�)��ʧ<x%����`����Eױ �}e*� vʐc����Q��������0��n�X��7ANuD�$/�-�
����Y�������N�
"�nǍ�yj�V���8&�.�zS���.X�B��c�4�����_�z�hN,w7z������=�t��B���G`S}��r�P]��8�؈��w|$��T<M�,7��YW��=Gk�VǏ�$��)x�X#y��v��)���W�j����R�=Q:�eQ�����N>��@�VK�K��`;ly�����;�X�/'E���b$x3������}9�2G��`䶛cny
���~� D�x�NI0�d�}-�6�K0��$R���f'J�? F6��=Q�!������y8���Ҥhd�bo�*o\"/F�B�T�x�`1��'����g>��&��Y�ȳ���& RXe�9�Aω��wG{Q�����:L-�z��:�15c��ɞ�f��3���{������mOkd5��Du��-&�ӛakݺ���ۚ�?/3�7��<Qd���ɀ����	�$�C���l�����3���J�7�� a�
��©=q����D��d�/<�>N���� :�#X7��)�[����(���H�)i�^@�,�u�#�P\�N�����E-j�ɪA �{�7'�u^J�O��I	^��5�_���4�?�؀�=yV���]�+e~�uvH{\� �=�BM�ڐ��yzf����[7_�X���8�	��G��ꂴ�F���$��A��X��NF�5D������o��w:�&E8z��&�L�<z�u��|��8�ﮢ�²�;��<�i+*F��>ϭ ��_{�?8iB�7 ��̬ qEФ`��}!Jp�����ȃ���k�$��:�/⸩]��y3 C$EG��%����:�2f�r�rʇ�,xg(AtI���?	��@6S��
���i��T��MS�׀}L
;�g2�ўtoM��Hh�PP�����x����6���Y�;��+ ��@

mmM��`C��i㳙8ptZ-�x�}?��~1e�vܬi��y
��9�����{�6X��f$�~��8��-�/|z`(	���W�lF`E���S>Xny|YU���*���k�12H��L���J����q�X��+	��ź��Ļ��&��YN>|�	E��*n���NPh�j��9
Ԉ�f�������V��%&T��"�5R_*)�p�	�h.�
h��ķ'L��Gۀ'�^�/]�%+��`4,���-��CO��ލ|6(��@ٙ�8aK�!~Hj1�.ȶ4��r��p�`��+��A��J70�P���?=���%��s��4��S��|],B�/��@�� ��������z�v���T�h�y��c�Ʌ��k#��s�U8 ǵ����H��݇x�9]ѹ�˃�F7�����	_՞���e�1��d�+;�v"���k�Bj�O���c��%{3q2��3w�4���R��1&T<]����&:��䐉��9�����]��w���34z*����^ ����h�T:S��֞�]�L���KOM��M"�P�ebLf	+�x�p��~�,(��Wā#�£z�=��A����&0��6�����5%[cu���Gyi3 ����{�t���u&J4'P��3j�T`���BH���r�0&�]�n�8V�N���$��-��]G?Ǘ���h��X���JΑ]޵'�M�q>�0W���]�-��#����$q���A&	��a#o�<��k4� V�<�͚�#��jt�'��!���� b�i#�ͪ��H�!e=T�	O!Ջ�E�bp(��e"�W�7{�� 8U���mY�gANO<[?MK@����ȿd�rՃ3u�G:�]�2�	"����^��qt�%껌h�Iv�)��~:M���Qb0�N�����v;H�����ByF�&:�OS��e`E��Y|e�;���r��'��V=[��ę���4�6��6�k�ū�²���
�j����ݔQo�YCd݅F�.���2���ۥ�IۛDq�]	x
��pK���a�V�M�W��M-��(�U��ɓCҗ�i�h4�PK'=u�m�9���;������Q����JjQ�l�螕Pl�t��=P@���#$�ϗ�i?�aY��ڪK1|Fl�^�����Eܶ�I�6/3�og��㬜E�n%���Gv�qsT��@-�Pp+��4Ag+R��d�rT�cz�L9_���f肨�v`��N��i��W�/��|��_���K�a�T|�^�6�����p��`zW������+V��-�ї�y�Sȹ�����d�h�7!ޢ`��Ƶ�(RhyF7r7��._>�u����G��!wy�^��4Y8iT����ӗe�H�}dG�{���%�6[�
`wu�o� ����px6�\(�¯��x2�
�F^V�����@�Vv<��֒h[�0<������!�+�#"�U����V���@�t/�5���3�����Z���{�*�BH�@&�?C�! �nв�)$��&���ߋ��-�8,�<���͉��� �Q����<Si'�yW���+�E�ю���$bs=��'5}m����LPD����$����Us]"D��-�����P��+�R����fON0ϕ+��q��*ΑI�FiU6�A���s��&��%���y��y�Ԓ�O�Bw�fu�t���9×�ch<��fL��T��=] p����1R�=~�	:��6#�3��|���]����#�b�c'ib�GY���N�_::)��n7�lܝ�+<���`;q���(��lڝ���D��[i^���F��T��T���@jGP��)(����@��Ä߿�1�ߔ(�A��W8c&Q�%�$�߆4���W���*ѕ�F�Oq\
���Lp���t{�4PCf�Ǥ���w��$�F�Oü����e�%��U���T�wg�唊T�+j	�@FW2
���ɓ�L���H�(�L>:��`w�+4���C��E���u�6Cm����Y�B0+�KQG8�9�=����2� 9��C`���4=�Ϫ�o���O���,�<�ٝ�e/�J?J-�����  ��e��4�_�gaN�ݕ��xN|��N�����A�,ļ}A����fvݔ �ڈ�WX����\3<������3���Fb.�&����]�u�X��:!Ñ�x�bJ"��Cf�-j��,��2;0H�s(@ ��:%�A���-p	�lMp6�����h4��؜B�,�h�k�i%����j��7d��Q749n`�qx�$�YM��	��\����h�x����xT���5��5U�E����-Y�Z>4�R^ ��s�������!G�%��U�����+��q���G�z�]ԍPq��'n$��&���v,��dX��l����тMh��n@Ç��:_�$�>���C�\!����@�e��'�I+sS�g)�ԅ�_"�}�h_��'D��GA:�nBE�S�-GDj��vKٵ1x�	a��6���?�[��
�����x�;�cV��c7��IY�����hƏ��� ��Ϭ��ϊ_B��b�l$S̝�vH��+틴��LG``�t|��fQ�3�����5�Ǖ?�;�j6�XTN�=�<,0�^C�vw�aƩ����*I˜��uRr#�r�|��KF7���e�p���%jp������R��-W��~#��{f��;��=����z��|�HSEh�ߦ5��c�y]7�8���,(Wb:��!UjKW<Ǎ��L_������� �cA�?���j�p���6g���������ٚ�H���OV�U���[�E�&��^�٪T��Þ�"Xa����ă�#J�f5��T��O1�	����>�R��[�r2����igܷ{$�Y=y�m���C�)���Wk�����	����>�T�6��5�)|c�@1�wbg��5��P��M�&��1���Pg!� r8?�o1��>�-��8�#�!�Ř��w�^��cÞ�%3�ȴ@p9/�i4�&�h�AVo�����r"�m��[R ����N�߭�B�@j�y24n-t�zw�Iun��.�t���$��:�?�f� j�z�^<�jچ��F����攔��h��#��u®�,�nNU௮p�'IOS($�0ӽ�c�I���|�4h�
 �F�C��ڛ�D[`�i2ΗN3Zg]�ߢ �B�����LO��[����Re9���ye^�ch�+��a�H�3\��}S���R�=�����O�O��'E<3gҌU�3�RY����k��u�h"���L�)�i��K�d���	B/���7��F짠�+���������z���bh��h"g��EX�`�� �P~�)�UO&��:��J�G����Ym]'�H'A{6�����+A�I�7_Z���M�6܅�Iwf~sk�3�x�HX!���Ձ���+��|�&W]�+9O��5�?kP4��!���w"r�}ڣ��վ�'�O�+��@3�.b�S���#�?E�U$o}a�Ƞ�haK�|�e1*������3 ���K��u�T��V#Qa�t�
[/EY���3�=gd�g�9h+�zժ��/�l��(W���qȚ��ױ:
�-��'�@����Ro"՛�,կT��B�B���:��d�$_�O�lTc�*����H���D�ͣ���D�%�=��_O�|9�)�Y	-o�u#�Wd���(��e�'���>�'0!?�>=bâ��y��DYtF�ۃX��-SZ2Ͱ�X�+-h{8����>�;��?�3t�9�_�DC ���řt�F�v�9�h]�t����J���J�հ�<7�>(6�<�1y�nkMv+�I�
����J�  j4	E-~ʠڍÛ�J�ub�y��$�d`��Dǆ�Z���$��k�&3j���pC�ן��S�q$W�acJ��p�� ���My�u��=-MA��[���kZ{�Gi�5'����rx(,IT,c��Ҷ�R���@vxG�i�;Gu�I��U-�*ߵ���A�w�
�ճe�SZ>Q�a�z��)��CƓ\������q�v�c��!������Z�zu0[+(�^0$�*յ� 'bѫ�2):���5?�{ܤ���r�p��� ~jf��'g^�c�v%�L։�\02�t�θ�i�X��<k��\#j즹� E�;���]��k���Ċ#��4��V�Wf��I���F�k�l�\L�-U	�P6e�\@)pk8�޼3H��Y�Dti��2�'�yr���!���d,�^a�Y�Y�	+As�1v�3e����@>�W��<Fȯ��s��E��B~`?(-�!�m�f/��.1�IM�&_ �oH��߼u��"q�ᇕ	:2�H����0�9BG��Ǫ��m�s��Haq��&;�!� EP��YfIp�!���2^ '���Z%DTO�+Q��"R1�������gh�yy�d!(�y]�v}����(L��Q�<�ߌ�LR�Xگ+�M��s���
|ˋ�����嬢K�4�� }�uX�~0��!f�|[2�$-5����0�/���)��4�q�푄���9�\7�g�l�����}�϶a��R�a§��/:$�I�]X[Z��5�eYısrN؞Ae��G�^��&��^��7{ �|!��Y%����80L�4;Uq�!�]|~��`������I\Y� J�oL|*R����S���k�u����t�w��n�*-�T�1�		EҚ��=���Yq����z���<��T���^^x���
Y��#��DD6ߩyW	�
���
;�O�YYq&؀!�?����1`c��/kb�Dס�`)�6�lM8ިs�'m2�h;�!����}�]jc����2���wk��3_+�.�2�0�7���y@P�EP��3ג38ȞC9��f)ط���ϛ��}��]�(�S2����Վ4;@�=�獌Wb27i�Q���JF������Hܻ��݇a��y	\�ŇfZ�]����X�;�)���<	E��6��Gᢪܒ^��<,#yZ[o޷;��(Mfn���r�py�Ns����7�3�ą@�J�l_Ù|�~ީ��}��כn@��|l��}A��YY�r�zh��Q>��C��l����%�@2>�~vb�=���}D�S��=���*+v�#}aD��t,���� ��H��O��0g�*��Z�Q"�s,�ǜ�*�D'qW�ʱ~�$�䀨?w�ٶ߽�/��:uo >��4��>wh0s֟,�,n��;@���/yBrʹ��r���_���{��*��o��(eR��	����l���J�ِy��[����:VQ[d�]�cĸ!2�xmӼ��%n��bTr?O��Cyˍh3���|���o�	�3�<Q,�� �(��2�A�aiC��� ��w�Ij�zZb��{��1��CB��	tj2^��"�|G&\�F��h���O]Z�=c��^�V������O�H�CQ8�j�H���c���E�_���7����S��vb���(��0$�D�͓iVo�x�DTl6�[9һ�8��i�a�s�U/V��S{_���E�Pt̫]�>��ɚXB���z�Ȣ� �`��U� �)�c���d����}x���ɋ 	��4�9L�=O��y�{�ѯ��$����v�Q���_-�T�tT�i��ӈ�:��%M*{]��ïӝ�iPc���S3�yc?dɰ�p\<Uq���[��+����LV�5ħ�s���" �^G=H���bp�3��]�
�Z�c[�̫���|a�j3/!�>�)P�,�����3
��h�>��'�G��` ��c��w�{����*(-��t�>"��<l�/
�#����s,�`�!jt����Z�Xtrl1��8ހQ��/��z�h�L���W�H\�y�Js��%��Ӿ�u,x����������h|�4`��fڵ=����Ԏ&��n�(<-���Hn͗*6ܡ�p��K�[�: fQ�2��#��4-�4�f����vu�If\W�[=��tx��r��2(*��}�~�_J,L�4M���ȫ�Ot���e�rp_#7��+KojSS(�{o�Դ���8�< y���k^�4�k	��ʟc�%T�&����j����;EXժ����?I3�u���{�X��/��N�G�,`����7��� ��񷕆�bY�O(a�PϚN��oZM�b�XYQ;:סRb��,���Hۍ#�7G�T��������j�E�i�.j�_�Ռv��]�v}��lVc�'�B.�}%��"�{�?\3�I?y�_@�/=����K u50f������w��Q�^���������Z�ʾ�	C�r6�6�URN�nT��N����ࠚ~2��`h��~����:�N5��
~�k����z���Dn/L#w�t!$g�Ɂ�oy�x���%AbA�ф����dJA�d.�g�)��a�����N,
�������\"tj9�+a)-G&\`���c}�
l��X�Єv����Vy�B�e��'����pS%�]�)z�+�:t}*�۫B`I6h���s��^�/�mؼ*t�?�g�U���\{B�&|b��R��i%ϩt��p����Cl� �;�Ҹ�A�dr�,OYD<�3�}1�5�G�à��Yo���j�a���FI��d%�5��E4�u?���\^� ާI0�K���[.���������g�o�I�B-�껰Z���6mmHa=m��R�l>���J����t܄X�����y�xǊ�bH0e|�=�4}��x�,��(]����� $�H%�d�V��{��ΐ���@��J{Hr:9���6$�+����M���X��~�4G�7�o^m�\"��|�U����.���`�j
 YU���߮C$��H�˪��#;60c
=�.��,���U��?[B��l5�ͰU+����j z����	$��$�Q�H������8R�r%�v����0=�������x�E�e�9D$���F��Y��A����O��a/=s���;�x7�|���v��v������TkuQQn����o)2���LM�o��U5��e^|����O�;
b �~����0��Ֆ(DkP�����ԭ��}?l��j;/�-����X=�yQ��2�M���M'���i{�;F-V؈>��~�Z-�.�-\�l)��:|6r�I� )ӷ4�I'�>����/�	�sg�BQ�\%+�<���b��7 8�)8��s�J���c�ǀ��8!��}� u��ϐt�.��=��v�u�K��q�����3a�<{WQY7NxB���넔ܰ
c#�n |[/�Uo����`�E��)�1��]���x�7��U�%<��uη��Ē��ʝVJE
�d�����\-0�?�{s����A_����#۶�
��oZ�/�!f � :�2�nt�'IWy0���h��[�< [�@4c��F���ة:�e�9�?Y� t��aI���Zݰ�an��k���SC~(]�7I�pBh�(�g��	��c��),���u���8d@\��I ߓ��)!S��EQDa��Y��џד��ѕ��8NP��x�M}v�C�2��qN��7�K���[�s���p�0@�t�=�_��b��`jv�c��g0fmoR��t��E/DfGl :��g3�6�JH�vf�9k�d��#T��z���������Maԡ)J�d.���6x�8ko��}q�k�@sL���|�R����9l�(.�|1[YZ_Y��?��_򳺥�����������gPa�k�q�������茞��ݟYG��G�=� ��:���MH�
��y;�(�&^���>��^z01=�ɢ���b�� P8C��<�-��܎F� ����T˄{�c����e�5U��	udH����xRښ�*HG�qY[�-��ؿ�NJ���M�{�d8X�v�E%�(6x�vzd�z�����d�b-�p�$��VtV�e�\{�m�[�G��T{�?����6��Ky�P�G�1��sQ��;�,��4`�Կ�v�'#}/�?�Vc`#:�O:+C��Q bʖ��݅���͓�6��R��πH>A'	�U_e��u2�(H���ț����]�����x�F�g~E�ʸd=aى�@5��5b���������pa�����Sԙ���q��WC@Yk�j�R���I5a(�Z�:��[�|g��g<�Y�}4�����zS(���ߺ-�ϝd`���+�:;��2|�l���hf��8�-1Ѕ�lm�g���N�X�qMtat?����:����)�%�A(w��-�S{:P�����`$?k�Yk�><��Fƿ��Qid��9ғ6Aa�+���"v�u.����d�n���Z��s)�
�x�~4��/hMu����kyrJ�Ĺ��`���5����/&G�>����mH�Yp|�yȃ�֔:5jR+�"�:�k�SV*��'�h�VV�u�b���{���o�@R�x¡N��b���".[���1��T�_��,.���OS��U��=��O�OP�����	��iM,�(
3��77�G�dE�:���zPv����3�.�>�=����<\'�n�Ϥ6?�sӠ"m:��L�Ԥ ��|��#J��)Nk�£L�W���>I���Z�˦B�����os��Rd������mqP�0�N�F}̸�W�l��_L�*��w���R�V�v{�c�\ބ~ A5uh�P���}����zE��X�J�qN?#o�Ј�b^�1�4̴h��-�y���C���g���x�>���ՁW�@�.��d aq��cT�8�@����`bQ9��n����){�Uv��f�?p��M?�D
� d��;�^11cc����2�{�NӋ����À�_�<=���7q�BY���8??7-�Q?��w9����Dj�yT����;Y�8�);�N}|w�����݀��_�5�,͑��J�ΘD�>�ӶϮ�:Dx_���!��`��t���>�4��FҐ���.A�	����e�qIQ7F|�Am��Mb��:!Ĝ���h��g�{����,��3F@�߹�8l�} D���])�V���e�!���-���c`���Rۚ���%�B�R[8 �pp"�Ċ�c�M=����Ԥ�>�K�^�]���s.@�8q�.�Q� V
�`)�$*f��&&���b!�$�߷fe��'�s3��Hj�p,�o���7��u\�������#��گFv,�ҥ����)ZU��d�������67�e
�E�Z0�B?<�a��QX{���RC�U��$C�~ҟԈep���6�"L�:)SL�(r�<����\ٛ��A���y��ڴ4�%�@D�P'���i�jq��EFK�>&#��A��<�.��K�yuח�y$�a¦p�N<��7����O"���`܉�s 
�/:��{+V/�Ht��y�>j�G�M)�_,;���A�쁡y��I�D����d$*!��!݄<��=,vs�Y�?8��O[b�Tq�+�o�}�Ns�20k�R�5��б^���?�m^�9Α���ش^�&���nÀ>yw��y��� ؞o�x܀ѨRq��d'��sߥ����ⅰ���):�G� �\B�a^�T���m2��k�Ho���P@j檡����\Mͳ�;�7��Q^O$\�|J.߁
6���aeQ��3�gi,ɽ	=����%5V��R��ڦ��a3UY�J�sp��q����$�ǒi�@qO\tȻH��T�<ߢRO�*�n�W?b����Y>�{b�M���Ɠ�>ak2J<z�Uw�l'���_�x�l`Y�S�㉢�14�HؓW��v��(�w.b�'7���-u�^)lGo�j�7Ȋ�)7Ň��y����~C�����}q}47��2=����Wg�!qxG��l��$�=��C�G�����@�[k?fjM�\�9�l*�T/�>>	��x�y������w$�d�^�����Cc�V`����3��w:����-�?xt�"�j6�����!��m[aZ���v����Й���bbx�y��,Ϯ��F�����f� h)5�9�!mBP�ɉ�Uɨ!I����,$�u.%������Lo>4��,Ӕ4>WH*�^:�c�a��g�&��?E����hR�p]����ؓO�1��@�j.|�l�=���(���U�d`�@Agъ6��+h�g�ܡ��L�e�X�3�^+{�ߓQ��d�(��X׊���p�7��t\m9��qBM�r0�7�Rb�~��o�&��諔@�{��f0��l�����9����1�2:_d;�5�"�,X0a@���U�����#�T�p�Vq1��v�Ia�ʌshP�&�ǧ&�pGNی���Y���F3'�9Ǫl� ĭn��	9���]�Y��W���4���~�X#���݂LM�L�/����h��٦�ܪ<���C�mq��FeJ@�WYx���B�'�������*-����Q���� н�����T����*ǽp������/�n�dw�-#F�0����ƖįP����ù�V�l����<C~���,�s)P��2���N�߈3I����V\�K�%d�d7��x_y$����H�c�a�ƊkWa|u�\x�R�3_���h�����驼��F)���m*���<$�/�m2�\"`9D~ cX���
��G_�+�4㙶|�&����Hc� �����m{�l�b\8KƑ)A%�4�y�/��P:C��Q6d��µ՟z��ϸ�2�~Bӗ}�~�T١�*k�Րu@w^���S_eݘ:�T�?[��J��Q?����wo����f�ewe3�HkB�C�2Ax�2�̠��-A)��,\�� xD�_�2c���7�o߿�%;��Q} ��J�t�T�_��b!��2{Qx�F
�k��$�l��:�iB��ү�H�����vN!��B �(����t�k����x����r(1?�},��Uj���K#��0��$O$�ȏ�D�)hD�A�a��p�^��O�t�Ȣ�n<<���J�k)�Sm�������,��[l�S�l��C�`Ȣ�Nd����J.��f�z�lO��VH_%�=<�Ѧ1b�u6�3�_9�f�2�@����6���nI��m\�*�wI�1��]�*�B�,�d�yU�<]r��2@Ov+ ؒ+Hp����K3]��;v]��4-�����[SH|'ҍL�:~=�c:�K~�����:6��$��r��T�5*���lx�v��$��?�9a��x���>����pw�����d�?�iiN)�F��5��G�`>uڥ��.�sԁ���zt�J4�{�&���8	A��b�L�|�S�υP�e�����N�X��<aHn��5X�s����o�Y�_�M�		��|�$%Y8�N?b�_U�F!_u��ĵ*���/��n'���M]=as�3YN��e/�J��Rv��K�'r��r�I��K]���Ub��:�\�2���h��F�M����{~�p�L3�E�9D7?1g�A�����he�Mb�l���^�&]��r4R;����
��觊�"��fz%c����L�e���K�?�[����=��.q�]5�}`e��KS`P� �z�w���lҮ�U�n�~���<�$�"y��.ғ��6y���"w_!���W$t;����i��h���G�Y�Q ����o�Ҽ%�����"cC�1
�
˷�w��1������*��X�?�gp�ǆkl�]V[��A|`�Ӻ�sf������E�cpƛ{	�#Il�!��(��\E\�m�D��q<�}�e����Вܿ���J(���c��
�����n>��]�1�Š�
�n�wz�Rʫ?@��\W_�q��d��/������}�a�j)�+�PP����n��T�k�z���D�@�Ѥ�C����4V|nNG�W�QL��GGWC�keE����L�;��uZr�����Q���Ն�U���|/k�e{�����@A`p���~�iݏ���6�����S0�iZ���l��Ƈ��0�>j�����L�� �.���AX]�d�)6fHo�����'MtSt]i��@��9��[��_V���-,��E	�A�5釢F�[� �َ=)|�/�6?�7��y+o�gH���!��6CE�Ⱦuu$M[4�2�$f�����mK�,A[%��9�@�ʊ+��ezH���'���YVf�t�=T�۴�����(<�i��*�\�~����%뒗�9,������X���ZF��LC|�MI���Պ#L����L��7c�(�Y�"��\�7�����F���h��1�8���t�T�X
"��랶�b;z�P�%�Vy�2�6Xt�[K���s�FV��HvS���jN�]��8�0i��nۘ�sP-��b���B���l�����G�po��y�d��A
�t�J7=��^��7�o��f:0TV&�K��с�=�SU�U�Cd��ig���E:M{wS�@A�&�{�x�*�"��4A�Ck�2.{�ME�O�ģ�4c^�z�����>��pU�Oe�c&
��I����Y%m�V D�o+�,��/��� �Yd#��u�6��c6?��؛� W��B��x��B8����_1����T"�'x`�{��d�0�g��W�2��� ������h>׻~-�}�ҧFUiG_�ӬL��G	$����H�SZO�Wi�mq"J��9ya�,��A��@e�y�/<D��1�t�x���/�R�ɘ��0��y@�>�/����Iv�$4�#I5�xZ7�?�@w�c��U���g��l����w6�����k���ņѩ�78�c�l1�J/��õ��I�~?	�dj�����R�y(Zf��ICƷUڪ= ���_�
vRYo%���ew9h�j������]v��5��"�-5�����²��@��J{��۞��,�e�:g��-o�~�J	�!c�����龍�y�6��|�g���M�-8e&Gv���� P��؎|a�(Fͭ��R�}:!t8PYÎ-j�(�u���Gr7k�_���g2�q����b����121��@0��H̪�C��2��d��ן�E�%*��WL��7y.��V�sbdǷ���pS�i�p�/Đ�T�~ڔAF%�Mi� ���{�uV!e��m�j�F;�
B;��G�X��ԯ������b��%32w'�ƫ�Цt���t�#����B��׀P���i?w�:ԀaȾɌ'	)��6x� ��F��Ӡ]��lx��+L�ӻ�8���F�u��������?�N��rv$eS��~���A�z[���5��t���پ�\2Tz|'g��Y��;7�9��+�&-�t����xa�ͫ�_�'F`&KY>��p��̎�B��x���úH.Fw��7(O�(�pԋ �+6����nIB���H�h���F�TK��ʳ�y��qP��_&�ʏޫ P����!���!4mol�+z���;
�z���t�aPҟ;����x�2Qz��vNp��=�{����۬�#�U�n�Eenڴ��l��Q>c����	�IB��~��+ρ��o=��UX���}�t�r���i��e;1�c�������A%3B�"��fC�����pgB�E;���U�7�Π��c"�<�7y �/�9+��5�+���afy�KJ1x�^"�eE��L7�]�/q(��'6��L��4���
1�"�B���(O��sM��C[�K�����G�Ĝ�<KE[�ӝ'W����YW�/!z� �>
ST>P���^� ��\��b����S�or#-�;dH��Z��*B_zo|H�����2���6��J�Y)]P�;G���	���=v"hD[Vb�w<(�6�n=V[��8ј�G��cm�AaEZ�b%����!M�Em}����"l�9��:l�<���
������f��(�hK��� �q�mD^c���*�g�`y=(Q&���plڌtK�cq�dӨ.T�1R�T��O;C��t�p��|��w��5Z���HjM��:�Kz������nb�VH��ƎDߋ�EE�xذi70��ev�^ÑzU�u^��n3���ǌ֓��n���P�ܕ����57|*?��]��uŜ$u��8�?*���֘Ǳ��j�+�[6D�]nJ`?���Ipq�Pe���H���{G�C��Z~L���M�[���K�µ/�rbP6� �淋��uyȚ̿�&5#�T�D\�r��b�n�i. C�EE�3�}���m�T�!�K���L
A�����v	��
;?=��1�����9���(�Z�κ"BF_�KŒ�қ�iIb�!�ln�"��jL����*�E�/PU_��IPa��	�!w��\�'��3�S�byuoP(�9SLű��n=��t�I���i� N�>���RB|x4��N��V�YQ����ZS�.f+��IG-���[�ӕ��j���o.hM�cQL]���a#�=����ܻ..��L��J��b!.��ךr�bp�5*5�����kGB�-���n���5-R�qd��ʉ��'��Z*3��@5�ԥπ��)i�=��v*y��(]���6f�����xC��\� �9/m�ǐğ�����j<ܸ���ح��ҍ*l>����>�@L/�$ʶ�Ѫ}Ô="�1��6ښ�B�f�)�^�fl�d�c��z<�b8��
#�{��E"7$��αF0Y[��&v��vH����@��P�w��Ȇ��̬pq�w�'�<���	D�W�E����J)_I���mp�N�(��܄\�� �@�yg�f�j2��g:q�y�$���0��J�H��-cN���1a@��uEe$&A�%��h��S ���ѿj1��Y���)����h9vK�=��w�rb����x�!�Q�W��d�".|�ɸ !��z-��L���0��Ut[n&j-i�U���oᙙ�  3W��(��,Qv�?�g�tLj��a�GR��-��7��f��<b3�:�����]c���/-�@0�P�R\�l�r���j�]�5 �lx�9���fGi/]�\�
�-�ck^qWE<s����$�HPe�A��C��}�q�:�%����*����� �Ƹ�]����p�l�9Oa��6�F�T�%�=�y���}��i[r`��l�U����K斿8X�^?}#5`�P�9_g"I��B��a������V1��3�Ƀ���=�R�	�D�Ӧ*Ih��X'�y;|iy��9�/�c+�؀��������=����~��|R?���b�΁�S�3ϸq�J��	G�PFa�k����󫗱7A8�s��}ɀ�6*�_9��������b�6�!�j���d)���!�> �g�+����L�v��tC��^�P�SY����Z��/*~f�]���R��Rv�L�~��?��bL��C>�7C#���tDy*[5UԔߋC�D��"�������M�Qa��e*�n\l���O�b�����\Ԫ��A�3���&	t�=F�DlU�
�`N��u���x���Rc9��vV�x���Mg'9>
�:����醺�k��n͕�w�2�����I�9>�j��5WZez�<��9����5���Ə��rμ��|u�L�zn�����?���Z�3[��H+���G��p0�.A>��ޘ�N�K+�>�����RWc!�'�A���79���q��oπ
��
��V��t�܇��L$���8����������\�]�1� �����g�A�4�����*����-�Rj�M6=c�r[���K�՝#[Ң�ʔ�W���u�_�>�4`{z~�悿��F��V�K�P����P��!�7؎�����l�[�$�Bxݣ�{��B�p��7�̽�S6A<Q��Ψ
,ۍ9���0>�L�R/�F��L��B��D�f�Ӭ�������nQg�W
��?G 5g�������je�����8��X\�4!�^�(�y!ޓC�(�z�Nlnl��!�7w7U.X����n2�)�T_�v�GϮ'JlDŶ��7y�/8<�'�(,|����uM���������5�ʌ���V򯿓m� �ޝ�U��[DP��5F�Y�E1�P(��'�?��F��;79���@��{�Q!���6��],��Ӈ�����s�����N+�'��d8��������B�T�����X]�6~������=��܍G���&����F8�;U�8Tl}�B���w-? ��t�����D-|�znY�����P��݉���M�v� m �܇tG�67�r��:�e��s���p��an�O�x�M��Wi]y��'2��ck�"�o���Hr��d�zOc��a��ז�f/യ��񵟉��/7X�.#v��xh��1��7|9[:GA3�H���/���|g�&�6�'���"5�d�O�;����y�d��:Q!��[y�ԑ�B�3�ZL���Kz�N��PXB�2�*ܓ�����Y�:4��].�֋�i�Q���v�ǧBO|2�)�)�Jp��~=�fy�Fm�: k�eHAs>���g����sJ�Z\/4���"}V���0ร6 |�#���ob��������IJ�"d5g����P!e9���<�G���٩4�͋-|W:�s+�;W�A�~��X)��p���|��^��pd���	)�" ���$�6i����a!�`������ךﻓK:Y=_��S�K�I�R�s-��^*�~�]4).�+| ��ԞՔm{J!jA�H���x	��6Y$.)aS�{j�ei$��	L��؈�ߺIY��2N�~�,��b,��{��A�z&�yї;Q`��F�ZQ���#T![�>ҕ@��z{�u�9S;MJk9z�����sn��m��vӡ��0��ۈ���PztcS��E�'���}[K
�D,e%�QXvZ�]�-��|�Uȅ5a%i7@���(�w��U��ؙ�@
��r��g�x-rvu�����Z*z�Y��_BC(��2�c�r>���@��+�z� ����@+�ھ�m�������1�;6��q]a��*X��?l}B�/k�ک�dr�T�"�@�S���V���iY�	sŚS�&�r�龒 �@@��C��#�k�G���H(X��,#��9�2��U�Κ�\�0�u�I0 -�bᨐT�Q��&v�,���w]@�1��	-=�G�	�s����P(�)fZ���	_�3�i"7͹��q�B�`k9��77]�e��[Fv��k*��Fr��'L�W�8c˥Ro��!��x��:�E��M������.l�h�BMŝ��hm=�Vנwð�Y�ї��!�6P6
�*�n)t��4GJ�"�lTA[�;���`��S��P��w���gb�F�c;=����y�s�w��a���;�rh�ħ�0[�S�����r��[��v����i��Y}���`��T������c��;Z�	J�P��e��!ܓ�-�~��'�9�K�S���3��9$����"�2H�V���(  �Y�lo�{P`�F���N�Y�>5�4�J���˗ܪ�.���+��i͚�n���W��O�ܡ�D��v
m�
�v����]����-\�Pb��0�K��|àx����9�&KJ���s�Z)T蟵���}b��L��m�4���9��/Ts�G��/R9�t�����qS�5���b�*��Z�B�����Q�/6�t,=�F��l�t�8BO��vAL/���J&�u�
}�a��T���{/�7�.�2ƥF�7o�\���aB�&�Ц�M�\u���,A�'q�2�����񌳏7ʮXN�ƌԼ֢��:���42BP!u)��}��E�.3�]ڷ-;m�Q�A�E�OY)�F/l��6�:�9��x���5��|�}zX�95n�Zv�Dt�_4���W��M?(���%�!�_Ce3B���8,����yn���9��<�k�ʛ���-Yi�����ù�n��M�q�l+�����)�Bϒ}��=g�F��FZ�[���U����>x�d�Q�Ӑ��c�oK|ߠt0ɽ��	%�ێ
p�����!;�e�21��@���������%[�^u0��u0�**mA�,�12��G�/�a�bFw�eG�V� l60~^Z3Fh���D��o�����7����5��=}���?�q���v�ʂ2�%Z�[��O5��}�dX����n��t�VZ������gk�Z��+�a&�5wl�����v#Mz�kI�zZ�m2�;�$U�Y,������nbvp���!Ő\)��j����5�������'	��b'�4���>����r��G'В��^���$����g� ���^�:�P��;g3��gqج��>NM��d.���ou`�E[��>�E�<�	�X�tg���_<gpO�j��W��a����
�����\�ݗ��_1-�]�O�D����E��HS�#����� �''���vT!j:�N!j6*�q��9�Q)ߏq��yI��W��פ�Js���[h��$KE����s[� ����^�a��,1~��)�3'R��u�F�R����y�Y�~��lCK0���D��$���A�&'�pę?�e{�Ɏ��)	��V'�D1�,S�b�:z��
J�\�M ��HT�>0���*���9;�{�B��pnE�Υ�"U��t��H�wi�G:�ځ�D�w���WY�� :\�S޴O�GL�̤,׊�1Y�?�,
O�����{��3c�����rb][/�a�#���~��'r~Hh��v��Dx�k����l�)[���m�����K6�pf曔������eR��&Ⱦ��J2��V�p�ۭ�T��=ғ�9J�h�'5��<�e�X�K���	����D����y?�O����XcL�'�z2�[�һ�n����T�8N���D��4�c�qɪy_LU� �r����B�g�I��Y$3}�f��]S;��߁�a�
𚢾��r�,/>��T�����b���{pXs�d��/�2x"ҏ���Y�a�~1���ڔ�v®%�Z���X�T���LB�	"�	��C��tٔ3i"v���cQ�3Yq%RuB:�1T㦉���WT'StN�����4G@tq���ɍ�;;gi��`�󬥯�aI�xl���%��5a\>�=�p~s��1�ۚ�r�-���@��P��0O��lT�<�p
!9��)Sh�#�����M���%e�L��g��A�b�)B���JMs#�ۭ2T��;���r�O�rL˼��,G��J - ���ؙ�Ȁ�����)�K�JyC���F��eaѨ\��a�T��#��c����kI���i�Y����U�js��y��|*�JM&��w����s���v�$��3
 ���Pp�K�o��� ���!R�� ��<#���<x8���E���3l�몯@zT;�a���t�D'`��鸲�B��	M^�obYE''��Uz����#�|n9�d7�0*�{:�VH��qr1��r�WB���3��?\��@�>�^�A>?�p�����E��un�k��K/,	�o���6d��=��Kw��P�ⵏ!E>����Gj���
�P��tG���QU}砝��z!�W�q��a���g����w���ϙ�{��a�E�"3�\� -�d�s[�෩���6�(�x3O5�>��L���L�Yȹ�T 7l�{�����%��[�L�ƷֈXG� ���t��<��Q;����^U]��K��i%�-ƛ��DV�|��p� o4rmJo��������a���^M��Ќ�n�O�VS�����e�:0�ع��v �-O/���T�_ߊ�Mn��f�̴OZ��!U �Z`|lQط5�H��	Ӡ~W���J�����x�U�w"��!�Ͽ��ĭS��n��?z�R��"���y;�@J=�޲D�u��Q<���
e��D�a|	Ŷ?G:--=��Dq81N����[����WW���s%�w���ȝ�����S��5=n��Xh)����9wC���ՏD%*NT��ܖ�@�[$#��ij��f��5Z���x���R����ܠB'�Ms3�D<s{t������B��n��*	d����Ѣ~�;=�\#���8�N0�Tj�:��#ⓘ(�6Β��Y�fb�}(l[ܐ|��a
�a�L�W@2�'j<Q��0"l��{8�W�/��*�����PǷ7��螝,p��%D>��A���A��xrR�m.��GJ&�J�+ű�.E7vE}�یIw�s��~�npY��Ta��9~�� @��
N�5@�M�7Z�(�����!��k��Й����4�7.���N4Hk=�[
�C��
�A��{?������LL49��a[��H�쏅2=�_�A$�E2�Xw적�%�zZ��m���Z�JA����5ƛ�(WtE.&��	]��&��#-C�:w�یN�� z���q��.2	i5�g��Y �w��ՠ�� mE�a!b�?�����$����qrS�O\�س]�+/�,P��u@G�S+H���6�������p� ��rj�ߗ^'"��-y�rG�'���_A�$�.M�g�����3��-8�#�q�X3������Zذ��Ca��V��d\��F� ԣ��˙˭���|}}�v���Z���O��E x��o$���2�Pj��GȵAŲuR�7��k��gi�)��o��]�|nȾJ:��AN��&���}���~�t�>#wD�"�����F �Qvn�g�Ui�����
�^|m�J�V��E��L%���B��X ��M���x �E�E����|�O����n����P�.��f�4%sc�S�ߧ��⛥%�m�����4{v�c�:�UXcC�/I�av�pz!�w�A�։�+}���E�� �cB�rs���<���.��U���4(�c��l�,0E�i�\�#q�W���	���ۂի�r���pI���d<�p�@0r/�8LǪ�-��]�ȭq�5�B�C�x�aPb^Bݗ5Ǉ�>�

^nH.�މ�M�2�cB���8]� ���&?81�It�Y������}�6-�?#��ds��
ޔsp�{$�3'�?�(��,�H� o�� �h�S���O�ғr���)
�C���4I�JL�=H��9�v�cz_g�xR�q��� S�ָ����"(�g|�{�QJ��z�D���=�?�d�I����I�WU�� ����D���k̈́S�j��qy�<�(��.��t*p�V\�`��b�4ȷ���L�$E^vA5̨n.V1�a�%��n����IMk��khJ��v���uT&̒kK�l�K,��FO�C���D�	3�%@l#��m�[r�_�Zع-��^䁦�<�T�?�424��80>̶�s�0�����2rԧ�=zg*?�s�n���g����9�����?.�]�ouVc4ٛz�5৞{R;��WK�7���3���)	�M�1�[K�U�e�(/�%��������@�&�֋mzd��R��F�KN��-"m�Z:/��c��5Dm8�I�$�._3Z�h1�La^���T/�=��7�Ą!GK�#䛈e8�����}R������+pw3
�m5�x��ك�nˈ�	`�����佂�r��?�x�R��5!{�B��{	�PS�����+�����$o�ٌ`C��O���A�yX�9J��Uy�mR87>F�FoG��f%1oC�7a�ٶV�Q$�t �G�!�"��k��+ͅ�K�X�1����j���˺f�0�3g�
�2M�@[��o��w�3,l���E�^�{wz��X��m�'�l������:9�Ds��b_�?�RcY���o�Jx���6`ު�|���V�I��R`��6��@.��= �˻b�g3���@��<��%f�����1!��\���/�r~X��	I�&�� f�TCou`L�im�]I7/K%�rྒྷX�-��4�%��U�yY��0���F���]jEc�c��E���y�����d�w@9�i̚�t	t�a!
�B��޶�e�Yf�co�5�@V@[i{�����Xဝ��	��*��E'a�>�څ}PRa�6-�K����}ig6A[���V�ۑ=�nL2�+���q��,����N]M�&W��+-��ŽLn��8��9F������{
���P�{Mc����w���6 NK?�FNU�IQ�k�1�fR���/��^ ��|����xj���̖L�/*��행�So��n����h�zy�O���/+.�)��ٚ�I�� v$�ٰ��[ ��� ��4:F�^�u 6����r_,lQ:hb���¤�n���y���p�������k�`�MM�H�=�&yM7��4��ph���1�@�ʴ$	�~?�تf.>݆^�G��	��$���E�m�8�qd��TbVRt(X�������}p��7N&q��W����"!��cw cL�G)��u���'t8,��h4��k�z�Ds@x1�,�ͅ9�o�Ȅ��|��Ą��PgY�<Q��@�����_vI}�[�ul�S�������`����䂪�?�Je@O��'�-ǆ��i|쿯2�"�{\�|�P�z=���� �pSC�C��L�m���:�g�cJ��NF�p�� �3��_�T�Z(�y��!�i�=�;lD���󏆕	�W�ɹ���Ea��4����]��Xe�p�(���_�J -�%2�;qf��G�ڥ\��W"�tgs�ܞ�����.��έ��O�{g����v[��4�����]4q:exQ�ᝍ�F�o(+~a�ͮ�wCo�u��;�s��lly���nk�d?�H�*���K��������u֠�E�U�w���^�=���ȧQ'5�lL�c�~9qk�x$@l�ठaF�@���o`o�x6��u,�@��+��D�Z�	)H	pD8��(oܜG�y�ޓ�!uɪolҽb�3f̩����D"�d;ߞM0�y��t �������fޔ�_�*z n�[o��N2Y�IN�8�F���̘�P�6�����k ��f-�eX�y;!/�n��_�yO�(r�i����BԔm��F��z������ R��d��mE$l]���/;
0��H�g��JR̒���	c|���#��v���6�d��q�^B!7�R���`(�F�Р�{�l���)�<*P��v�UA����[�/���,��s�H��xw핀����d������5�(��~�dC��e7~���;9��[�@�Sy�l��^򒹏M�0�}p��Y��:YJ|�n��-_p���B�gc�:L� -�³����_��o1ZP��	D�4��٠��!�Ǖp}Ju�lYrX{)4�qg��b]�
T������J��G܋��^�5*�<���Er+n�NZ7=UP��ρ��mׇ҄��X#���-Y��i�.<�V��	�� ��!D*� i}k�>BJ��d��:%�*�R�o�H�ί�����`��쯫U%rh�����-��[��F}���Ǽ�Z#a1�9��p4���Й��3�R~������ ��Ľ�W��6�֐[� �[u��Ug�J�1��;�	�E��٤(�"0`)���]yx�?�����La����?#&W��dFG��fҞ\�O��2�b�\�֪���϶"y�ԖRZO����_x]D��!�8��n/'�e����*4)O�Z��?���) I��:��}�Y��'p�|d=�P��Y��uCe(�RQ��n��'��wX��$�N
 6����
m���L��q]�v7iHN����-� ���_�ٱ@�%��F陊�>h{�:��(�Q9����w}u��_���/M�݆���}��@]t*r��� ��Q+��'���7�Y_�oҀ��)
&��t3��Ta����B�0^˿��%\[Q���4�3�i����g���F������i�Nl�U�D[����5ǍK"���n��^���z��H.l�	:���ۢ��p?��^,�)�׭��Qn�H���}.�[y8� ��]�0�ۯ�m"Aly�X�b����;%~�.���S�b���|m�!_����꺳�\�Ԣ9�s3�A�F�]�̜�T	��@�)D2��5H��$�Ս��׮�t��my��ڛ�jhp��o�a�8>m%���׋��yYg�d����F��[x7��t��Z_�l,�9"�D��	RS��]��8���Uٸ�K�l�k���]$�_�Ś�Ӵv�������cX z����q��i}W�b`Oh�tɤ^@���ݬR�-�+6�L`Xt�A��JV�F���Dz?�.�|�|0�:>ˊLV����8���O��h�+EM�r\9�DH�7��Υ~z�ߪ��	n�*�!����`���`�,�P��p�
�\v�j�m;�n�h�,<�~$�r�l���D��:�j��d�v�U�\��.��0IL�ԿL2X(�6c;�⼍��}�^5��5y�	�ڔP��(z��ڡ�۷"�QC�x2PP�"6S� �2��#Ea�пL� �VA�c��`�:�X�H�1*��Q��#���¿vR̒+�)���R�ާ�&�*Z�/It?5��ʤ���G�
$��j/����-y}v����D��7�Ϲ�����v]���	Hȩ!9���^g݋��"P�4B?s���-���W�=P�iN�-s4��?o�q��{���7G<Q(#������}nL+��� �{�\o�>`ٮ���j
���u���1���%�{�8�ՏIHT�3��Ɂ/c��>�>�OWg\��(�)����Ɲ��Fy-��s�����ɴ�y�Sq�e0�ҝgʑE������N���b��4�z+0��}��.��w������5�v	[A�oN�k��F����d�Ԁ8D8��Hl���Ml�g� 1/�l�Ņy���ه��ʚ�z��sK�W;'T��MxH#[�qb���q-���Wn�~�7�>�p�9��w�)��q�,����e�"�p*a��{���@0�P��-�ܯ���&�2�5�E���lU�B|�袓�8��al���G��hR�T&k
��
Sl�{��������� ��@��1O0�����p�K�ˑ6����뒲�56p,$���:� ��NySȗ�s,�04�kIl��#X��%nJ]��k�����m��ww����Yh�+�-�w)g;[��|EpRN 90��Xdئ�#��r!i�.N�Uy���tY?9->J�y�~���-[�,�u�VmZ&|�W��T��]͕Flw��,%��V%8{��$TrC&��U?^'Tʋ�Ǡ��ݱI���s�A��-f}j��(-B�6�,���.��Mߐ�x�?��X��1�H�<bv�)����R	]��B4�*��z']&����v�V��u�iqEq!Ŗ�:g�q���"�c|�ǿ��)����ほ��;�� <���e���=0�#�-����!53�a"", F=B�5��"_3��� ��`.k�<�ca_�:;*i�6Ź��>��x٫'�2`����-�U��W���_�1:-��kB���zp�� �d�ԙ�K��3]��O��%n��TYף_>"G����$�_GU�L�zt��rPhK�-�s��[����8�q�3��R-n�o��r���_�w$W�ã+���:�s���|���f�3~��o�O���<z�'��?�X�XH2��(����/nwG�2.����yԴ��Z�В�/��:N�����)�)hEQJ���&��B����=�f8{bg76�-(��{�K�d��|~X�+����!�S]�2Q�C|�"��!o�..1��9G�ցkp�����<����!'��_^Ṅݛ��x�������#�bL��8$e��k���nA��Wc���!Ƶ����2�lk��$��H �۫,ʼ�������������a�)��K0�������C���z-�0�vG�r�]�������OeQ=���b�|�TX�-ViE��50�����E.���D�z.(w 7� {�Q�˳�&z�D��V�Bھ�No)!������ ;��2����'�Q�-��7�+	EA�>)~�.N��A��i�%���`z�����{�*"O���f`/�Ȱ��#"�w�
ݐ6􋷬�@�n�b�M$>��p�
�x�+J�(����8�=Y��'3�����B+j/�T�:��F���l�o�ka1]�]s��h5�C5_I]| '�Үo�I]g�nSjZ/�����vx��_��	i5Nz���W9�@~�9�g�!I�c�N��ff6L���/��͍d�&�m!NI��x�A�H/��kU�� ��9Ӑ���%��<�ju��������6���:������A��E#���d��!�͸�X�s��ZӁw���wd9�{/O�ķ6���_��G��HZy�+W��<z��ڱ,�h�0�8Ƕ ̇N�T��N'��e{xE�j`��9x�i�8��[��$k��Q*J�EÀ븋�`�5���\HO��͙9���̔�}u��i���4��U.�_*g���ˆ[&�󚓭\Lk;]���g���qIIRL("��S�9�O��Dq�{�����pz&d�-!���쎆=��>�(�R�_�mu���O������>K�XL!�^��A���R�9#���B6�������:����)²���������.�lA��cYL�;QlB��E�����*T�A��	��L0Zȵx{��(�~j �0�<-kϕ��|P�-%�B��,�J�y �s�s�{Qb���/1�7�>J\�I���B'CY�îi߆2�t�Ұ����st��KBl����zg{'`X�>T%��,G�B������-����̭}F�O�a�M<����V�Ʒ�8�f�Abk��eA��	'�-�H��+�9�����fZ(��~����Ql��m÷����i��Pҭ�m�T�S���]r��-Ϭp~srMC:���Ҳ(v{S
hU�I�~_�yH���ݸ�ׁ�kut�^�R���'Q�)��
�!m/y;�iakL�8fX}P��>��ઔ�?�mM�b�9M��ژ��z��{$�J/V6R���!��a�)(��>��hF��3M���@��Euד~R����A7Qm8�X���l�ο%e0�zsBL,A��K�eev�/k���V�`Ny���VI*͡}4�W�GVH5�O?g�&cTr��;�m7�M����3I���*��������=�3��Kۘ=�O_wnʕ��x넵9>�ʠ�5IV��lq�)Ow�`�4���<=)Ɏ-%ʔ��`�������(����	b��{	*������OC� A�O\�,a�=�9h�i��kM����_;.�fb�7Lf�+�S��p`�8��պ8�fo��~NC�3}�01'^i��[���o�gĥ�PE�ݨ9bq�mP|eU����������a�l>	k����3���}a i�r_��V�ͫ��'������@�ݍK꿊Ϻ^�2�ZUBE�T(�鱴d|���f�"כX�[����d�:�bA�J��B]�gH �W�PR�P{n�G�j���P�o���}�(;�S��ᩣ�:���D����f�����n>颋}�_6���O_��w�)��f��� #����~��,?�n�!,�l���m��d��iH �>4!��i)� (�x�Hf���n�x���ufm�4Q�P�ł����`����7Z�a<�֩���X����?�̆����@�g�T�%��uɀ=$�k���΅jR��s�G�_��"��ݜ:�5
XE7* oX�}a�񈑍��n8=�
>�a�a��;m��b/y���u��ak�*��6����r}֤�o�U��jTˌ2_o��� �+>�`��	�����E� ��K�OU��;��_W7YM�ajq+4�8��c>�ː��> �OǍ�n#���%�ߊV��	�)O7{���>���,g�௅��]g>���N�%�W�/%6����<��z��b,�Q�t׽� ,�n�F����N��?T��#)7��O�6�+�������I*�GH}�a\�FD�z���c�ta�X����5:k��<l�s4'�Ŵ��M!�i��#�l��sl�0/���L��������N��kV�1ܰ�ԝ���hA�+���'�lHo������K�b7W�D���@����;ONoQ��*jǔ��\��PAb���*S��1�g�	�:n{lV�C�:��+=OU�H��2c9 ��.�!2b�N�0!�3����(]�����ˡ$��!�6�v=��?;��rR�9�qD0�
�j�M��M2OAE�P�o�r�k�:%-v)=:}.�5��8�L��"���&J��r���T�ݏ\��9L!��+a�%�x��	��g@�|t8D!'n¯@�S����W��r�^N��Kt���Tiu��+D4�������H�$�P��w�g0XC�0�C���s_��sWD[8���ŝ�J<��v
5�5e�C��^�Hd��� *�S���5����q�Cl�~����F��d>�����-��5Q�=���
�`�}�Q�s��R��U�xD��)�=&�9������)��(�ߪ��p��r5��ӽǔ�8c�;�i��p?I�9&�[�"�A3a����N���+�z�~.w���O,���o����a��`ѝ�z�#�S����9y�B��FW��$l��g��LX͡v��C�7�ʹ��~
�',��`}���lZ$��w�B��v$��A�28��������!���m��vu��f�Y�~����0��b!�ƶ���u�tr�v� �h1KW�qh��O��Ť��C3,X&��_�le_S�u���Gq�|�_���Ws;HE21�px�T��<:dho�a�Ɖ�~��\�Q�Ma~���D��&�.��l�R����v�5��0Cr~�c�����j��ڒ�x!W�i�B��MFCv'o Y��b R_�d7�؎��]C��*:�x09ɭ�����9����'Q�WZ3����+�:U�89N��`P$*x��5'x�:6�B�W}�ְ�sڻ1��J��RP?�5s&.~45mY�M�y��o2=��{��s����a��3θd�z2(����z1ΥqHW���������4�V�м-)E��6���
 ��en��!��j��∉W�%�67����'�F�VL�rK@���5�xQ�Yi�:��f�F�=�^|C[Z(�<��;
2���CV�OpdRy/}0!��b� 3V�qe_��-Y����s�et���˚57e�d�.i�`�{���4xЄ�mw�j"�N�����^c�ȷ;��|]&?,�8s{���3�{\����^N�'$#�z��3ԒK������q���T��t�}N����W�9�v����|�&1E�1��5>i�Or�	�:�(�)�/���K�&������ �x�� 0p�u�f���zi�z��G�$���M�mIsFW|͠{>��nS��w%���5D�n�9n'����0��Xʆ�z�/�qP���Mh[��gJ��X~�h��q	�$�v�V`�и�d�:~�Ɗ����&�PREi4�C��*
D��������9q��,x��%��6@��B;�K	ϯ; 7M��{�H��/�v�K@���Zz�Bx���o�K"�sl)D./�<�ExE(�=��)�lPݧ��5�(�Fy��_�r��}�����,�%�<�TXÿ�-���.:.�~����>ñH>�hp@KH�M��2[5�6j&V��S����T�~�w�
 ~聏�B�<���T��*�#�F��4E[̅m�$�Z�s�/O�.� .�'9{#��k�QJ�����(��C�c�&g٪}�,]�ڴ����]Aj�B����d!2�kM�}4�ƽ¨M%�;�J ��uu������P��F���4�{�Y�;d1>qʚa�2y�'.g����!���T;� 9���Ѧ�o�jγnW*
A���" �|��D*�X�	/��h/��Q���J�٪W��0��~�
��up� ��)��h��IՍ�L�4��CS�C�+�t��e1}4�Q�A�����__�n�yepaIF��?�;�)�`���ٰ��s�-uV#yWO&ЭoVp�B��Z��C-�e&��$y�r�MH�����W�:aJٻ�#�(�ǰ��7P3Z�5nܩ���O�+L��B��G�f,�;e`�����7//	Ϻ�٤�O�S����L�\�L(�M�D��c|8�3W��e@T���~����X#���R�ۡ�.�)�2v*Na�bƠ�����~99��h��jX�0��n��
�Ld�r�Q���I�3T�[��4���Q���%mյ�ʩ�ͥ�*�Z�{XMWw[��f�~�|�.&�M�D"�2R[>��.ݲ���&E�4��.��ʘ�e#���{2���1��P�l�*��`����_ ���G�ƺ��l�/�pW���V�ȝA��ڌf�*ˊ]������ً��ٻz�>A?�F�	c���zp��:���xЏ�K�~D�I���g�-�i-�M7����7���&V�6���QW��:XL����������Rf�|.�#&����#� ��1w��o��$���$�£߅	��:��ڣ
�?�5м��`��*�hə�`���0���t5���0X�a������V�ͬ^���I'�K���VQ�$`������H�	?�����E����v��
�C�`Hm��r!�Y�Ao�{��H9X��5J��x��Ќv�$	��mM��#3kZ���"��r��	+�v_h�Ɨc�b�Ǽ�؜[��I83�CLD�����Sʄ��a�lU����i��e~]�(m��"Hʐ�f�9Ԭ���3đ��
�X�����b�/M<�6��6K� .����OK^�)cO�ʍBR��/GK�B��#����s�v�EK�X�pS���H�>u�p�_������w�_���o7�IS0�}����{���i۾΋���"���ٵ�~���1Cne��{�Mˢ��߬z`���H;���%Cm��{E5�F&T�h_B��V\T�ET�����[����Z3�Ӗ��+��@�>���p%y��j�����0��é2[��/0�v>>��yy?��#�\��� ?�m$�/"��/�ym2B͏i��ZT���
�(�����Z,�U�����x���eV��o�
c��[��rL�+�Fމ��V�`���~���V�=��8����^����$����gmSӗ"x�\VS��:a�-9(������U�6��	:-��r!�!�F̰�� �K(Q�u���؃� RXH���3�Hz2�截dH��R�u��<�Uj���1]�^n�0�*f���]������;f��2|����Ia������n�vH�v�Ni^H1��.GF�������dm���(�eu3=��y�w=�b��W��%~u`빋��;��&�UpI��6�M<tx�L���5���T��������o����X�a0 &u
p���B�{`�e��?�w�_��6ka@��H4�L���u�O��Bwh�g�k��9�h9�m_["���U��*��8��O��b���G ���e_�uS���(���s���aJF�5��!T�	Is?k��:M]Q�����D�a�F.d�e1+|@�K+�W�>)��Y�U�m(� ��x�'�PE[�'�e{���x���L*�`�D���B���AG���"�v+xr�7��Z�*5�9m��Z�m�H�;�=.e�k�ܸ�C��NlQ.7�(zX�觉��v=� �g���O�&�)�b�Oӵ��@�3��v���!\�)��	�}����q@C���zV� �Y]��`������=��1��H�-2m,1�hg�1&��&���2 =ѧA���Te��*���{Ⱥ��gq��Sc���_�-^��Wn�V݁R$s��rj�t���bGǂ��'�V�2u�a������+�D����\2�nk4�-�D�����t�R����e�Ĥ����'��b-�)z�y��۾��p'����ߩ�>�[@��[��,b��JA����v��ʽ���{|^�����Һ�%��JC�8��2���9��j��
��-�9���)�Y�p�i��h�P�G\�}�,�*���%��X^���/c�8
�7C�����=,tl*ނ ���o�I�4l '���=����ı�'�%��%�W���U@e���Փ�6�p�m��H
���'D�&0Lx	�P�/�M�O�@��J28<3vKy����SD^��w)����_#ź꒡6����c|e�^��7�6��uA�������t9\t�l�`���<�H<C{3����ܩ%M��s��� 9���!����x�(*x��8�J�-YEbiBvY�Y�Q6^1Gg���BG�`��=c�� �b�煩��Qڨ����з6P�i��@ 쟊�bmf�r^\��a=�Z@�~���;����F��K]���t?ǤJ�o`n_�S�����u�����E�N&���E~ΠVt$WcEZ�Qh�=X�B	�3jko}�i�;�K��H�����<�;ʦ����[��9G2�ǩAB|�Y���u2]�s�gLr֐�ύ��"�t�Ii�?TH8ج��˼�%�6bD��X+����z�u�h�m��{��@\����,=��L������ѡ[Გ����1}jז�s�l��<�xXG�p�DN����&�a��ޛ�6?N�s�.�Q��u��ڜD�6wpۍ�6|��w��[�=�T+����W���B�|%q��%˫qO���|��o�Q?�ke��af{��mQI�=�}�5����2�k1��@�.�6۪	��@v�֜Z(��4����Z/�A���!ޅ_��~��U�%4��z�C�Z@B������l��ö���I��p ����üf��)��
%�826�a� PJ{������NC�ছ���������؟Y�=:M�F��B����E~�=_N�Y�C���?hp|�����f���0}�iv��"��Ϝ�GK�Sy���Yk�N���PǺC(4����oA���; �_"���QZ6�D:l__�}lP�H�G�����G K�[����������)��G[D�3�>�������|��g���><���!)��y/�-�����;eO�����n�IA%65��^)a����O�m���,���T�+fU[�M��2�}=�R�y�4�AB���f��a�/Jjx�'gE�.�US��y����Ѷ.N�ܹJ���~���2�E9w�ӕRw~K*~<a�ǅ�5�y��6ۇ8�0zq���	Ln*�����#qC��*q�+��
��+3���H���������s��3D �!i1j#&Ј�0'��W�6�sw=�V�����5�i�:ֹIe����vb�,��S!Bb�α@�$<Z�ic��1�.=s� �Ȝ�V�N�6?z���_����� O�*2��{�*�92��o��r�������;��N�UUCo:Vh�e�������=�t��Se{zT��Q�md�[��mH~�p���"��g�/S�Uǻ�<���d����SS�
xKey�@�-x�����;W�_9��3�g26�tE�*�i���d������j�砌/S^�_� .��^�Ϧp�������l;)z��q�'�x���o�gJe��.%\�te&�C�]�łm�֙6�c+^��m ���D>�>��4��0n˚�d���Ca��t�������)��(Y��:��(������C�\±MB'H)�o� ]�u��~/R�Q4�zϠo�\�&<R��E��r&^�=ˣp�P_��T��	h�.ZEҜ6ഹ�|l���H>C/؃6�s���ˮ���b32��
7��#ͅ6�O���4��RY���D��i����*�����9
�̱���^zm ��X��oj7뻶V�p���"����3h8�����H���Z�y���������;M�O��O���RLұ0�[��_������� NW�g����Lg7�!�>�<#3[ɫ�,2]�|6f��t|�<eI��!:=�����f��Q��4׳a��zԽ����H�eSH��,S�g�����E#܆�g�,���VS5"�"|�z���O�	x�U�x��0z������N�.�	���}ϳ����>��� 	S�l!q�ѕj�2���q�y��u�Ll�0g�����{ݴ05�I��	8����[b<��%#�߆���6�O������l�K.8)���Jޏ)r��Ί�����`�u�!;뱎��yN��St��]+�t&���<��Z|��M�MM):!AV�1�5@��ԫ�Fz������֒K�A-,a�ˏ��I4n���
�D9oI���2ӻVfn\d�˹����DtpH5��'6Q�G���jsUt��TS�Z�oaFh���`��V�x�s�gF
WV+8�y(������GQ'��I�m����v��3�s����p!�	̗A�K5�nO#Đv+�0,��/(?���腨��"=�|�v�P`�L���p�}���:�'2ŀs:��pfo{��D& �zK�H/d�]���Z_��Y�+k�؊���$b[�v'x�<����f?3#���P �o
��.{�f9�!<J�=D/\K(�d섋���V�[�x��'+��=F���7�X1!7�sZ�E�ɟ�:�Sv�$�G���	)�xяs�[����==�5I�"�=o �0f^��Ӟ`6��k��z�۩�Hn��J�7	)�Zh��(��7R��ݙo��^Q�GU���-��H���#�O��wa`���5��I����2$M1:ï�f��t(�M@w��fV�B���|�+�1�E�*���H�H���
̷a��!�Pcm�O����IkP�FA�N���r�+����\HvĻ�h�w��sg�f]��� @�\8�N[�U�������&��q;E?L�4c*�p�l�jl��W��s�f-�*�j-����3ßN'��%���*�d�t%�C/�LOԘi���Suw�#/�*ۿ6�C�3�fS�"dQ7;��*�x" ����>���l��4􁓔c����pmLL@~���5I��S���)��ͦ�0���I�mo�zlq���&_=�0��b2jW���:������_�Ian��'�˽^��⿬�;n��.�����v��(B��D���ߑ���T�`*;"��=V���K��d�V��몦��."�/Vg8`�A����鬔�����";Z���~������V���dB(�UX�<4�uȾ�%��XH)n/�Q�?�����OV�=�ǅ� ��Ji��MO�A�D��6�ME��w��`^��FgO`'�߉}~��-V�fR�ŸA	�)T@��Hp��8a��O�eO2�����^XZ��&ܷ�+��a�g	���&`}��섋�Pfx"P���N�t��Ӯ���g|3Zat�#���?m��������4�-����~˟��l�(�T�����%�oZާ�|�O(\�ց�(\mM�"��wt���u5D���������U�r�4z6���{@��2�ᇮ~$�d�� ��
�9Z >�2�@�jP��?���&6��G����7��ʔ8h:��J���xf��>��s�x���H��^W�R�������i���������
^sa�$����0� �����5�������-c�-�q�-<�0�x ��	�
0����ģ[j��H"���1X_�Q��<�)�Y�RW�<)�>��&&��̇�CO(�zd�|sa����d��c̩��[�������_,��B�3)o�r�m�Q��J�����o�Ձ���D$}�^
�l��UR6D�}z~�r�$��U|�r�/lN!Q���*�ӕ�e{�a̴�FV���OV	/�Ǌ��+x߃	�ћ0�����"@�I�ڽ.��m��C�(�Cs���j? >���3�fe�K�s�P5Zn����A�&��o�s�����??&0&��Gԏs:�I�f���D���ī�.�Un�U�������w~��#���	� ����B��)��U�:u�_���e�]&h���.ÂJ���B���*���c/v��4<�T<�S ���W��
��W�z3(�Zl�
���rs.@ ����+�%��!q��A�չ��/��# `�R���+�L;N���C���7tK���e�BW!��X�����)��Z�@]�w۞cnã���u|��@y�2�L��h��Fv�71�F�y�E����{({�����������ގ�������f�7zSOZ�z$�N!��k;�M�P�Җu��Vj$��j���� QK�j;���
��{�؋�A��\@�Pw���o�ժE���W.��R�M+Y�J��{U)}}��kcMןPГ���s�0��%
��e�]�=5o����alX#+�UEe�`A����gB`�z�P�)H>[wG�]����y)Z�a�^TM���<�b�@�g`�̻�:��]�Z��|d;����p�¸��A���1�-��(L�gr�0�V�o��a�m�ۦ��i�G����K���E�9���w�T;o��w�˪T�>�^#�����)����C]��'��&B�K_��"5�<���f��3�{'\��#O'��e�����z��D�}幡d�	Ij�%%�z�K���{�ǹd�� �6Cљ��Cd���n��%#�9����Ѥި�R�Xbhu�5�h���%,rÅ���#� m�
^W����T��zS��F��|�9�և���#����m=�E(V�|��3`ZM���(t��$O�L ��NT��\�x�d���0��~LڃG�W	n(�8����yNk�g'��x�uP�P��	�U�[�b �R�|��h����~DU<#�B��I^�?������	�9����c�c�62Z1�b�+���lJn�/�M�����i�,���S�ﳰk��"���r�=�q�Њ������k	��]Ǝ��X�	���\������!�4���בtA�D�}�&�x�x����ج��Xj�Bɚ�Pz��G{�59�0�!�����E�˧{�_e�+��B���#g+%��j����ϞQf�9�#���{�+��$U%�'Ô���H̔�b��ݒ�h�!�]?~??�O
!0I��f�qIyp�x;�B�������O�t�$���;�E�*z+����(��%��D�n@���[NM����7�wP�ZO��9�6>KG]��΁I�
k�%�pHd��w�9�X|q��9���{K>�F0묒�ya�������M�o�!�H�,����]۰�>��Fl�#G�dF��� �ő�|�JҬ�/�����|\��&H鿛P~]�K+�4D��c���J%�.�pE�<N^������j����\٪ZcEQ;@d�Կ1--ɦ�zc`x�x�v�wb�_�Yз|B���t�6����/&��0D�P�a@�D��ٙ��^�X:YN"v�C��{0+���Nf@�?W[.#��4\q>B�K�~�𩡌�!����|������gi[@>� �|�P���c�ݵn�8�۸;n$[i&{,�m?~�N'x�)����	`f pf|�q�O�y�u�cz��9I��"N�b�&5�)����[�RO�f�v��
��t��R���eU܈���W�m-��r"K�꫹E���Q�bg{p��?_�)1�V���=RS�W�A�	4��X��&+�7��q��_�Τ�����g9=���x����<��9/�ѻC=��SN��Uk�o��j�����/Q��U���m��X� X^�+����s�ژe;�sV���2��FU���R�ȇu��1����Xa����Xy�\��Ɔ�Qy>�546 ��!n�����6�\�γ/�����ZS���duyE�y	�N�ќI�Zee6B�?Yc��6T$_�����c\��=�����Ϊ�[n� } �B��:�.m�:�N��{�{������L��>j�̆ڙ���)��H8��l`�6V�𺅽:��$",��_f$K��eLc��pcD�yh�W4�Ɍ�3��
��YNx̯��x�s����k���7�w�"=Mn�=�Ǔ��~r<7e�����4[��л�����}^�y%�R[����x'��#���Hlw}�a��+j�g����À��1w]���{��<�,f�je_���49���&V&�%������$����̵]�������� ��?�\�Pad��W�ly�a�h�	''B�R���� �B���I�^�2�)��K��ΙeBX��.�C�1�'��x{�"Y���Q�mӗ� <?�sU��o�Fa����n9��S�di�>QB�b��)�fE��y}��V�+��-6�x���S�Q��&C�T��:�6�����95 �����&C+�Y\Q�C�"��s£|��̖WC�<m�/�]E��1E9z9�v*]\��O���L�����9���Ք��J���,v�s�W�2x|Ps̰m���O*52����ZM���O;�&Z��\AF�ϻjt;D2�*�Tpd1o:eL7�Q�M��5~��`A�7�>_�S'׿�Eຖ6�;�����UD�M6�'���=Cl��;H�b_�����[�I�ү|sc�$�r�FG>!��mAP���i����� �ҹμ�]m�gcK]��w�ߞ��[���ѳ"'\%��u���}]��%���<�,N~,p��Z��dz��C�E+E��Ͷ�*��I|�
�md���\��]�Gl|�O�xf��}��X�� dW��fod�P�a\�v�D�h�^x���r��������i�R�m����`&�4���_Q�x�ȭ�Yj��Y�����LGu��Z��k�0ܲ}/{��(8�,p9�>�.��.�,�T���pb{u{�7fx���~��rLTؗM�	�g)a���J�����1p�� u��ǟ��5��
�m��Q,^%)�>�{����Ɋ=�<���G��4�����*daM�< X~����T�f5�y���HtUA���&��|P0[���{6~�T5�O�gx-��=9~�-��y8�2^� �뱭�o��2���|YT���6��B�������@�컰��x�?k\u��'<R���ڊ}^��)>�����;oZ��ļ�j#�xY�z�?΃�MNeGq�����W�
L�����k�_� �2s�
�X�'�k�ad덤l��k�v� ����<q��[:h7��FsM[G*þ4�Ψf��	�/N�e�z�*.�e+���%����٫	�΀Hi�>%���彊���luo��B��V�рU�Z�ټ�r�r�����PI���5U�]���������Ӂs!HN=O�?u���U��A=�!e/�Q��;��(Moj�� �$�zQ�RZ��G?��`����V�9moa 8�}ξ�a1���w� n�8v�'m���[�M��_�\�6rkYpěM��3���g�X���!���k� �)^����
��i���%zj'.���7���b��or��dU�FH/T?H���Ƿ��N�����u ��	���}Z��8�����s0�Pi��;z:.VR��>��$��,��p�ʂ�V��x�cL��P�=?�c����ϥe�3n�;òwEa/�#��&I�^�%Tp{:����?��m��w�;����A���7��u���O<���֭]�Oj(�n���e)��>qSr����(0�&MY0H��2\�o�2�h�C��~B�:p�ڵYe��.�L�'��Be��$�B�@���[�ޏ�l6W)M.��Ɯ��`�WB�X�Rl8�{�X��o���$��R(�x6?~��K�aNhq[����Y޶/�5�?'�P)��k���L��SDT���-�i˟��;��,��T�\����0��A�l�,��3���ho�5נH��r��b޿�P�(s!Z:u=�m��{8�غ�Ͻε�3{���RE��`n�k�ϛS��9�����o��.}62p�M�EE�Wr8��ĳFܙ*=x���t���ר��G�iL5��E�\�r�֝�(Sl1ޜWA�$��f��g��Z���Cb��Y�+?TN� ���+���mS�]
Y���Ķ�(��9'T�y0p���T�W�PG�����4xb?ƈ�����=v~!��1�"?/�&F�E3���̲I�&�0��\���n,��AB�a�9�33��8���g�ĳ`W.`��6�F���!ǆ���ƃ�)�忱G������P-OS�zN˘������W��-d�YN�W�#rB�Ȅv|��Ɗ�af7鐬�Irlo�1=1fA��#yG%H51o��V��(&+9#�؛p�)��*F��J��W�ƃ>�o�S��y�{������}2��I㿢v�����A�Z���|��@��u"��蕪h��%5�7네�� �j��d�>���Ǖ`,x;�ր��n��H�C`!��t[Ir����Ҟuы�|} ���cc��G��0�B��xO�&�	+O{��wZ�Ǭ!�Hɟ^_U�r�[���������T��\Nֆ�XL�B�rR�u��}�&��Kx�ՠ��J4"��>��R����4�O������%�s~�0��[�P?mbz!����vT�hfvp݌�V��oF0��E�fЩDk`P�wr��B+�=��*��}y��Æ�鳱�ۀ7�zɎ:�0<~�s_�ݏ�/:,�k�c�
�����S;�6'qgz�0`Wڲ�� �e~�OPN*Y_(�}OnQz�|�0�"�4Ā��Ȇ��N4�Y���b:�N�X��ei�����(H��<���D�R��r	��c�[�em��Oz�*4��I�!��z���jUHV��CǷ�&�.�%��m�r�o�[ҐB>�d�|�aȪSdӉ������a��w�u�%Ͼ��C�(0A5Vh�@�j�V�[�A+��HY��b�AF�8��v���R��kjbV��V��n˟V�,�{2[�~�m'+�쩺�GM�N�p�<���A���,f�"I�-��~��=�L������B�S� yIʤi[T�	E���lX&��: ��k�OG� �����b��n��q.C�r>�䥇8Ǔ�iT�\�`,P#�S���n�1�e"H6��v<�sU��8q�~Dn{v7PJ%` <�ι�ȒDğ2*�w��et攙<�0)��<1��p�l}2@�ռ�P�f�H48*��wyi�F�P�Wn (Y��V%2E{r�0��n+/����3�<�i�8'lPD珁�8��~tA�>U���%+fŃe�Y`�=��¼M�Z ��O� W{����X�
�fSg�~6�O�*�͓U��wl&�R�pW�~�>�D�S��4��h�c=����������%����(V�YDL�]6mpc�`(�8�v���?y�#F��l��� ��8�6%�b��-�]H��q����a�ʞ�OU-�0�K��K��f���Z(�3��&)��{Q�jW��mީx�c23Y� ��L�k.%S��͋���|�I���~2�X�
��������T����7�?m]�l�nO��x�+�� ����h���
M���.������N���!�sS��;c�z%�|�u�>t"���a�PRﰸ�c�#n�)�W��[x�p ��W��d|�
�:*�jL8�[�3&�o�C������H�3/)>��#�D�wFF�����0_L��>8[Z�|���ZD�ё�$�k�HaL�sT1�X�l&��
K&(���z������:õM%�!�����򗰭�j�d`�x�0���[T�7�LE�^Ϙ�CC����:]�-�[�O�^A%ѻ�zkݳ�-̇f@WƟ�p�H�FO�#r��Zd����
�V�MX�ӈ0�8������c�����V7��X�)Nv�/�
�4f��f*u>@�v�`�����]�g0��)��0?������x��%@;U�	Α�cv;�.HY�:e�ΰi�<�
�lȦ���'�*���J�����
;}S�mf$�/�4Ě	�7)��r�U~�Dɻ]��XV����WbU/��M�R@�%yDb�w9My���r��ɼ�{������_�JD���W8?���"�/e�޼��j,�&����21��G��y�~��B���4iL�H�jgo G��]�����d�ɧjY��[$��b߃��_�,=�;W���.�;~��Iqr�`��}�jɸPOGW���w��Ngk���¤�[��2��'��s����p��-���^?x�s�5�, ��� �C�OS����&�����Y��i�"P@a`ST�JbH�?�ٲ~�O�����F���� M>��Ey��C�뫍;��X$�r���o(,��>����|�8�X�j���G�c4๔� \?�P-@P�2T��{��r����j��7��H[�'1.KJg�b�J킹N^��	��h��>��S��+���]r^�h�Ph2=���B ��~�iB���3�B��nY((U-�|�U�.��9u��
0^`y~ZY��L�%}m2C�{�e�f�>^��Rtb�I�#�����.wbe�Ǒ�{�-���2�O�[��'�rEY��5��`Y�r-K��\��� ,]#��]ἆH�#����E }XZ-���xθ���nh1���Y���l���'���se���ZE�B[�析�$eu������q�B'�K�@��A�ǌ��e��p���V͍<�>
A���D�:O��R��ÅV@ο�3�y'6��B�\�"�x��Iw��xVf��e�L�γw�Q��Y��`a�z���7�S�f��`e{)t��9Rhr�[����x�96E�ˡ�3�äl
l'��!��4� �W�u�\+w�\��4]���I-e��>V�6
�r܏A4RY�����d��/,�-5�	���k;#�	�3�'�;`�)m�;ѫT$���=�.*��h�쪘�1=��D������&������w���3�P^*1q< �:>vJ-Ɲ���;	f��9K��شz.�ڕ��6�E�\(�^ύP_4�$��y@t��S/?�x�t�����;V��pU�$�I^͕ˉ`�e&�)Z#;y�<~c_Δ�t/yt��ڞW�N�"�B�H1��TD.�_6�5�W����h�Q�����8�c��k$H�w^���U�?/Κ�r�ћP��غ��-�3�{/6�53��n@�	D���''��<��lRb5#=��K01.O(�BS@����@y�L=>LCü�yo����E�׫��lLp�5j$����k�<5H���xM�z�]������&5��6�����{*�B�v�4Eτ)�1t�4�4i�k�ǁ���?�Ҝ���Kɯ���oe&G5gɑ����{��M��,�w�mk��i�����R�k��lED7�ñ�3�_���{����D-o��t�s��Zk�R�����2bs4��X��
��ӯ���Z=:�'!��w̞�U�jN�u�]!r��!�+�~��J㒁�3F#�T�r
i��:�6Go�nWt�%�X�3w/<�%�az��w�+�����w����A���t�����T5�;(�{ޟ��Z���R�YN%Y�HB���;��h{���[H���K����}��^yԱN;~���I�g�U��胧�3G�CΡ��e��JP �D��n���_N#�ͥ����Z�O�2�{\n���&+{c�U6Z��ߨ^͏��ڌ����C��x�O-'���ŜK�ek}Q����_tr���{��͖�B͑�Yr��Gi��5*$f�$ڗ�{R�q-��KꪤW�s�z��Ts�dC��n�+c�Y�%��d��ĩ^�(crP�����pؗ'Q�C3�5gY��F7>���'�$
����ҩf��r^��W�iș���<�o� �U�1��f����J�bcC�Ak7}ڌQ��ti5N41L�N(5�ǃ�ί��kU|��W}/���KlqH9�#҃e�N9{i�����3}����$�	?�+��פ����=&�H����f����h���a�j����1) 0IG�،��X���O���DT���H:�%/D�Щ�̇
/��N��]���KD����ftk�����1��}�V�)<�n*�ʛb#���OU���)8�<�r��}U��ПÏP��!D���K���圱9�?ǵ-��;�.ۑJ�Y)���Wf����bcx|�@���|�Qw(�z�o����34N�#��97�u@�C�d'�4�
�,A����o��_�`�SI��4k���Ht��}^Rjx�N�/�*𡖕O�S?B�
�\r;����S���Q��H�e�jD
��+��t��"���o�F���ƀ
�ߦ�.�oaSŗ&}˞�)����Nݨ��������S���?�W��ƝH��d	�Q�&`�(1�;�W ��ɓ����Q�b��V_�Sh���H'X��6E	4��J�$}�x.`2�M H�=����U1�.NЗ�[,E����cq�a�P�њ2��'~d5��Q�y!�/�se�J��1&�هz>�`�8�釠>l�r{�� ��B�����Br�x���4�s@	է$���\	L�U$j=H�(@6>�b��� �^+�@ÈG���9͌r�\r�y@��
�9E�$�څz�+j�4�%aݑki@�妌OpjNn�����/�>{���sjЬ=v�:�'i*�� ����T�G���Q�qB�Z�=Z����������n�xLѦ��wG�� ��?���{��{aS[`{��3v�G��g�7{c$�!�h:-���W��z;��m���  �_	��};��yԠ%�)l�^0x��ݖ�X�~,�k�b�G��I�>�E��0����R�{�w�#
�Z���$��2qWc_��ޏ��k�
�̎�V`�H��������������$��f3l��u{��'m	@v����q�c(�m����E훃�~�.��*X�	���,�&�zpң���W�m��Z�'Z�r~SDz��.���uuR��I��$�4.�r��;����4�.ѣ��t�.TF�g��3+�q�y<w*�-�V�)T*!:��`n����X� �h�� ݣ����
_��xޚ�{R���ni=ͼ�s� �ѻD�ΕM.$�R�l����7��D��~��E���H�>��Y������)��[ĺ곃��,*�t����&M���!D�ž�eeG�r{�;������g~����nq,�}Ԗ�#O�j���/NQ`sO�e����P��)2�>�K�E���0![����ؙh?S�&����߮��B��Fl�.Su`�?b�^TZ]����M�)����H.�Y�Y����oЕ�.k{)/˄�Պ��I)�����R�~�!0���bWK}�04��מ`�J���D(54�-=��yO��q#�'��[��
i��y.��1�������[�$Q�g 򅁸��:}U6�:կ	Gs�������ֵ}I̑K|?�]*B�`�l�fO�ZoI�z�R�Ul�y#��1"]j|A��ͦ-&��{��5�}�R;�)v�,��:��}��J(�u��d>oⰞQ���<N猝`���KM�q�:������wŸ�cO��'�ؼ#ų]�;�k��7u�R<����w����x�Ϝb���zg=#�zJ�#�"�/���s��l��<F`b�Ov��o���2�+��1%3kz9s�
�PFvu{�H�ӳ[�ّ(��� #\|�*w��(�5�����
��
vL��vI♽e����p�U����nP��yod�|J��	p7���c�Z��"�p38������:�ԅi0lT�^5� �`�%�����l��\�W�E��8� �&��P�u^���Ҡg���Sk�"�H�ת&�LF�Ϛ����%��i����"-B���A�e�7NK��t?���x�<��nD�ķ̃�T������M2|�k�P��~��1��#v~n��\�B�%�g��qP�$b�[s2�=?����CA>*���,���d����$m[ͅ�����ZP`�5��v��*�l�p��f��v��"�lk�ž��l(
�[��~Z����J�?{�����W���dk��������t����|U+�J
������U��XMX�W(nh*�p���d���N �p�N���~g���4�$�m�a�2Ȭ�������R��j"�z��#���}wI��g��?��Θ-i���9���Xߡ���]wz/����C3�衢$�>����L�|ʦ¿�(Y�o![bQ��
 �F��ZFI���N�$GN�*6QJN`��d0���m����{}Kt�3����j�*�x1]�h_�L���`���N�@z�]��"�x�I�BE57&���i���J��eZ�c栀���4K��x��/��r� xg�es�f^�C�y�����#̺�~B���-6���y��?} V��+��Yս�M�o��uQ������v�mn�L���p�ʷ�x��e ��N����.U�C���k�JP��.�ˮq�����՘���$����-�rR����"���`);o��N�!d0�XV+��-���xg�B�� k�1��z���T�]��h�sZ �#_0�	��I~��,pkPe `��kœ��IͰ��RVA����-Z�Y;b������*1ͳh��:m0�O���v�	K�?��3������ ޹Jj��y�=�1_4�GJ���c��.��3�-�ji#Շƒ��`JpK���~h�coe�M0����J��������x_��~�!�ok�	&O.��m�{\�YQE�2;7�d����go��i�&�b�Of6�U�肽��et��*7��7^E�	"�F|��@<��[ҁɦ��E��C��R�S|՝�t�,~�wȕ3V��=_:�׸*rZ�Q�h���ٟ'��G�5�N���|%7=��1���F�a���8�?q#�&sF��y7�ͽs��D?^�QTK��N-|����,c{\yY�f%!���0����Y�� !��+؃3��ڙ�y=u�rn��Io��e\O���eB)���>z�'�S����vu��:��ʄ����0���G��F�`�����w���H�`��?<[���Ovo.;���-�qe<�-51S+�}#��pQ��֎�ɔ�ܞ��5��q�U�א�t�����\�#��`>9���v�b`�t��I>�OFfV����~�;�z�He<3�^_j�%͇�QA�yڛD�j頃��s?��GU��T����67� �����U~�aɓ��D?X��T9�PkHL�L��UBƧL瑂����<��S�G�����78��x������x��)��I�(��پ���̆�˜��R�9��U:�Z��,�`yR]!�y��� �e�g�
����հF;�|�*�Y�\g���Yy��췾�'#�G��|
!L����Xz�}t�<��AĂ����OG}ի��r���N��$�f��"w����}���9d�7]+����� �����mr˟���c�� �e����Wc��}'|s�#9`	2�� �$�ԃI��Pϊ	X�W~솮���G��W�i���i�n'g��G	,��g�UK�6����x\�s��a<r�����nhxT������~5�H*E���0TZcڱ��ru)�)������`8�=ߤk�	���U�ՠ�,>Du|�E� L��lķ����j;�����ub�Z�.�d�îK%����;4��=�X=?�9m����{�lG��ne�>fc��Wi�
1~k"ǡ^�n�o�v�d��i���Jac�Ugh�F��՞5�saf�l�K�����XvJ�����P�'��|R�LGǆ|�-S���a-M|;α5���V?�t�	7�C�ҴǷD:��-�|\;�C���������-�x%�u�UU��)ZK��_��b���HM��:)��e�u��].8��N�������D����b�
�p��xbl5�=	u�� �s��k="4��ƞ��󐾑Le>~^~>��;�g$U���߫�Vn.��x�k�)�րq܉{�Iz(/��9�Ɩ������2�N��C��1~&�Sd�����f��mj��p}���f�������.ԕ��F����8�Ə�r�,�-t %�I�ޏY�^���٢^������֢�\�My�D1�|�@d��(�n����Hk<��l']��`W��/�a�sJ>���o+h"��C}�M�M����a����xu��y��$ ���S��"ܧM�K����7�S�Ĥ����1d��D���ʜ�c=�����G����Ճj��+a֛0L��T��_]PZ�[��Ӏ~����v
2��y	�9�E��$��w��Ex��ˢCd�튌h~a8��	)���u�xU[c�+n�`��/���cZZׁg��TB�'V|�>2��h���9Q\��+�*�g�_��������:@2׋��0S�-��d'�	'�~�V�O��������*��/���+V�7;����eI�F;�j� �);���FOC��+ޭ!�Q�٦5���}�(gw�%Jfk뎫��ON�-�P�˪Ir��^.2i����5�����D�ҏ)�+��
hqDD3�HGn�5��2��zG�Ƃ:<���j1t�޽��k���6�P�Wq����e}�9��B;R��U������� S�f�I7M���2�a�����i��O���2p!��9?�_�af�Pk�A���p[x�2|�Eӹe�av�v�w��c�HhD��$[H?�Ӕ��� %]B���P����g@��`�ч�M>�� ��4u94!*�_�m(	����q��(�q� @1 q:�@y!bs�V�vUi��j-#����
2�� 3N<������T �+�S,�a*̨�"Ł�_�	�t:l{���ʡ�y*O�%X"\��7�㮥_K�ߥ��4Ҁ��-��p���w����+0�9�5�[�l��ݵ�D�0��S�~I�9GTWa�d[�q{�N�m����?�ޢ9Z��%'6���,���@u�V���5Q^e�E��WJX`�!i .f��;��͜�O3j�Ka��Z��L_�F�k�'K_��B7���"j`���#���&Xdz�4q���)%�P���ԯ���������$���ơ~���I��|DDz4�kpS�n�ع
���I�m��3�nXН4��٣�Fvc����:`'�n� ���t��6�y�U#�vM�[2�+�f���wM;�<�Y��ߓ!XP�6�W_'#����^�f��k`��Ȩ������ ���=���gc6,�}���J�����4��6�r߅9�M�/@�x7��x{��A�Z|E��h7���f)B=a2S�@��ĩN2��|���(^Ҕ����G���?1/�C�ݑ�ԕ�R�.z�܅쎧C-�:EB��@��ðSY�'�w��8���'~��U�Bs&-�e���!Xj(һbH
�^~@6��uFn&"�i�w�L�R�������L!��Ґk��uPT�0�lXo��u���H�Q�ء�vB�A�1��C>W>�/�JX���?uGj��K�G�cv�K�i]S������N؍0�!�������҂���4)��q�F��{}M��]��N�a��Q����������#U?`��˝���η�cu$M����	V�Z���xr�C�(��o�ã�L��@]�s��F![Ԃ�Fnzn�@�.N����T�f�E ښ�x�&��%E�i��.��Y���xg�%y��A�[�;��m�a'��ZV�w�aO��\�8Y6� *��r)��x�/���R_�N�,�Ѳ��H���>��~� G��֐�]�ث`��ن�4��k�p��c�h�zN�ZJX�	�X6,�6��}o;T���Eޥ+�W���:H�ʩ󎠒��+�N��HڱhΩ4��ȗ��h���1���K��3�����I9�f�˱��m�?-���m/a���0�����nRBR���ӓ�����g�r�`�b��@Zt٤�ŵ\�$�����n_�Q�!��N�Ҧ�fv��a���(�	� N�?yy�@�e��̒���د�6fT�U�D���Vl������u���z�
��ӬdG �w.9ks=<biM�������7���G�E�"��+���	ڪY���u3%� �g���$���z�
�LEZ�08�fܷwo�d!Erm�*ɢ}s���(� 94��+#��D��s˽����`]s~�")����Ʃ�?��$�Xl0A�͋�:}H�x����ب��7��e�J���`���XZ?5'�Mi��6��z��nd6i�p�(eDp�\]�0���7�u)��$��-�!�(���"�� �p}�u��83,�(]N��-�/m�J�/�����,�|�(}��Ԑ�=���U����������5���鷤��M�~jqv�6�������{�g=�i�I�����԰V2^��&M�����L����Uà�_�`���$F#�C^5�2��:��3Ppqk�%�+�׳񱤣l&v�Ր�*���,���K��H}��!��Q�m�	*��`in�l� �h�^��BO�*��.;�~ǯ�i�hVI	�M��\r&S��^�w�O|k�̬�#t�j�Nze�}��w��i����x�1���}I.���M�o�Q���ɻl$�yI�tc�hZ,b����x�S��ob��x�LL������e���p�s2l{i}�(���%	��,M���8)lt#�Ӕ�QUH���|�'����.�(���1} B��6�}���L�xm��ڭ���Ҋw��U�2��@��YkV?s�^��>�?׻����D
D�Rh��J�zawL<���?�����"d���Þ/r�=,q���3�m���y;����v�P�[c��I��5p��qi�A}���<��:�$���"K�����jU�>dE�Ϫ�Ycm̖�F'	Y��{r�l�u]%�G�iM���1-Ҟ�y�0W:U@�0�%q�\JK��4=H�s��*��:���
��ӺD�����a�2���6S8���
���}�qށw�~=�[�
P��Xw/�9���^�~�>�"������u�����<�4���w.J��\�[~��-�%�`��M�̿��l4��jH����5��a5�����d� 1]c�����6GĤךax���D{v��)�l��{`��$V"� �n��h�ʒo�ZQ��+N�{U����G;��J`H���H9��ZN�3G��gOl�q�+y���vrd���<99�J�T(���e�9`'��`�'=�Q���Pɗ=t��Kd�2�t
�>�mǒ�=	���(7'����Q�f�m�߻�a�/��z�)��ҡ�z8�܂6�W�^��gH|7��k%2d�����׿��ⲻ^G���y��Z۴�}'�ؘ�~ޣ���晊��ϪH���U����\�~�Q	yQ�U�e��&9���Vq�X�I��s-ݲ�5 X�.��?����IhǗ�s9����kRH�ʺ[�
;��/��N��E/,�)^���"M"m�CيQ#4���W�p����ԕk�r�&���f�H5�$@$��#h�`���Xi�QVo�;̈�#��l��ԣ��wg���9;X��ߕ�o��H���	�36���ƫ$��C�2��h�?�n�S���1����t`�u�0�i��<�#�J��b%�q{���_�I%v�q+w��|��K$��r;��9�Nƍ��,�V1]���C�CS�Ϻ(6����&rb�]%9�6�?���@��{�}�X�࣪t�lSE����oH�$Jɀ�1)ɛ�'°:����&�#���|��Y���q7v����´u?5�!�6�v��in�����nw֘�Ӑ��`M#O�>y��k�U��R'���Q�\5�G)?0�tq?��2�[���Z�m�+��s�ny�?��X�Z:}�g�2&��,;�8d���o�����9�B<�˛��"e��#�玳�]8M�)�;bX�I����|�Vͱ�$o��Q����>u�����_%�>�����ވ_�s�l�N'�F��Ϟ7�'���<5�"�ɭ�@m����N(c��R����~_�|������M�O0��_�	�!N}�U�x*Iq�}@+�TO[���k���x[�#]��c������|*:{n0���G�.���?V�W0�'�:Je�kCY�@���k��</J�8�i�<�>j͠e_Ea��݆D�q�EY��yzMz��?,�s�6�b%�$�~��A�Q��Ẉ���N	;PY$M��d�y���Y3�&@V�.��V��n�f?c�fi�����ۃ� �����(t?�#�\��W����Qj�֋� �-�8��t�۵�ߙ��ʼ��V�f���d��r�"b[Ц&��̇��ޡs��
��Wc9,q6s�x ?���a#gs���g�9��m���S��jvL����
#�����+�	ri�¤��2�#��oL7���r�-��ԕA)O�K�>YNf�#$7n�=��	���6��]�T*����Lc��m�~����2�6�nd��Y%}���
��q� S"�e\"<N��qe��e7������f)��#=�nv��D�l��c/e���w4�#gBE�RA^d�>�K��v�߱� �'�̄�ӓ��_�2���2u,�MwC �>���K�����'�1���J�B%.d�}�:�뎨6 m�,"8P��`}����N�A.�z��R_����?3em<�F�`�"L`���g�颉9�%���h��&~�@�̙�rv���s/�8�	��Y�WX��GkmA�2�nV�}$�����uv]��M]ޞ3�e*/���/���H4k�+k�l��2����b�����x��y����9�f=�� #nm%jA�����աP;��u�� ?�(�?��8����.q��hq�Ubo_�'�t����	�(
��I�6�����1�ѕ0+F��؇	��K�uP��	��P�WIm����%�r�]�I��x����cXnZ���@�����L���cԲ��&�.�����lZW7[�֪D��]f@~����O\g�=��tTNUd�޾p?
l�6�~�)��Y�h'	^]99_�Ij�h���#�������_�;ͻ�D�P���?5�8?U�v��ݾbzW~eU�[�6o�M�X�ҫ6���2Y�Ғe��w3��Vp�0�u��}z��Ͻ�ta��O6�"q6VGb��*�>v�zd�6��B���fE:��6��5y�@b���E��/f
<�E�� S푊�pG$��\N �^�6&z5ܟ��Z���cv�,>�)P��Nr�j�1E�:���>]�Nmf��U�)��j�dO�dJ\�(#k!t,��P�; �[�"$�V�/�r�*���`�*b�I	��������M��c;�؝�I{_�1�7-�E�W:��o&�}*j��6�nH\�L�L�e<��%ю����C��k���.������x�HZ7x*`���À�A�c;���h�₿��A�~�1Ӊ=�W����5���
f����l68��)�e�Nl~Ļķݷ¿�����k�ZD�e����"���/�ҷh;g���9@9���4�y�3�j�8���1���(���+?�x�����on�܈�o�-��2�}�x
�&���N����"/N**�L�zO��<����V���g�E���Z���S��T��z�|mq�R+���)�2�(��[���C��Ƌ�%|F�y��������^�J�MR�9a.2lH�k5�ee�_H��1{�֗a�;fJ�٤�s����mf���+��`���֪"�+���
���^	�,r�w˶_��zQ�[m����6�Y����%��Q���*����(�Ɛ)������`���c����Q���-�
�wCԙʖL ��BK���pv�4��C�VV���.��|��.Q;e^Yx,
f�ݶΪ;�sͯ��.0�4�D�}��g��ö.\MO��������"G`��B0ADy�-�L.| �0W<?�u|2*A	\)x��Jn��?f����k��n��u���N�N��x�,�۸�����8�r��qKs�T{XK�Ga�ll���~ӏ���0����g�&:�D��J��S��P��\���k���ȉ:���m���9u'̈́�3�3nqۙE2{�vn���x�E�%&gj�F_�ŏKb��ّ�y}X��ǷP��𷙭?��̜�b�T�O�i�n�h��,�cm�p��1�=7���s��O�.?co�a���LL|��I����=�0;k1Ćz�ZP��x�fW��P|EV�yw�o�\�!F��,:�O9;�U���twf�Sx5��tx)<�A+�!�ݴ�z�r8f�I�� ��)��l^=�:���.j(OZ��o�S�p,�.ke�.�6ճ�R�-e����<��h��2 �&Lu��lr��Mr����d�>�����4��g�k�L�������/&�rB0�|��>����q��ڴU�EI����EZb�}�$�lY"h�Fvw��G�B�0����!b-K)�( P�vqÊ�ɹ���_�2�$���](XP�[�����d���Aʄ�95��lҀ�Y��ඬ��x��!��Db�������P���Q���"�F���P�����kH��r�Ŏ��T��%�%6}�������>���C#��)@�q_� ��j��?�;�(����M�.��+�c���1(aCE��(U��w�e��  ���>�}���<Z��ɸEp��S��dsP�<���!�o���1�(sir����%�t��p�W�$GQq�Zy`�`�Gr�c������Y?��t���#�d°�e�+3��2JӰ�Źa�q]B�����U�~Z���M۳�ySV����+���>E:����І�RB�;GϷ�eر��P�ʳ%����蝞wc�����b�ѯ���GSf`�=01��H}C�|�&,�G}� [-��5���(i�IZ���̸J�6�����!�ј�iDc� ;����N�D�(q|,�����h��}i����^�"�ƾz� �����1����D;I^�(�t�Y�u��b��.��αE�ix"��)~Pz,Ʋ��`��\�|�r2)H�#Qw �I_d��c@�����a� ����n�?8s����t�1
��҄%7��U�2asM)�4�#A�I�绽�u��{?�	QG}u3��t��	=�oy(�����8m'�O!i_���1)���o���V���
�Oꭺ~�F�z�=A�#ܧ ����{ռ�+�;ҝ�s�Y?�F߿�����vZ�4����Ywı��'�,Řz�JD�̾�[���2�9�G�D'��)��s�cpq	2���\ʵ(��|c���=��0ꕥ HU��?�dw�3B�.���Å�a{�B�;G�|����������{i>A��ʂz3n�T`�����Tm� ��1tT��-�´�wZ�C�J�Ew������k�����r\���J O����Lr�m��� �nX:O�N-禓�2?>���H�kT�^g8���`�WB7(4Bu���d{e��̫I�7d��\�/
�د���}ii�jt��c�����O�3�je:�! xY�7%X��fŅ�	�s�������&]�o��
�(����!^T�0���l &�{oWJ"��BX< �\�ͮh
�4
� 7 �rƹ���L�,Ki��_i�D~��)�oy���;*ng k�țRsx���b���M�^w�����]~��L�D�]�*��D%,�u1#7ڕ����t��ǁz�sN�m�)M�� ��8�]��8k�L8��_�[�Oh� DQK�	�%�G?����Ԣ�U��=5n��/��C�:W��&�'f!���2 dA�0s4�.�b(�/���"Y�u���E��Uc	�LE��ty�a;1NvO����.љ��"���h"V�
��~��6WϺ�FS�����#8����s��jQ�'{�t���*�=��=��&q/���G�!���O��Y�����L���}�����R�Ce����':�/40ybe���3!�A���Xl*�{���};܉���/SJ׵z(F#�e���%ڌ`1�ty�c%�=I��b|x/ۣ��"?����tv�UH庛��C>�B{aN�
u4E�#�9����%"i�֤#2���gI#�rܻ�?��-�z}�(r��?�v:.S���z�)r`c������9�,⁷8��%M���H�v���L�^�kS���b�(�4�>7/�rvu�)�Gf	K�L��C* }��A�[oG��(�9~��>2��̍���k+��/��t����-������8QA�v��I���Q��&�FɎ%������(�C���r�J�A���<g�c�<����E���(���A~�}5�iD�Ʋ���vp&��D�f�X��V󑦯�W��wQ@�%\$�`&�Q�����z�7e"��7���E}&���W���C )�� ���Z;��ߦ/[��%pzC����Ax���}��T�(%HY�Dm���R VG��a�d�CN�$�?� �=.�S�ށHěY�I�<�cj��M��z�5eU�2\��&iX	��)�/��BG�X��R`�����R���}5��5��*�������$ߗ��  Ϙ�f�}l�S��|ޠ�B�i�L*���h2q��ʬ[=?��z��F����f�B�ia�w�A��N��.'�����+uN�Y�A�c��i��Xĳ�tڡ��C,E�s(qO����V��p��=�q'O��X���F6F>�m�5| �7�S\z�
cNpglT&��b���e����q̑������7j������!4�G��˲�p,d.�O����n&��*:
8==q/$����߉\X�/�x�VHN�� &����M8��5,�o_�T���ϒF*aOTH}5f�2	�=%E�R ��*�����t+��<h9�:t�8�5�$���|o��W_�c�ؓ�}��"�x��!P��{p|�|��y���v@\3

��Z@�˃72��!�×s-���M��T����ė��僚��������@��,�0�(�"#ɥ�I[�]#�e@7��eLMZ0��>3��$`��~��?)u_V�_c*�&y���x��R��Xs��R<��`mxT��T�<^�Tnf������R��+PQ���>�%��[���'��>F�`����<�$x?�1C�K=8��'m)ۄ�4H~P;��q]��|�Mjׇ��C�:v$%`��+@z�����i9`��CU�ޟ��_���v��[q�I���X�M���C�h������|����+Q�92�,N�]5{��?� �}E��8�Ebi����jZ�|��m�^ �Df�/:���'�Pc�Epf�߃9𽂸s�F�4�H���y��4�S���?hJ=����h�
�'!(@ )Hh-�]�^�f�2���E�(����+r����;m�Ǚ�n)5�����xy�� 3
�y�#Mx�m�e�z@�ҌK�u6&�{��I��\�k)TQ=����]����%��O�]q�{������:0x����z�]P�bM�P�5 �l3���-�'?��]I+�N����]M->�{�$���oRJ��y�%�+]�k@���T�M���gj�F@;6S� �.�o1Em��4J�|��J��8�e����.��^���;
�?g���<���;�{�i�B�k�x;m�m�s*)�˼T�W)o�{��m���<Y�׷G�[@��H �Q��(D���$������?p��w�HY@\�V����W�W869��f�P�֗j #���R���{/	���*wn��N�y&(2�?1�r;��a��g%��&�`-��P=ޅb�6A���߽����[���b�|��\oi.����L$����!�w�G�/�6@������c8ؠ)�߭fw&#|&�V�ul|��e�a��/�	�N�3��Z����2H��)y�.6���k�o�����q���,e�QR\���j	P&���.��͠J=�ڽ>R�F�rU����l��C�Gf��ֺ��m1+��H�}	���W���N��1π��RO�rKq����=�F����7X��E:`��}����"@M�Y�f��?I����94�䤞G�(��³���KoW~���]�wg���?S�x��o,ڣ�P8I�,�͍�	!��O�u\��2T��.����N+���M��k��(@�҂C��hx�K�*�P��a�09����W����^��h�C�v��U�@T��C�y�3	Uo�s�X4�DFݦ���v���S�({��jbi�X66�&�X�d^V����gY\F�z1_��߈���	�*������͐$���GZ�3�O] �϶��r; ���y�'��򒝿]l㠨<����t<����J
1����=��8��p�׋���e�f�o|�]4X'PtP'S��#I�ׯA�R�{I���x�Ӽ/j���.��1�\^[w�w��s���I�ϒq_��P��l��+�k� ��~��n��`2��Jx0������S�����Q�X��S�ȋ�o���"v6'���)�s��}�Z�3�:�[5�������%�\/&���S�zl\Mp]��ي�y 6�h��������y��;)��.l)�~���[D�"���Q*�3AF����Z��EQ�<�9�k��rpB9@�� $�2Fl��a������c~��f�z�70�ӗ;fdO>D��͂��Xp9Z�N=��iLfqǞ7��G���Lc��',���H8���_j,���eW��x� �yM8)* �>&1�s�� h�n�R�Dm������@����%[B���߆˵��=�,,���@<���]D��W�A���1D��&Vl9�SV	���VSG:�dV� a����@Y+N�o�f�+��&u�lM��+Ǧ��qz����~�2"_�֗z
'�#6,Ms�FQ@~�~�t�<�%t�WZX�o�DE�_(�޽e�#PM2rbv�~��A[3'�/�	1(�?���
1�fk�m��嫣�/�/��$-Ї��9�^����L�i��˱��$��x��C��N������Y�D��EM��/#t�4�,�`&�h�>��L9C^���^�*�3�sy'�
��O3�]�#`+�_{{��L�W����CnR�'�NЋ�W��i�%kk���U��f{������3~Ľ�z��`zo�n/��^�~���7R����A2Km�#�U�D`�������=�����u�3-}��T��V�/A���ܚ9zR��Q��vvt�Ý��-D�6�2�ց`S�;�̶觊���dŢ]rp��hk�.x')q=nqX�Ձ�z���i�'�^ߕ� �Qi�	F<�L�O(�C��%�Tb�m��[,�ff �̈\Dc���|L�,8�)�B�e��O�����5K��k�"��۵�a�j�Yj`sH�[���H6R���h����n�c8�P*�*@D3N���`O�vߐ�����rG����ڒ���b�c���S��9
&�»���4��rj�Rv{y����䇇��"(p��ю�bl��p��B�A�D��ʀ�����J�YY3���}g~��R���G���kU�ѝ�-���=�Z����X�m�cQ�p*L��D��*�Q"Ч����ݧ��V��c�>�D;.V���M�?h̍^����,ɥ�l�\������p4U˴��VV�C����A��-������{\�bO�����y����S.%߁[�@���?�t,[A�WQ%`"d��j+3q֧8�
V�>�� ���/_�C��~���A�Ub �O$��PW�a� ��l�Q5�{��4\#V�M��@x��|W�3W�tI��n�Q��	�i�-�a{�;�u���`֤#דpԫ �<�*�}�7�M�NI$��=���u�E��x^����c^��k�8��fu��w�?�S��~���<Ju�ο{W���T�辢�&w�<��܅�!HǅAЫ��;�#b:`e+�l����]���c��˧F۵0*��hN��������K��a�W"�F�	K]��;E&~��J�z�i�Z���@X���:8Uwg5�W�P(���Bv�@k)��C������w�_��Q/�b��R��h.-��x��Az�D��pHd��_������H�L��ց��f!��y_wRZ�S�)x>�"��#u����W�`z����D^l2m3��%����`Օ6 �6ڌS��0o�ה�1�4N��0��ӵ��K2���J��$�ɩ��UJU�H偠s�Y�F2}���^*��;*a�@ 9삎��Ʈ'�RY� ��jzvPW��/�И�C���$
h��1,e�0�*���`��#L�BΈ�p	wi�tW]x��;�!�
��Ca�s#O���a���"��L�h旵["�v���Z�b�����0'l,{����J!�H���e����F(��I+%\Er��*i_햌>Iu0�&�1���cVU�Y�~��UBcf@��fs�lD_x���uC0��պ�.v���?�E>-&İ��qQ���vG��V������M��nဟIn
:�����N�t�T#ΞL�t�ӡ�+	�R\�[�,�����U����7B��55�/&W#4;9���LҚV旺y 0p�����VC=fYK"�ւc�Z�k�Aq���0�,��I�k�ǃA�d-��t�7_�S��tv w�JY��u�=�S�+2LW���' !c�xQ}0���\��S��o�)���z�ES:��xH�,AY�ݗ�(�u�����N�������.2 �v�g���?ӝ�a%��ft�ح^�{�����h���h�:��:i�b�"�9���cD�LfN~�+W��#l'#?3銎�FK�;v���S��-��\LӺ�k֙��i�Ь-h��/�\k��\�����:�M�#���F}b���`Yl@G���p*F��h�߳w�O!����}Ք��n�I{"Q����%k�й���^�
Q=���,q��d��SQ�����,i�����e ��pQHF���h=Ip�X4Ղ����T� 'U����d�k~6t�b5!�1�ߴӄ?��up>t�X�ֈ�Lg�
�{»�����?���$�e�<OGv���1DT� i�8n����Nj�?�I-��"�(�H�J�tS�_~��<�Y?��^0+2f%r':6��ծ�/M�;������BЇ�d�h��þSq�5W���6E��P��J��뜄�S���捥�l��|�G��7�A�(�Qa����]V'`�/���d
*���3��N����Ց�S���]�5�L]�E|1����]��;��@���z�)+�U����{��y�N����(M,E)��jc���v+�>$�
9X�6������H�f
�z���,�>ez�{��S��D�2�,Ȗ���z�N̔���ᾦ�)��<I,n��W�kE�	.n�����^��7y_DO�(�>%�TP2�cX�q'A���Ψ��+��m�D��ב�J �	�3���	����yx�e�?�VC��W���>�ɭ��Fx�+hU4�6�(�$2h7q��[2���RE^�LvCz���3��w�޼@�����ɦ����u�R<BlS����a�3ȡ�C�v�|�� +)�VѠ"��Gw�.���v�୍����@re,�%��!ݳ�>N�v�)��$��O�M�Ê$I��k<�85��B��V#
�,>>�R��1r�1�� ���3�u`��\����'���ف�E��5cmTNS!0V+\ϱwR��mk:3IV��1#��Y�2fEItz��1͡(�_泇[�%,��P9�{G֣+`:�;�6H83z�ki�zr���VD�	���g����L2߄m0A˱[���0��Q�9;ԙNo�}W�/n�>oh�Z)�S�)�"���i2�4T��N�V���s�����o�R9�M��u~C.)I��l�Z��'��.t�"�����+;���ZeI,:E>���uz9Q$�	6[z;Q�z.6)h�1���t��.~Y�nV� ܘ@*.��T�i�-[S�&�ζ���uЉj��O��K����^�'����!��,<�!Gq����k�<+�Cϗ=�@s���efR��i�,>���P,2���l�0?>OF'��P��������m�S��h�. X�(kli?�쏶��,���G���-�4���$j���{�5}5��X�M����p.�B ��_<�urضN.�~����$+�v����
2�\�H�������g=��k����V��X��L���5���n��֫/�nZ:��5NVϝ&\1_�USVr38�2j[��z?:�^���i�XQ�	×�sHm��X_@Y�7ꚄE��[�˼2��@ɨ����Vz��r�z߿}_��!|��|>�Cy��J��3N���1K\������$͜��X�H2�h��gȴC��B��5m�)1�����Ԉ� �Pe�b�;�1�� ��.�!j�!a������N�#�幟�ڤ�	��O�ZMfP�A_$�s6�+5��[�+�t�=�Nn���qO����RV�/���vW�&��u����l�R)=������"ԛ��uha%Q�o�Df���`|h��f�D�	o%��@���$�
=��Ϧ������N%I;��q�`~	���%9t�.�m8}2�{E�Qh�W�.��7�fK<��\넡]�԰��? �Ť*��3h��<�g��z�2B�J@3_ڮ� ���t���e4Ig祿K�����M��Ѓ]^�ѓ�N5��a��W�� 7�S���"�ZQ1��h�	�fK�������	�rN)��JQ,sڝy�}�;,�F���?W�N��<�c|ā����$6ʍ��ɲ�YЦ��o�bz�=�ѕ�/y8vó�E�'�44]�6���ȥ1D�1�&�L?�m��D����,_�rs���o�F25u�u��%J+��!ϫ~Y�?��	�J&B��Yxπr'.�A�#�d�����G�A�h]���K5�G&!5^���^x�����jG�?j�@N6 ���Z&�j+��,ڮ�K�a�,&�	�X/��������R#_��M���֊�#Ϭ�/E��50G�M���������"?BX&���8�G�B��ܾJbod>��x�A�QJ�������,�,=B�͞R���M����'�qM���x��Q���^�t���_d:gR�N��/θL�I;��Q����xew,�W�N�|�մ�aC�.��iڡH=q����f���$�D���:�2��a��`��)��,+��C���B�V���y�I:Q�zz���k����(u7ʊGIQz���7B���gxɍ�0�@��"l7JF���3O8��ͱN��h���rv������EL;ܛB�A�Ȳn�F���%�4�ԋM�fo���p����px�-0n����(��8i2�A���W�^���bw��j���\�_=q,g��J�G�W�R�-`q�Pf|�nb$��TO�碱�R������g
^�R)� �_�q�r��-�����` �����P¬	؅�'�M���1h�iJ"��F�l�h��8‰�=}������e�q����yM�{�):�I�Hp/�6�5�x���{��1h�B���K|3��?M<T�jE\�b�OW���#ң~��,��}��}�	G���)	��b:���}Mmrm�-a�2��7=�/_;;�"�@d�۹�|�_�Q�l&
�Wd�*cĻ���� T�!N�����Ĺ��� �=*��χ���Ѐ���+ӎu���<Z%EbP�N��w'� �tds�V�8�%�6�"��C�Iho�x�CV�53�P�.�GQ�>-��r�x!�FF��l;1s�2ʷy���~+�:;GNnL;a�Pg @m~`� �{�Z���E��O�O�tט����EUYbRl��iZf\��6���+����"�2e���x����5�6p��(���b���72t �����YC&�He�fK�g��2��
ƾ��ªn�����̪�4�AVs���+3f���=���E\٧Y��)q��19�����G �T%���	���0���1�v��U4�X�"�bJ5���!R�m�b�`����Q_n����!��Go�&�kޤI7�	ʇ�?���{�8Iiˋ^��`Bō��p���}g7F�vy]�^��5����7L�_��"`��{�ԑ�?�P����pĉ\0����%S<Xo�V�����OOLJ��Rt~?�E4\49�Ȁ�I�{T�	a�1�y�M�.�5�Ҁ*�}�s<u����r���!��ޢ:R]� y�Q����6J`� �@��H��4��JƜ�����ݨI��g�[<�aq���� �nmb��;��fRs����a��n}�ɜ�p�sB"��O���w�s� A� �wZ�5��Xɒ��P	y1�2���}���5�`��^��s�/��3L��>�G��Z��oz����M������#?�HtF'�A�6�3�$Ǩ/�&lr�u�����}����ԍH��-&�%H^�qA,��̟)�6��r�5��cJ��by
�$�S*�N�h����K�����&�����{�1��i�����w�f���=��u����J��7�}�]=�����_�=�47J�'�Չ�Ph�0{��U���@�;{3��a6��J;p�Ep�'
�>�����,$[`�5)���u`��u�8���`�v��2�F��M��R����Ηi��`�Rɲ���0@�tς��)<%� 4�~>�*�6h�':��3j?��扨T���[�ZS�F�H*�]�g��Lo��8���������С��:�Ty�0�p{�Ad������"�q�q���������H	��@4?� X�7����azTh�+�7e��:�\����w�|`5�]6Q�~*�����`�}牺0[�d��+�aI��R��]C�������V�b#�i���]�jj���f����+�e�7��$&_�Re#�~�r=�V:�H<Lv�I�L�xVV�]���O�A�<͹=C�r]h�	B�!�06o/{���Z��{fJ��L`
��|p�}7���-F���4ݝ��d�d�#J�>ȹ.G�P�fjd�ʳH���U�������S�_�T): $�
�n��}�^Vp"��餑�Su����.��5����5\<���.��-�׵��E����D�����b���幮��l*��ϛ� �Yg"��h�ՏB���K�����ʡ7"=߸ђ�+��A�ǲ�`�C�8��Yg ��Ӑ*����K֥x�9}?�Ix1�~)h^+l�9�Da��B,��(W& T�t��~h��lnjo=
(+Y���{m�_K"��R��Lc�$�%[���������5��PWViM��u�r����]	}]�i� t(�A�e���r�q��i��2���{��z���Q�-�q��:��6�8PQ�tn�_	�X��q���"2������}��0���M�������՟�TF���)+�n�? -2W�EZ��ƨnp�Sb�� _�J7Q�I��<��w��
�Y�=�u��o��7�L Sp�Xr �~� ��
xpc<]�
`A��@2,�����+噰�.�R��9-� F�(��AEΫ��)�9���%���ƹ;|5�^~�qI�����KH�8��ݎQ�Ӫb�|5 �֜���i��Ɂ��=X�[�k2��s����L��]6đ��7ì�����i���5�?����I{b�1���^	�r^2��1���P��BG����=9	BS��ĥԈ��/��N&��������#�L3�m`0���4؂�;Ћ��ډ�<���&�"^�A{���'J$����[7��įy��=_�
��5]�Ve���B��	.��P���Q<J0Id�|8NV
������#lv��M�`B��0��͍s��!p����4�:�h��&I�~��z��[8�B�H a���ԁ��mȟdwy���
_�
e$�j�>�b&�4lI|
����	���eZ�_� .�V�}��-C;�!F@4�]�4�ɿb��&�a�Y�w���b���- ��̨!A��C��C4"�/��"��{��Y������q/@t�V��?%���2ơ�)��Q�~��d���k���;��Ϸ��sįC�W�'���$�&�?U���|�S�;��c�G���G�1�㖖�.�up�"H��P^��@�oG�������r�h5��췘�0�����p�K�|����^��^��;�_t�V�*��J��J�V��R�:���5��
�go�z�}s�mza�qN��5�M�����2۶f���u��PL�+H��d�mF���ܧW6D]�����^"iS��rA�X����z�j۵�%��9_�Z.b���c��iZ��,��f؆��4ʧ!Mkg���-���H0��6�e�x��o�϶�QҨ{���/̟\�5m�|	�d���G}�=f��Wb!¸٬������g��ӓ7���RI�g�����i�D��O&�p�����"r��9�۰�<�ep����<��έ�����t1�O{�G�ei�w���Gr��݌�AͰ/�͵T���J�&��G�E{��zN�M�J�ƺJ��L�����s��#l���ܯږĆs�ӄ�~~%�.����NkSǞ��A5�y\%:�������0�v3xM?�n @��r����~ �{?�3��l�'�AX";\���bTфr:R�l���>����{�W��Y�u�[uQ'��u�{���Q�n��?z�Z[��b�Ĳ�L��\٦b�`�;.��"5ށz<�,kAg��c�f�\>�p���16|��g��;�K@7��g���[�?�F������BS��ί�@b$��L��nܷ���i�تG0Ĳچ�
�����Ax����ci=����j����A�����-o�B*Lܬ�7��ϑWp;��X@�US��c�߶v�%)����4��	�vÚ������/����S1AΎ�J�������6��D���YI����N�Յw�VZ0��/�q��C�~^�c�߹"�{ӹ�|"#���v�G�F��N�Rt�BiY�� i���Bd��
c=��\���8n�*���ғ�Y�a?��j�b�hsJ��T-ۧz:�:<Q�@"���#��Q���$�R\�+b)����������Y��\PX��� .[�$_�D$���D�l��v�h9���I�� �?��ICB�R�|/g��qLA*?g�=lx�Rc�a��o��]B��F�}յ/��[>�6��Y����~ѝ�g�-���bCf�r0D�1n�&�|���A�-�ɿ�o���EvNch������w����MZUd�1hm���w*��g]�w��3�p?c��XLVNq)܉�
�>gAg&��#�Y����-J.m���7v�	��X>�[(*N�m 5��b�ֈ�?<�� �I?�nxU��ڇ��(�gڸ��//c����z"���[/��C�sZKd�BK���i�|�m53�p��hi	�/����a&�~�mrL�ie*ue�L��y�L�J��SQ��#J�ɞ�����.J�[� �{�]�곒C��;w�Tl:�+;����Ya��|V�+�z�[s��Oy�\�����rE/��WFe��=���ӗ+�Z����5z~�� ƌ�4��X8 []r�`��`�=\�M���׋E�|D��P�w��5W�_��T��N��n��v���ڑiӹ�6�4|ǧ��CR�^�#�ϝ������x;u��S�d��h����	���T��s�<����t��N�x���fx� �5m
Ub�*]��z���yi|i��W����+���Ȫ�LhB�a��@�K�`b¢wLdT������Z#��VV��
��Cԕȫ}�﷩fQ9�XLl�P��l�q� �����.P�﹏�}����跘41AM�%�l�̃������i�~�;��@��z	�R��Q��V�&��ε��9S��XL����l|�G� ��4�<�6���?���+i��6���>I���	 �Gef�̽+�����M���Ļ��ao���w�/�����k]wP6�RL>w7w��:a~��<��z���mr�F��;��Nh$b���:��bZ��3�ˢ���͂Y?��K�a����l|yn]'�}&�P�yӨ�iz�I+B�O1���!.y&7\2k�9���2�$�v�J�lM�)�cv����U�_�W�\3������gy��?���aF����"���v���gV:�s}�OxfT�\J4Z�M���!��X�*\��C����Z�����đ�J�m_ �>U!FC�iv��Q�h��H���s_�m*����+�̥�	����@0�'^�ֲ�<&$��R��}��~�@&X�w�o�^�8�Z5y�(�Z���绁�!��2~�)������~�{WV���='Tӓ��3�gN5����Z�}�����Vww���yr�;��Ux+�L�?pK�!Z�����O���[��7��)����X�=�����ë��M�$$w퀩c<{�?����^� ��c���;vY)!�G�J.�� ��8m�+����>?�GB2K����1��	�	�n7+L�mŉȿd��I���^��s`B鉣�����G��EC�~�f�����" 5����C΃tK�QQ ey^7'yX�ׂ��1���Ҥ)�H�: .��W���i��8�e�����~��LܧY�p��5M@l�/[ޫ��r��L�����3���i4���?�Yb8D���D���Y�|�����|+\mq�[2ޑ2�\������_�pImϞp��%韖��p���� �}���[ۯ�c���Rv�eߞ�O��5�Sd�`H�a�۬�C��^�=�1�l��ܛ �O���;p����K�|�RG3,ϸF~����Y.���,���,P�Ǎ��?��n�0�̧X�*��}���$����@����+�����`�sT/T����Û|F��_��%$��g�Aq�DW���s��\���9�C�0�&����~<WG�c�向�b���!����/�9��Y:}[����ȫ/�_���7-<R�D]�%�D.�Y.�W`�0D��p]3��I6+�E��!.x^}�
�b���OM�-$lP���G࣒;�q>�{{}������웑����^���R��I�{y�=��Q���B`O��hY���$�2@������?>Fidw�f��jL����$-�I�l�ILJV���q0H�6an�*�>����T,�60������jhTG-��ύY�Ƅ-w8#��h�JӺv������Ѽ��t��^���LF�~����j�8�*�����;�d�f@���P�����c+�I�= �"Y�a�v���"?2�
��b�k��]�IըW|�3��bu��:�X���+�E+�
�d�c��;����mF�l��U���5c,;Y�N'�+ᴡY����7 2ĄWO�4H��FnM�l�@Z���̒R??���J��X�+lD�VkI�{����U� �O��`����9�;��Se@!�$
��� -�I�;?���LUM)�.�{ݝ�F!���ac4~��]5�s��ݫ�b�n��	*�A�pA���<k�@�z5_xkxߪ���1:aF�&J�m�/' �����I=��� ���fj��?���/m��+?^a�ҋ�'��ݾx36�lR�;l˞�2�w?֢$���
w�>ጬ
�a3�K-�$�-�w!��{Z�@�?�.�V)~��|��q}�bhp�K���\ĲK�Ԍ���W�D�1CўJn��z���W @8�іX9U��F���jíϰF � @���IB����7�/ b�|%��4�B]��M.�q�#N��pKA((3Jj��f��]6޳�d��6Wa#��j���q�;��ʋ�Du'��5����ɱTmS5�ؾK��ѵ$&�O�0��e��2 [fs�}Z�_&�a	#4�c��)@鍔��~����$���V�ݬU��4�N�5����T�nh3�!R�,�[��]������.��R׏�dn_�8VV�)�-!j-�`$�� }��C�RE�|fV�3�M"CL�z��b֡��[=���}����8Kz9���$��,�|(��D��������Li���Z���IJ�`�m-�P`�o)�K�+����b�t��u>5�gD�w䱻9r�3��m����,	�"F�G�H�w���?<�̈��b[j��J�g�X����d��_�� %O!��׃�:�zh��cN#g3f�K��CJ��*������A&��Z�+b�M��s;r�U����Gܰ�Ịm�6H�H��Ӥ[E��RU�qA?2Eb�[C\�^�:=Xu�PS'�͵�~e��:'
��~���g�������GY^��4Y�3R#-�ah�7,���� ���D�P(Wh��2V#�:`�mBҟ�¶h줺�b��\����ۣ�c�ݡ����nGvl�u�)���Ǳ2E4�	�Xi�5Q88(�ӧAk/;Z�z�T�\V:�i�)���hY���wRp?^��/7����Vt��/��Ru��6��*"gN4Y�-�!�� ���B���\,vwS?�%21Z�ɤe �;l*Z�&�7h,����P�T �ZK�dT{����̪�{V�:��V ,�\�J�_�8(�UҺh<!Fk� cU+��d���VW~E��%b~�Cj$�,`~51��8~ە@ą�����R)��#�I
��y��.ƨ떑O�:UX�_F���a����g��O��}Xx�b^tU���N�ؘ��^.3�ĘwT �Oq|{��t�tYR]���4�A�Fai�ʜs��	O��}�g A��lBf���k�ER�[��M�5\�b�Q�c�� Q��9g���9���78O՚���5�'���2�юG��G�] �W��Ѯj����G%�ߥ:�=l6x�q��B�f���=��$��L���_*`��t���X1�0͍�-�قm�8��*��+���߀�D��9E�Pv�Ԅ����p��N?(nA�������Pjё�9:+�-�M�Ҋ�|�c[\�?�*/��Q)�4̈́����V�Ϻ��0�,��M�v*���:W���j�	w�x���w�dμ����@D����~a�T"$��M���PF6J��VH��O+��T�ٜ�=����J�� pkEBo����Ӝ�]XZ������㊊�"9��E�R��Ϩ0��z*���Q�UD�4�U��Y:⼧z�ۻm���󶗔0������������TN S��'���g�zу��j.v�o�.��n7QbD�8��
u�c��&��*1�������!�E���y�)=گn�4,���r>����h������
��nډ5��< Q��I��*�Ҥ��]����O��4w��}�v� (�7���I-�����+S	1���&u�u��e0��uj���[��}��X1F��;a�$��e=+%Ty@�ɤt�Eyn;f�TF���S��CkCFGa{�6M��|׎`"������6�e�a �m�O5
p��,��6Ύ��@��͡uM��8��N8��x�)!l��n�*�����i��{rW������\�ļ�-�:����- x��r��l��R��5�j��yJA@iM�veP��r�T���Be)M1��Y4^~͛�A�f)��[������&��[��x�n~��ܼ锛X���Ō��yN>#������M:Ւ�4¶L:�c-����k3�`�"�9���u%�T���]����/��X�ѵ����0�*Ǟ3����;XD�|��H��X�J���p Q���V�QZ�|��5�3��k? y� ��V�&޻�� )x;y`���Gyd��R�ySk�"�)n�ý�)�����u
�r�n�O�yZB#&H���7~��������Ɗd��T'�c@!�Xm:(��;Pe�!�ģ�):H/�q��-Js�e�I	ܘ�	B�����M�=�1��9�҂�`�����j����g^���UEz����oW�M^���'�]'zq�3'(Ox�9��J���.�8�ޔ��8*���|��,���	��
��8�?�������ef���M� �t_ddu��X@I�e�R��˗Z�Z�~f$5�Q����v�o]�V��Җ���O��fxE� ��iQn��W�_���C	���_��n,�__n{�����H�'ly���ҥ��v���<�W,>-��oKP� ��A��*��O�]��B���2�  �At�,t�]������ ��F<s�@:�
["�(M�*���!jt�F�ͰL�x��c�����}�Cu,���F<��i3.H��4���ҒN��0��RiA��^}3f������щ4�9rbلX�[������-t�_m�����D� 	(�z�|�s�z��ȋ�p��nΓ��lbaY�>�����P ��m�V���>&�H[j_�e!�Q�<rni�P6����85mC\{��F��y����O�cs�q T��%�P��rϴSy;���׮���������1-��B�dQ�􁡅+(�s��~N� �m��V���������:˟�q�V��LA���@��Z��H�?�I�/�=�������"j��i�rR�q!�GNR�rvf�%i�e�lG�4���ү�ڰ:��Q�-�×��K�7�e߂��
n�����":}� �C�8!��xp3gA�rN�:P���QJDP`�#n�e�;$�IH?#q̀b��|���&[�������<z��	c�ͅ*��;�z�¬�`�]ە�?^�\�Dm�Q�#~�;dl+Xk�,�ׇ�D�]�p�w�z'-a��Mi患GpBG��雡�4�"���1�tt�}c�����w�5P��aY����4
��'��9��/թ=<K��$�G�P$Ȳ0Y��/-I�"��ἆ#>�&��;��J����-�ׂ�T����T�Y�G ����n�� 
j�4�e��'k���k�0L" ���� A��K��S]:�/._�6Ez��A��J� �� R!�уx�J��lI~����x��X�!w\�~r��1�R��2��Q�<��i� ��^e��\��֦�` � _�)�4��c��y�@��iZ��;�ʧ�Z��-M�ݴ8bN&��b�Fx��h��}�7��l��������ZИz]��=�.�7]۷���}�3Ej�}�!EgW��;2��5Y7�%���V+�*��_����b�ޡ>���HG#�e���]d�3�m�AVg��:��/�~څ){"���kI���a���� ��?������/�>����+�0�M� �`���t�7���l���(�)�����C���l���-N�[�}�Vtyڎb��1#,3����� �5l��Y�������b'C�3F�
5�o���*mT��&u�:��<�5��� ��=�$��e��F�F��w* 7�`Ĭ�kG}I?���i��yLO�/��᧵ǔd�*&SVk��L�h��G���g�`�RS��,���|l>�}vR��|LMѫ��Դ7�
b7QȘ��(���9�텮���1ѐ�M�A�g]�.lc]}�o����N*8�R=޴#��y�,J�ռL�
1�:�9%�!��s�v�EëKO�(]Y�*f� ��%�m<�:����J�6�M`��E}@��b�k��rO�F�bF��/���-:�	%l��LAqy���Ƙ+��k^/dm�e���%���W.<�彜%FR��cO3���<{(:�kz�;��ز�:��/׋������=ԡs�s�u���?�7����m$K��w�+1�A�x��y!_�`��3 �W�	*�T�N��s�����tȜ��*�� �"�fv��dZ���*Ko�d�k��%;��d�����H�E��4�m2�D.��)���
O -m��/�V���e�
 is���A-N����V�y���5��K��O�QGg�G�d>�<0�Ɣ{)�I#���D�wް�$���R���#>:l@��l����;q��E�+0���'���CLI�Gg�bV�9��:Q��ݜ����C�!��S�/�#� �[Q�pYk( O�A���?s���C��5�p�%��.ɿ�[=WQ���h^ �O{�)���X�}���^f؛��"uA�(M�Z�|�f�B7#��{�P_jF�&#Mu~��j&��U�50It�D������O���<j0����ΩK��n0�����hغ�j�
ձr��Y��m��],���zXF�S�ɱJ���yH�QjJ��� U���/�`ۿ�1����0=U{�JSUp���,w�$��G�������ӊ'�sn���tZg���Y��i�++8�� ���Orޛ��2�����+4�Q� qkr���)�{�ٰ���kt3y<οKif��O�K%P93u��W��}�bA�np����Y��ꫭ�j�E ��M�y<x!����{B^r�ьmc�Y���n�ll���R��K�Ըv��S�X��� �dy�/������\��E�iL:zv[�@38�\ѝl�4(��6>t]x�L-�.Y	���X�:����MF��W�f�0Q�5�*C�c��	�(D�h�Ϋ6�2S�%��%^��p��L�=?�I�#�9�fG;�	��H�\�5 M��$�q�ɩ�����K%���PE�)pj������i ���oZ��)vP�3�%�	~��oI=`���j�K׭�!_�/��O�Qďu��W�{�^��D.d�U���{�=.�[�4��+ԕ���i�<�M��!���J".MT}�t�L�&ʿ{|2�TiYI���끧�p����i|
��$���_��ː��e�%�Lu�<x�4ck����~���t���vJ]��9y�ݞS�F�������E���
�P`Z�{���Gr�Zg����7ZW�����`�M�%�����vnz&Ѫ1�U�P���ꞷ���$s��	�>(�����N�piE}E��x��Ķ�X�*Up0낧3��L���ySħ�[7m�X�]��'T	RK��#�FE�g��4�	�@P%���n��	��a�� �An��䂸�J�b�n�h>{9�X�b�7A6�%V:,դ���!�:�ÿ�_�KJ�l�>��ۤ�s(�*cpL(�$��j��U9����_�t��:<� �'Խ5���)9f������6��̤4e����<�'��n%��u�pfA�I��x�1[|���^�i�yL�r���T�g
Jpi��X�LF�Ux��T�A����������	���	5�`�i,tB����u��ؘ�Z�!���T�M�d�$2�p��J���$�G0WX�ǻ^I�9��u�LE�'G.:M���:�P@�WX�n(�G�w�����ά�∬�BR@��O��>�����Z�q�Wʼ0G�����[�l�m6�yb��ɤ�Q�Y�T��WfH�ΌKG��lhKl_?���jej"������@ڤ�V�1{dr��3!h�wEb�V����P��uɏ�6��Ė3n>�u�%	v���'1�Qe# �"�w�,��|�ɛâs� �yqig�,.l��m�>,�] Ն����a�.1�N7 e�}�!��e���s!�'M���nh�Qz��.b����h� �0��b܌��5\+=CѴ)x�n;\���/������wU>Va��������SWts;sг3u3ߕ�C=�������9&�m��hS��}�8����=�6?�y�>��a����:��Z���M��n�Wu+��mb�0D%U%k]����M	��٬�![�����s���`�������r��mSx�1xxh�K���TR�u~ō����y�.�jڽ�}�G#���8���}4��Q�f�=�?����	
�O�4zI3���@1Yq�_A���L��A���K�f�K���ݿ ���|͊3���f�����/C�$lfV�(����a����w#��}�K�1�#�AJDtĩ������S�I�c8�D=9oU�ؾ�ԍcmhi�n���vK��\彩ϝQ̙��p�,��]G�lЪ�,w�����U��9���TX���P+�@���x)q��6<��@���k��RN�ڹ�b}����eb�͜�p����KK��I��F.�>���O1;zG0��C���HW#���� m�WF�>��F��%f��=B�
�\Xc���x��.=��<�U3왟R|9F[
��d�k��xH���O7IKJ+�Ʉ��FWG>O��A�x�1�t��*rm���P��q��Ͳ�ϖ[/>�\n�T�j�Y9E���Ο�5�u�z�� �L���ϠR��� Y�K�Ƶq�!Kv�&N����VĎ�c�5i���"0��ۃ`f|1�ըM�0�Sf�ol7n���=\��i����WO�G��:��LJ�����`t�C%��u��/�i�W�5^ ����,e��6;��Q�#�FKZ|�����2��~l }pFQ���J'��i�.ǟδ�wS���nq]�QL^y��Au;O={Hŝq���g�8Tl꿪I�Lֻ�<�)h���㐃"���D~�v����!�w���1v�D<�㲥z$�b�6����o��;���q���ҵ����wZ�Q>d񋏄��S���7��q����v��D�?��^oB�՘��>��`9�
b�x�p`�={H ���!2:���Dm�X+5��B�~�s�q�|��ro�?��$�)&��B�kԎ���OF�"N�r���y}u�X�n���jz��KMT����-؋�����e�1Ϟ%�:@]]�y���фמn�P.�v*@��g\�����ֲ�P�b�d�i�4D��Gb��h�z9ѹ����\�=i23��'�+{=��s����q�g��<���-`��>#�X}(@�3��4�-B"ǥcy]�F�h�;�w/2*���,K~U1G�^��
a�ó�7�"��)N�& �抸��M�L�U#�e� =\�0L�̪в-��f(�8*,ik�4V[�u�'z65���.=2x�&����*�/n;��l�t��׊��9�a�c{V�mR�A��T��݅�s~oA���2E۫�O���@�	Wl�A�i;�;�2��.�T����YW{���0Qb1�$-=\Q t�Vr��[�dk=yj��������%I`�Pa�b��!_>��	�h�U���u�,H�B��*IHib��ݝ�į��+ꪡ  s����<�����,o���vư���m	_;�d A'�i�IL��%AO��i�bϗSں"yj�PŪ,�չ�� �k���-�ඨtE��}�qx"P�{��G?�U�Ι~2��#[lƐ�bm����v��q��2�q��ʺM@�~n��n��o��sx��ƫ8S>I���1 ��:�$�e�{;���Un,a���"��'"��k���N~_nK��ńq��e��8oJ��9�E��ٿ/l�ͥ�U�[Lk�<(�J�[b��f͡c��t�<����_*t�e����)��&ʉ�;��/JX������/�Q5��j�+���C���gH����D=���9;��P�
���A�� ���Ț΂��0q�9�+5��5NX��?~����T���`@�`�����H]^n$׍�]��ӊO�h蝏'�N��g�
��C%���R������}[�X]��.u�tN��{��?`T{��c٣��B[�9�|8t�� ݟk�{9�q���p>P�!8>.�a6�a�B�y*�Ϫ�䲍>{Z[]�.��!����Hd�t��=�~�ކs�+��hU�EF#K	���͞��ɥ�[A=�>���j��E'�D������W�u;��-P�������m7*M��%SZ|���GY����̞��%�*����>c��.��G�A�EZB���S{�蝑7@fR�f�ۛnk���y����n��
�*��κll�w�D9����6˷E�Y�K2䈠;ɿ�w��6أ4�"j�=S��:�Op��;�I0��GOG*Q��\�-S̽��Q���u*�F�ϵx��������ٜ�I�&��1�Ǿ'���-�ծpؔ��<���!�fP�H�_��5���~�������aL�1+�,Q
+�@��T@���e�%��]u�(�5�:��
���)��Z-�NI2�ZD��́�.�uϣ;[+�����i�3߲,C���� t�Ĭ���y�-&��m�
c�x:����yZ�1#�:�#����8	z*��E&�\Z��(�ċ��g|z�v0�Ur�;|&j,tc�z�V�3?����<�.l����g䋐��#gU��a�˭��Gs����{��L)�1e�c��h<nxG�;�Cx:�ท�s	��x��c��21�]1lfL�4���I���F�x�L��Z�L�j0�Ր�� ���z �QXE4m_/I��{8ݤ�g��c��;RB��.k�d�oR���L��L�8ץTl���P2`S�V|�� ���ל�s�Cm��G��h\�&_��K;���(��x���5��>Ms����;ξI,�chW
4�3�՞��]��~"Ot�^��ׇ�֥�G�#�A�Ȓ[��ZJ_ǁ$�9FJ&�q�M�BJIR�1��㺢_+�g8������1K�!�����1�f	��F_f[��w٠Th P�A�_�~��L ���79��o��s��Uw߬��-ry�I��X@�:�&�<� ��Ɩ��8�{�$�,����2�i%9��
���2�"�oۻ])ǢD�a�]Y�)��j���C�>x�3{��8@��-�����o�w��P�j,��k��i:�ϥe��˘���!%3{~E*n��z"7{Sʈ�I~L��&d�(h���)$��fI�5�:�y�@:���ױ���#L��em�S��6�t���֞�c����r,����9=�����c�ŗAl���߮%m<���mP���s��Sg�tk�f<�����L���i�w&���Qf�0E���u\d���>�����b��h�V�l9`�[�C�1"� 2+�=�؉�Vf�O~�F�L�����mB�5�?axxW��At_
�w�g�Y�ԋ=%�緟r�	��|����F�h)�0����S�j���������IGO��j$�)6����՜�ya\�#��;�{�nq�ߤDҮw�ks�+����;X�\�1���(�xx���T�1�4��3�YD�f�ј��-��
��]��Uv��8ZK���\���%��7�<�{�ӛ�}H,q�6�E�p��K7ò�#�f��
���oYNr�g�9Z��8Z<�M�����?��baܮ�]>��;��-D��>.��y��(=X��l�]f@��2fP��Y6/�HA������γl���h?��h���ֶ��>���R���g�\����5�����> �:�i5�)R����5�u�G��u�{��2�n��c�m7���^ �ʮ<#�4n�S>�$�� �2�c�o���%|�ʶ�+"�̃w�r���$W�*�[��>�F!y�-7 ������Y�zH��g��a�ٗ��Jz�k�@�x�fjoqR�P�<�n��������u�����-c	�c�+~��-��ns=֡9Qw�%@�]��%�;���>>�X3����gEe������@�����ғ�I}Ü��[
��'}~$��~�*.����2�Da��\�J��.�}����נNޭ��&q�S�]A)&���-��,C�{&�.��}T���Ն����/}�5�]ټ���2�U�׭B��t��jQ�rPF>
/H�f�F��BlC�.����{��)�#'Cާ��Q�Z[��*���t|�����g�#���7 >;����M!�v�2f1(���,A�	��V���r�=��`��F��]1�W+�IYZd�ʋ��N��l�R���v����?�O�O[":&�=�Ĝmp�9����A%ڰ븑iY?�!�h�̕�y5nA�����w�q�iX��4Z�m{<�@�vf�ĂS��4��g��-Đ��c�#�k ��Mdw���mt6
p��!�����5��@u�:�_���JDx�k]�	�������)��>T��>J����:�h������m������2��e�>�0<1n){�d�ml:�.h���C2�b��́�p=�۠C�tٜ��T��0�%��L)�	��-b�u]���jia�|�KM����n��ɢ���&{6��,D��Ab�E��b��R���B<���I�,Nԅe
��{�|UW�D�<DDz�;/�.�k���fL�k��%��Iߌb/�T�)KC7�[:�0o��0) ��
�H��n�N�Ga'�F�1�{�G@�Q���cњ'P�Ki�E��b�Ƴ���P܊�W�(�vC���a�7(�>6��!{.����I��8��K���6\8|&4�r� e}�(X���g��&�Ht���:�]F����2P�[O��0�������˱�g�@�3pP_��{aN3��q��s=�d�F��u��*�rQ�� ���I���1���˥flx�c��I;lF�������ZH	�f�+1������ó����"�"�,�F���D.Ѓ#٫��(m4�=8t�c\
�yŧ�i�+,t�Ф-[�N~�&�+���ҕ�t�{4>_It�~F��71%��1B�֔/0��@J�N��f��M��|Y�'l?n�Ze��*�L�\����=Aׄ,Wa�k��D"SY�h4v[��pl��Uq���䷬��M���^M�I�jy�o��� T:;H�x�6�<}���q~.]z���L�!f7�e��{�4�uH�W�#CS�Z�_P4����d���W� r/�փ{͎Ke%3%�h0�Z٤��D𐰧���: �W���oپ�.LB��Ý�a�T�|+�g���;ϳ���f�O7Ռ��x�c�'����	>�8_�-K��W��`*4y��H����*������>����G��*4ܦ�,�5M�j�a#pR�}�BN�Kw~"�Җ<����?s�Yi���a�A����o��JFt��s�n@$lB�7��97�eYћ#��B����s7X�U'�S���Ɂ�n�	�Ҳ]Zl*L&��ө���ͼf,�72��;�	j��,������0�Px?z�!�c6���h��6G-��M	<�1��<rt�Z�B���`��vn�k͠5)��<��S��7'��n��L��w٩&,�7��������3Q�j�����Lu���3������p�}T	�)��H|zC>oIX�����t�v�^d�@��q��P�Z����l��34� �n+�')a�6G�'�ޗ�;#!�?��F��*Tc�<XW�r-+�+^/���S�K���͝f�HJY.�*\��1�γːV��*���^86��0�ε�+I�B�#���oɂ����t�I�b��~,��ek������I�� _,8���j\o���`yů�D%\�E��[�>��x��(�腘#�f���g*z��H�Tb�$c�~�7���V�M�ۚɈ���
^�!4����6`��A�B�s%�Ţ�글x�s������3D�N
��HĭٓL��x�q�v��t7���N�ؒ�_�H}�a{�02`gd�g���ݼ���;g�A�"X�z�A$"h��t�(�` Y��r=1 ��a!J��Uj�4i����k��|�����p���F ��%���`ʲWVh]N�7����!*�y-(TN�'�	��@ �*��9��.���3�ʦ��5-�?KmT��i�2M-�z�}��(a�p�ic�~�v��w�DR����Y^��g����Y�%�Ur�QJ���*d`x�g��Ƕ=�ĕ�m2����qe��ȓ�w���;?$:B˂ ����F�R܌��u��abaz�})�eY[/J���Y@=�<O�?�H��i�j�w�$��sED>Iw����t�ӏ��fT�2�37Z�t2���k����K l}=1��\�!�r��g���t��^y`_`�Sތ�z.qD��Mk)^'����a��}ސa� k*��IK�pP���E�K�ݻw�	�Mj�Ș�ͺ����H�k�k��;؞��q�A;�8��[���e	��r���-��X�t>>��sK�����Ƶ#��A�14<4�;���Ȁr�N�J�e�oV������%>0�S���$:BQw_��j�>Y��
��bs4)���"5ca���� 䁯�"/j�<�I�[W�8�o9�!�L�߻�<X��juc�a@��󌤱Ay�8Z��{�<� 4��D�v�n<�Z�B��atC]ˣY��?%	�8���g ���<��".w��!������y7Mfr��Ѷ#9�A�q�P)\�� /ul\�*'�@�U�g.���3xs��brϹ��v/^.
�|�M :����W�tU��O����~\q���w�����P��F[}��������cp���{��T!x��a�/Y��~�>��/�n��x%8�a�-�Jk����wT�����̗"~��=����O�#�g|/�n�Ԧ�%Z�(l�<^+Gqǅ?r�߁��K>A}�.R5���/SE��A,�|@���94'�_��4D�_؋D��Ϟm������)��c�"�+$�!� �l��w�ڧ��ȗ@ S-oF�p�۴�k�X*�h��\��PjڣQ*��MsX�F�t����S���2�Ы/gC�є��]|�Z;�ՠ ��M�A�L�̺�"2���C��_��ƾt����~�s��h��!��vu���Ұ15H��3v���!y%����m1.9o��|�_��a�AK-���|a<Nr2�R<���Y�,�h�*�7��0���sjv�g����  �)+�H
��� �������+WyT��M�*2<���ɞ�}➩9Oѹ�#�=��b
+��jFu�hE�׿)`��e��u���Т�WU�WTq���'�����"?�K�4�\<uL�L�^[BH�QZ�3���ꂠʑ�z����>���sg�b����JWd۠�lt5�l���8����>� z&�B����806��OZB��HLN�!��� O�'�G�7�"_)qϵO�������?�A�����#��n?y|�t���?E��9m
D?
���mxm��9��y �V�C����V�%]U�_�Ym|6)UM��+E��_͹,��e����.����8/�[%�Q��[��Awfk��n��� �<�����V���� 	�*����	���w_r�#�6۹$�w���W���ȸ���G��/��o��~��^�_V�_)���ta���!�"zc��siW�RM�^���o��dw�2P��&Q\tۗ�3E;찆|��zgz�	�����\��CL�ڞ��c�������1Uj�8�X4ãح��y�j',j^]p/�Ĉy񼣳So�1e�J��Ո��`v ���3_�Q�X��q���g3n�� �U�hj�� �4B_#�����(z� D�?��w:|>g�G%}P����jc|Y3e�gU,���z4m>�V��z��X��y�KH���.�.q뗊�rCxs�]	ɛ'��,ZЩ�����ʜeC�Хz;/�v��lU{f�M�(�h��A� >'�}�<�xv�Ǜ��5����u�Ү�ag��b��I�Lɶ�Ζ���N�db�3Ԋ-�@#L-Ln9��ݬ6+����m���'잤%,�p�J:�L8X�f�<W\���o�d����@e*�� �P�5�,��Z��y (��E�C�8���l)k��F6����Wh��7�	�ru���a2(��)eI���t�j5i$���.�] �y�l��c�{�6�rXd"�f����;A��d��q���_����Ri�N���>ԩj|W(� {9�<��Ǆ����&k�}�Sj��0@����� �?���֔�����H�~%br���c˵9JPg���t����	1˦a�����i�U�-D��,�J���T��GH)΋�(���:�rL��� V޺��J�w��~
��#��H��~�|�9)y�� %��,@@s ��a��v)��0\��_WZ��O�
�.���?���Z6y��gܫ��(K���E��GPs��B���(�pk����=�40�f����b�F �i�d�ǰD�X	�V_�,��c������e��ý9�ިw�k<?(:��0��Xְ�+��r�d�b���B.H�
]Ae�Z�x��r�a쪽m���R������cn��8 ߬�i��UJv��p�eT7�X����ߐN ����b�dJ��|D��w��ѧ{Q��E���;����]�ߓ��NSK[�.���Oz�lP���褐	�� sLFιR"����}�@��B�i��4x<ɏ��1-�TCC�����ɔ��"���X'L���2�K�h��Dj#�ð�q.s�9�<o����_�J\[�fY�����ς���x�^P+���ߟ��"�}L��/Ԃ�VI}CK��毯��`)�U̖��Ј����v9��/��FhKcpa0�le�A���Uk,v��b*~�]��*g�r�$~����~�K��Ƚ�O~�>��S%ņx�bd��t	��A�K���BXez��{[s5�,�L��1����+�&A��j0�qGH*��Bݘ؉T�U���K/��~"cp�﨏x7�X�m��n��IO��m%��&�u�e�{��	���x�v|����~ʱ<��q��[. /,m^�[��T����x)�O���p.=OH��Ǫ�R�����!���Oƕ��B�Y� �!"��l���ߘ�k�c@"'����}c&ši!��W�$��3�K�aQF���6�P~�D��'Yt��B��1ض����M����$����L>Rzd�a��[̮���!�� c��[7��5���*�ሿK�VXs��?�e��}�;���Tc��i�2�����<E�ʁ�:����v���'<�Jz�3R���	���L�yZ�Fi8��v����!6~�5�I"f��$����С��'�g0�M���-(ź��5��1B�&,�Qyf5Q�������V����y;��i?��G.F�����J|K��NQJ�|�N;�1|�U�l)f����u2�s]MV{������4�*��WA�І^��
�" SH�o�A��N����P�^E����a|�زη��c��v�@c{�����G���9�0�u���u,��%�:�0	���␈SC��-�����[�2tx�1���J�)r|�FvD��q`��S_�Vh0����<X��Y�W��m*'��7��7h�/��M�Goa�߬a]`7�j�ݺ@�6 Tc���i����n>q�i-�#W�=�p%ğp��oc9 _/�B����x6 ?v=K������ьc��Y��I�a~92��6�lu�Ҝ˥��*C�ߍ�֘�Z!��*��ǃ)QD|��keh�" �f�SЙ� sg�j�N&՚}�d�Q!��S��j/6�����Yb9Ml��NI���� �Y�}���w�;� /��!Ʉ��?��в����Ct�s����b��{� bH�xJ��ޭ=s@
o�լA���us͙��cX��M���E���3��B���f��웢JIn�_��1N������Y���y�)55���}�L��M��g+R��I%�E,(޲��Q�j�x���Q*Bg>�=Lq�w���zY����[d�Z��XA-��3]s���� E`���@p��D�^�C��ۋXZ��"���/}݉AD�z2���V���8�s�J��9�eF�����@�����+���=�z׸q)�;,�n<�����i�EX\�@�1ۅ���$�����#w�J*}�FjS"�'�9u"�(��c�R�cxp��G�w�(r�l/ h�.�@J�O�_�dc%}��4��]-Z:.����GЈ������tRY��L�(��������0�aRc��x���r��y%��=j|��8D�%aQ:5Ñ���l�������V	vK��N�!l9:����.�n-�U�B�0�b%u��{3]8p��4,
�2��W�5���u�1' �Ax�˔D��h����"}���2`*:9o�����Y��qT�]��O��Kd�S�7i���\�Cg�$x�u��Ke�v~��Һr���αlhh����פm�:�|/�d�RĬ��
�5%-�%;g÷�N�#6��D��C����Kի��ᇡ�ܺ���g�KL��93`l���mmc�;��0��ԅ�O����Ϻ���p��\����*��RO-�à�Av�E �t�l<�Y"�y�δoӲ�ڣ����m����ħ���	DT=b���4]��ҭĴ���{�1B:M���z>o�%�C^GZ��]������O��w`�>DaŪ�w�uSLX�&�!T�� �3�_�v /K�@����B0����8��ZۓP�;Ƙ5S���]_��3\��%��N�V+�c=��^T{t#��+�ޟ��D/߇��Z����h����|�"N���� +K,�Mh�@#A�KX��4S�Y��B�X��p����C3S������|�n�xt�A2�m���H����*zך��	w'&^bE�1��ƶ��E߅x�V�R��9�P[���楼=ѧ��!�c�?]��x�S�<I&
ݙL��
�������l�d�GC�o�6*��s))�FK�HR��,�3+����0�Gg�2(���g����.���^���1��s1���S��$Y-�_����v0N(��+ڤYIo��<���ͩ�B�,_�6j��
���p�n~����k�8o;�m��<f������G��1��8��&�u4HA��;�D}���dh����H���\��#gj@�l�qes�p�L2�q��J4FOA[s/ի�z}�T��q�A?���K�Y7=�h�`���tc]?v��]���WA��w`��#2��Vv��9�{���Rէ���؉o{�q�����}s�ڛ�T��G1��{4x�XF�-0'E8����z�c�O��\�����/�8�u��M���h�e�OBȴ�Dҙ��y1Qj���I�5�]�9E(��%]�I�d�/��RO̥�Y�n������k�ʵ!�L+m]��Oˇ�_t���7]Ry^���;ٵgM��X�;��9椕Q4�	:�?'n)Q=����6�h����cQe���q����zl�ŉG��'�*0l��;3���*-�"j���~�T��呋60g��
r�.�j̏&2����a�4th觇��v7}�[�5��oa6�^��mW
�qA�� o��jB����w\ߚ1�b�u�u�5��+���ݕ��Yz!�\�m&�Vfl&�q��6/���>�� ����sԿ0;ͻ�p	��� ��W3�j-�Q�ef]�#� ��϶|��Rp�!��)�ǘ�)�<X�9����q(6a�Z�?zg���?���/�^��C1��h��xp�f��a��7�Aбb�A�����k��j9��
����fơ~��SY*�FR��">����د٬<�1�Xk�{H>�	ӛ��!�&�2_�2���8��w)��� (���3x���y����yn4��!Q*�s����|o̰xP�F�i��ͯ�#c����Iκ
@S�.-q[�_ p'	��<Y$&�Q�oԠ�O9�@ӆ;&���&hp"���M�&�:{�j�wLPD�2�`���)�C瘎b��Ɲ�%sV�#��v�3����)��z��x�l��P*�f�@�E� ����F��V��R�6�jع�(1�0
�s��!���9�$h�pg�"K�H�W������|���TCw�1�C"k��8���0�`]��2�-E_�Ў�a�:3�Ԣ���ܨ�R$�!�QN�2~T���*ۨ���N�`}pg�KpUgӘ��f�?��@��xx ���Xm(��<P����Wt���@�O�� ����=�,��1�&�� U��?�z^&��4,�n�z79jQ�~�x�,x��w��I��*�a|�D�+��A���\�����-/����R9��'h��+Nj�¥\G�������^VB��EC����o���@�.Ft(iA6n��y��l����*�~����9޾&P���'���ZԽ34���� ��F��q�$zq�j�b�KJ�����Q~�@�����(�|ә��L��2P}�S�KmH���m���6em*ENR�3Ikt@d&5��a5�-��P��kQ��QuF))&���|�nG2�1��1���f*,��
�M51'��"<h�ؕw+�����{g��|`Ü��;?:ֺj0�_�h�r,��$X:;%nt�v���b-_��(a����p� ݍ�mP������ ��ŉ�ԕ��aK�JX�/���{������Zm�"�9d��1z7"���e�h����\�֨~�5H�gO߹B�?�~�0��C+�#�����;QI^j����[�N�߱��������Q ȷP��1l����4h;���b����ؔLX���Z`Q4Fʶ��^�ܸ�Y�1��+�EO�,&{����W�Io++���Ԇ�"b�@�[qN&�b]�<V֎c*.=Mq�D��)���hS��fC��V��>�����=�U8I�Ggj��oG���`%0gH+�:�]H��K	�'����;�gb&{[Q^�H��y�N��zz�p��xY��%�g�vO���o.����r������o���H]P��qf�xJ%����~u<~�L��Nәh_��o�k�-Ů<����85��Nv\v�~�C���L��K_�R~Y̧��!	+eT �tH��X��d�!D1�X�r�P�V�^��8���o��o�/���j��[�6���i1�dwc�:�E� ��Ü���w%^:��
���f�pR���֜aias���=ғ���z\�{o"٭k%5����~�N�x�\ 9����������J�z�s$�]�ҩP��EKeN��.��]րP���?��H�3;����$~z'���;~�É�H!��f���q�ߙ���}�;�ހ܆�Zm�_�/3F������=K`����b��=e�*������ܩg���MbS��~#��H����(�N�9��`R��1����	��g�漈9O�����i�ix}5��9�u+UǘZ�������WD��g��	9������%v��2��n}���=��t��f��a6] �Ӡ{��*T�,
������մ�D3�=,bT����
IL��V(���!�+u&̈́��0d�Ұ�x�����b�_�?�X徠�%�}���m��^i�R�y�����/�`�ʱa��7�/��G�a�
F,E����!�\�yg��K����F4z��f�����M�|00"�>�ӟ�.�@`յ�=R��<��UCs����q�����+��:<U���6��X�_��O��KwMВji��و�n�t@̧{�.����{4<,-����vG+�H{�����m�g����۞�(�	'
D~�T���@|`�x������A��+�Zg	�3.��D�e=�V��NH�{ׅ��v�3��_�!����mՈ�-2"k%v�(���@~�pa�����^���hT�Y�л�nV���yS��j����i�3��X�<܅5��B5|=��z!�o9fd~�f(�����j�}]M-��a�a��~�"'��o���v��D#u��:!V@F��;{)�wSbe^�/]f8�%���]���Gx�0%� ��q���i�Ԏ"c��~``�- .��QC�Ek�g�9,�J-�'u k�X���R͟�Z�-=i�3��^�ܼ]�f�$ٖ���3�06"x>�������������=��ܯ��HTP%����	��.���?���4��h\HBkA��sS�a���F��S7tt�i+�^.>9�ŋ`g�ē�����G�j��?�!�:���M򞳴M����<c��o��&�c�}������B��D��Δ�h/��K� ���{KQ	������mr��/�9(N՜�����Ȥe�pkX�6�l�ڻ�#��5���m(�C��t�f�װ	i,����}�,��-M���a%K�7+��K����W�Q�@�0�����{���T ����y�{��t�����s�{g_)�C������@���9���tJSԋr��K$	SRߒ#*?�!5L~#S0B�xĩ��~w{��Ps���i�(�B��p�f���*�S.x7� ��iי��@CI�T�	쳧��;�4�Ϙ�ҋX���lؗ�/��IEN:���:K�:�נ�\QJTh:��h�d�)z�%��n��&K�c͆���mJ��/%�ta�6|tq�hLz���D�j6�oJ����Zo��%�%۰D�����=��0q�IfJ}��zD�8���^g���P��
lVآ����:����9v����M�	 K,�g"��4ٜY:��|��l����v:bE�Mu�;u��IZp���&Aԡ��`��������"���1d\+�sF��*!5n8M4g)x��Q�ށZ�<� ���;:;y}lk�I5`�D=�I{z_���u1��2�=�!\cf[�\�����Y%~7�Ԙ�N�d��1'�X��_k���i�`2�Z��e*�]�����|S�q����
K\���!U�S��5Z=����R�"a��)%g F�w��C� ���(���*N�ΰZ���&����F��;w�)�<���;�����	�ڽ,�<z�,آb
̽;�ji�OI�Ѳ��7J����P�*]��<�Ж�@Y��=�Z��o����m2�~0�3*�Sgz����w��k3T��Q�ҳ��̮p�u�I( 2�8��Z�*7�I�&�y��8��䬓���)j7�l9j2�����a՜��8���E����_�l��������2�_��5Hz�S�\}���}�2w�,��{��������r'4��|���G,g���3θ�Z���y�;�/8-�� \#HĐ1�pt�C~��������E�勽�%ߖ�VG�'*
T��k���&+-\}Și|�x��{xX���J,�����.(&���	����k+J��H���6�#�Ё����N���45e���+s_6�$UF�:5�9d�	,���NI�1�����7x�D��ϯ{���I�ʺ�-�?B����}����N*s-c���@Ȋ�}v�a:���I�Y'F���������j%óH����{3T�E���Vs��z�^�lt��dn�����4�n�G �]�g�<n	�0��ҟ)�ߡ9�u��2¿�^���+�����	6p��j��\���]׈�K�����J�f{�8�������Jw��V�s���T�y��
����U��uo�m,������ҙ����z�0��n��./~�ʬkpa=ԠY�u-UMQ�S��Z��)���^d�ս�Yz�W�����x������"���c�
��񚈐��0���X�^��o@�+���^�^�GZ�+!0��\�o��� ][YzuP���ʒ���fһ�_n���Fh�Z8H�<�1vmx0EL��7ȉ��:1v}��ռ��wC��>l�~���^hN�u�z{kˑ|�I�I�Y)�%cԙ�Ud` �@��b=V=��ٲ�j��z�s�(�&sԪ=�{����JMļ�9�#="���'����_����*���Y�VFBY�6a���/�?\��/��������J?��ct�=��L�,���j�hܠZ.*F�=���{������.r���¶&m#v��=��ς��N������r٩�b;�%���/u�x��$���k��3ʜ���@��_n��!�A��!U8\�I7}�)��Jئ\3>��<��[fG�?,�`�J�X��x��0������w�E��/!�A9��W��鰔�AX�H�N�/��R���뾌;-%�Y��1�!��pu�	�P�}^^�ӏ@v?{�}7D�m���6��;{JW.�na.�]}�)(���=��ދ;��cT��|���Ȕ("���Hq)�#��[�k�(h�6�h�i韔��R{A��n�f�L�c|�ӷ?��p�-d6k:��JMoI��i��\����?X��v_H;�����\
����W|$<��1���17:w���wD+��S�D��<�hV�V����RB>��n�j��^�� �%�v�R7҃T�E�)���43;��q���l+��`��ӎ����n�~����/!��c������G�eEڂ�wU�޳�V/�q5b�i\I��!\Jy�@�S�&:eZ�U��-64Yl���a�`;ާO��h]��3CVi���5��q.�X��(,L���o��#�{t�z�fq�J���1M�W��z����Oz�5�^*�f<-������5���a��{{�R��5���� &(�!U>����tay�{�'�n�۟� �ieW9��1��+?z	��^��r�k�w���wO�U�>\����/�y8>0!�6����U�A�J��#֩��@(���7n��  �b�$���v �I���o
ws�)G)Rh�.5�
�Ȑ�� |%��KD+�:�U���������]�HN���-��K�~��`jm��P]�����)MU~T��h��7?,�ɈQA~mL�H���]��z~KBX ��kD���F�Š^�Q��p��C�~��P����Cp����Iz} �ɠ�#W�:�2ȷv+*90��4i�[x||��O�7�O'�*ēn����R�� '�]��15�@�"r�#U��),ӘTI����w]������t�!�n�sڔͰ
�y]�%��e4@���{� m���5�M̆!w�=JB�@��O@֜DG �Z��RZ��~�=���W�fg̝] }i�ϗ��җ�|� �jT��|1��7�b�,�I�*�-��n�~5��\�n�����,ѬP���>�? �w�-�� ��T�)����ZF���x�TU
�D�$$J�
����h+����HBB�i���]e�B�m_��1Ś��A�[�[-��k�Bk��fB��Iڷ���"/>nCHa�ު?0Gd"�m�A��[G���Kf�C���lLD�H�/��~.���B�%!0#�ˏ�^����q�CY��7z�-L���`�Y?�(4��k�����:���* n�j6��!��A���f)�0�\_���!��~=�g�e ,9�"��j�����[�t��KH?��ر��?c��1O4��W-��oF�H��Y��%%�=u)s@[�}C���fX�j���2���� cl�_TP$m������n6�ߵ#������R(Ȯ�ȍ�I�	��xI���<�bK:�CM�{��N\�����n��%R�]��s�#������i�Tb��e����[O�VtBj=���{��f50���;�i'a��?(ԧ>���,��,C��A�����=���Gl��n�t1�@���;mCy���G�\R;�D�$�\�3*�����-�zr��p���9M����.M��{n;NC¼�)�
4��C���fĕ��� &�K�|EW�e��~�D(��zI`A�5cb��w�H��D��CB5P�(U� "��q<���s������n����h��=J����ɓ~ �ؐ��{5�(Z�~���(��[Q���lkT�mSJ?Gz�Rt�o�j�Ǡ�D� }���s�i��ӸFHD�����'"{�q�7ط�h!��%���N�ˉWW��nP@bՀ
%.CՅ�������/;QJj����#V觶P��a�G3�sY�����&��\u�M���d�P��>�M+�
�n-�4��D'��}��(��	(9�iD�2�K4�7S�\�}�i�+ڃeH_�E�rp'�X:�p|
���cvřd3�f$\�6y6�&aƤFӿ%�~�PnJ���������9�i�j��⨑ŕt�C�ݿt���*]�>����s,����J�?_@� �ch\I�*5_�`���4%u�;z���u⿺@7�������E��ۓ�IUG���­#�Fn��8S)�����P�w�H�ˇ����bg�:Tl�c�u �8�/�}��]����)�U|q�t	U'���z>_Tv�qJԗ�&�5����`�e�d��H���	>*��|�Pb3عF�Q���a[K�3���A5�wlJ8�^�{.�l��sK���z�R�i��tsuY�3 ,���Y�[��\<[�*�j���>Z]�{�����I�/V��%]>��jqS*>/�@���/�)9Ԣ�0�2Ky��N�)����h��s�eNZ��+�W)JyL�E2�]._f�[��rm]�p.}��Fd�ɦ) ��H�d؉������և���2��7D)� �k_�E+��&3�ɳ�<[��RoH��<�	�W���$��� [�B�Z��R��d�w�2NA�h�������T��̗�Z���I�}�P=q�4b��4�u��>-X�{�SJ�i�ww���fhS=	q.5fVz�J��
2�֢:���]ټ��n�1kx�uq.6�a���ZBDs�Gâ121����s<��R��3_��`���i�Of�AC�.��p��꓃t��	;ϼ���:������{���̮�}]��� �����On~n���A����e$]I�Y������F�-�O�� �2����F62b��9Ѭ�ܝ!�� ���r���i�n�d��c�XA�<��A��w�&�L>��T��򜃙�"���۲�0 ��F��[����(2�i�BC�Os�8w���^����Ϩ��G�P���c9�A�"n�������� �~�ٞ�b�i�:�L�tlT��r�.�@�?�э3e�K���u�0qv�?��ƍ�H�Y�caM�M���������Z�bd%�k5 ��}ʑ���Q�yw�°i"O���pP�׼-uO�n��ܚ���#��tLU��
	 C�$�Q�ބΤ��s(�2?�Hz�������|ž�${�U��t�����'����]Zm��`P�i��:�N���R9��Z�j�#�R�j�9���=�Aׯh� ��	3�����q!�)j1���K�)�� @(�E�����
D�X#&�BqC=�)�|2�p0��qR��v�R���_���<����+�C^ăq�֫��������JWt�Ew�`�dJ�D��e.! `�R���Q\`���9|�_�{�C3�1P�<Q�II��';~:]��.�Q��1��p��@M5� �y�v�m�� iH��w��j�����j`��9�DfS��yfW�=7����]W��=�?�����<�ס�B.�ጃ}M��D��<� ��D�`��7Cz~��Y���_��Uck��bۧ��'R�Oq��iD��uO>��՛����7��N�'(Z�F���?�8�3���:��I�n�����[���'�B���m岗�4�U��]��)��H_&��S4�%��,8�5��}�&v�/� ��m3h���?ݠDյ�\��z�x�D�}�Ifaf����ǂ�Z<�z����A����r��ndN��R6x|y=M�9�ɍ��c�nX��kJ�ZF.{�A��2A��1�TB]M)js�]����A�Y@�'U�7"��5)G�[�X���<5�g��[Ŝc�_9\Xۯ��\��ť7��|k��L�	����)��@�>ɤ�\�rFs���o��FC��Ĕ$"��k��}���/�+�tPG�_�����!@�����ї�R�yF0�-�`�jwg�XGs�=�Z��0�z�)w��X3M=zh�p]6B��D�rd\v�jXuƙ��'���~r���F�Հ�C��x�|!q֙+��K��4��<�3T:�Md����Tc��T�a���r]��>� ���Ig߉J�.�ⵤ쨢`\��̾<��5)2��O�R:9�sVXS#!D2�6�V��G��@�ķ����
�F-���s0�Y▄	��0gGr�8]X����2"�9�t���O!(�ø8:��8�¤�s�9\9��Ktu�&k�2�q���P������܍�Brr�����l4�����Jb{��B��!?���%-�O��@�]������,��sJ�*�H�=QEZb�%�e�ƨ�-��T�_��N��\�@���r>��<��*�(o�4�Pv�[�L�6V����#[Cj�gM�?��N�d���h��)8���lE��[ɫ�Ik���s�q�O�<T���P��?������+��b��y��.X�]�����y`�������"g��oO���k'W�ԄB�ɹ�yz%�m���NH nz:y�$S�NGl,n�T[$"g�C(���sL-����uuR�Q�_@ZB=?�W�p��p�A �j2P��|q绱��t����i����LD�a�Y�P� U7��7�kP��+}=gRI]���R���Ҽ���mv��&j��j��Y���ڕf��M@(0%�m�yT=�`�V�F�HG
�g�4ʚޓW���X��Y��c��%��R��"�^�o��#���c�5F`>�/�0;x�K�'$#v�e��0QH���)6�HG�l�	�QS;�>Gmʷ%{��=��}J�������3�߃Q��D���7q���1�	5��~<�\˩��V��O�C�Aw�J���f�Qϼ�&�I�+;���m�P)�)���jl�|�pe.������]T�X���d����yՏ�=�����\��I�!JΗ���2K��㲭���1S��x҈�E3@C�+��}��"z���C�fLG0��~�'�Cv����x�՛<&�&�
WW���FRx������=o���.�bqm�,��`�3�=(�Ft��nˤ
{�U=f/�O����ǔ���{k�r;Z�����aO?��� 8�p��&�
� ���k�jb`wb���DЭ	џ��k+��A|�/Y���1�;��@w�qraꀯ8����"FQ��lUq�DHO���Y�Gpz��Q�����ÒpӾ�� A��+~�(��F�j-�J����E��MD	�85���LReu�dU9W�~#����5v �!�6�(^�H���WI��(Ռ_�U>�M?�3Qy�� ��ʞ� ����α����g޶���徱��3�oI���Uc�g����a�.x���rd�r��n��}����8��z�5:|^�t�?�*��;�}k'#�=a/rv�	���[���+�?��C���^F��,�\�륶�O�ž���T~d�#�8�0��ҤU���aW|ʅ�������_|��@��f`���\C6Kz�{�'ͶQ����u�����v��2��s�-��d�j�]��ؚ����@l�B�|+�rp�"$��{�ĩp\�@(�v`m�����Z�2Z�s�ʆO ��|g���q���"s�(O��I��������ø-i�KŚ�pӗ�p����v����e�;�Ji �8�u"D(PV:M�^)�������e��F��2Y��t��{�d�����S���o�h���]�7A�!����tQҝ�D�RA�7�ڑRu��_��ŷ+�xQ��#G�ǥ������O;��D�}��ʾȃ�[�Q��:HgNd -{:��˺�ң�?��r/�^�]���D0�<H�N��?|&w��V�K�C�m�j���o�;\戃wMĽ������I��!�0���
��Fv��Y���������Ƽe�PF1t3/H�0�a�E;:�?0I��՘�\��Y�ue��#U_j�w��gS!��_	ɺ�m�X�>����ҹ3����33�����?T2�ehCg.1��aE��ug�h� PH���~@o	�F�/�O{\5� �h"�����8�>�jĺ��<C����_�D���>A
�e#?��U�N�c��]͠��[	��,ٱ�9��*Y�XaxubneT�k�5�y�7��"w�}Znao-y�Bݎ���`��/�ºtʼ�Wd!�ſ3����:ѵ�8$p{P�x�0:$Q����� D�THy�ĭЍ7j�K�ƀgBy�ggsW���>($v6.�\�}�6���5J�O����U�O1w��@._�!P�q-�:C����/����<�$X�"�TOW	07@m�>�&�ۼ.>*,E��S+�$���u���:Zx�#��'U"W@U��@�|����#��g�`.Ґ����:�|+�� ���ڇ�a��c�FF���B��v������i��S��̰�t3�NP6�t���[�W�����!�&rP�����(r�-���o	E�/�.�i<��Ϫ�BX����l���8��֫��|f��*aX"�y��_�u���	|9���P����蟼��g�g8ٹ���T_��y`+C�#�������f�!n�/�*O !���S�K7M-G�M�̾0����Ls���$@��VV�V:��>�>m��;�yV�� ��!�.,��(��/�%{F��_94�>|��R���ڜqn�aRc{JȦ��e���!�H���{�k��k~s0FZy�x�3x5"<�7}HY�g:c�aѣS��O�i��4�D��RHTAlc��9�ۓ�u��C�^/2%k2�ۜ�zX��)�w	5�BR�:9�W�<���a��ui��v���;��|�9 6~�D3:l�\�e������pI-�pr����WY)U�b��{�Ql�2�Ue\G|:r�[�G����;�=�"�7~IG�i[��,��˚�}Y�`��v��K�b�8���xr�����#W��&�"�*B���֊�]P��*9�[�ڼ.��AdM��==�1�i���|�-�ٳ��o�5�1�����!�7�=qkj�h^�]$Z�/w�m*�ŢӺ�=�j'@��$�4r�^|@c�oy�(��zT�[�邿�Md�]۰b�*�;���i匶�{��@A�_U��v4$�lP�a�\<�V<�L��-N�:m�3p�kS�06b��;�)%#W����b*�  ��b�á��l���欗d�"�5�>o�U�W3[���ǿ�n�s*I(����Yn"2)l��Y����{�-�Ԭ�c�}���17%w��F��8����2��7H;�n��N�j-L`��x���9�ܨ�/b���hӛ�D8a8�@��L�?J�pa<��Tڪ���⊨�rFTIF��"rib /��������z(�띳�����iY��u�������ůA�@�㸽�}'��l�Y�H;�Ħ[���(@�̉��y�X@�u/AHr�ᒓ�"�߅��i(=(�E8�|;��f���{>���_�.?�AO���l�c$؂�c7���DXtԳdv�.
�~s��<R�b�J4�����������%��׺y�i1��.Trt�z�a��.�(�ʺuF���
.�Y�7|K����o��r)H�A�� Tsk��1,m#�O��? X#�8��} ��:�������p4
%zK��g��ȅ_N��`���l&U�s�w��3)��(�2(Z[�y!9�*�|�K�����a"��Ӄ��l�>�v\�Ojk�y{�z���G�,머qS��G%sBx�������0"X��9�n��1�j#��k�z�}�1��T��t�����G@�fx� �����	\�}؟S 0��G$��)�8:��C�+��\h��q���+b��+l��� �Q9w��Ҷq1�m�g�Y�i���� I�����8�:��O�����=�����On�XNt臯������W�.��2>2�����<L�Ϯѣ��AV��Va��t��/$;���T"c��/�˴�l-�j ���6/-B'���jUuck +�!JganR��x
F*@W�AD���:g��@�t�2�B|�{Uy����'��<x8Y���.����F��TȦ�It�� g���Y���'�?*���a� �8�1�x����)In�/T�i-����R�0L�N�#���W�kl���('%�o^��SI�X��H=�2�~뉳�~4��ޞ(a7Cp��B�ғ�_d�r;֜2�v,\�S���Ҩ�5P�ݑ��:��j,\5����+
3,�`�}�,)��KS��Bݟ�%Q4��R�Ls�?'�C�kĔ��qeY9�6r��U�!���:Œ��MTn2�\ ����mO�Y�2�CF��5�',�T%#o`�  �c5r�����SL� ����d�o����$xN��ǖ�Hg��zտ~Q���aU�����=�>�~�KD��C��Lˈ�K�'������z(.�#8)آ�� j��:zzObtLXҏ�t3R�|���	ڌ���+�W��_kն-x�%q���xR&/�;���X�=3n7�"G�c��X�WY������\�gN�F�,�0}ѳpe}:��Pq[/�Q�V�'ީ��P'e�!M���O�dk�e>VO|���3z��h�ɤu�M����Z�gN�ge4�G%S��|�P����)�!���5�͛�Q�����
.Uu3�7�7�6~dkӆJ��p�b����G+9�:�h�6e{T�����~�]� !G3v��v����oĳ>�`��wZw��6m���,V�P��r���^[b/o��_0Gh����?œ�}��m���������+͉�t�V���"��.M
]�&p���H�4^����	����@?5-�[�/{|�Ҭ.�+��/�Ff�2��ٙBJh�\4Ḋ=`�=G)j#հFU��)~yf0E=;�ZW2K(-
i���c�P�����O5��{óc�a������Ac^�ϐ��'�PY�0I�T[ ��#[^�M��_8T��Y�r��[����?t)�����m��4ǫ7��|Əs�p�7(��;jD�Y�j��q�\$�A>�t�����3JJ@>7�f7P���`�7I]�@�Wd6\�����_b�����Bjį�yN9v�+J@'�<��ñ��d _9�0!�l�������� �1{QLW�ι��x�^H�K�	\D�1@�_������<I�^%_n=��h��VGާXq��D�!����'!�U����R�X (҃ob���X�=���t��"1*c9y�A)ך�t�;��2R8*��v�y��(�ʾa����B�7�ӂ`��u}t�황܉�3J�V�<���$�����z��gV��'�@�8���"�v���J�uozZ�\���|/c�#���ʏyۚ�|��yOAk��7���X�!o��q� �C˶���.&��<;]�O�]x��pҦ"EqS�F�:X,)ń.k�K�d����8���i;2`*�:�q"��3��G� `��y��k7���Vմ����d�Q�gx��M^�E閊Yh|� �J�f�;�ɧ�G��l�!�rg�.�B��BL	b0ǻ߶Դ]/�� ?4ؖF��:�*�Z�`4ӣD�
Ie��8�̶LK���o�����22�$)`,��c�2���;�w����j�U���ѡCfVQ�G	Xc�#lq���|.���t_"� �D�iW�H,��*�X)h;{� 5{b<��[~���m^ �;����[�$wR�l�c�rc+��޳��nyG��gQ��_-��"H���<},?�q9�A���}Z��gn��6��[�-J��-�U���v%�sL.���*�G}'x�7`�K:�ݏ I����4;'<�xv ���6u^8���]�>��,y��^��A󑈗y���q�@-Rb���t���5�����Ye�ݜ�9�V���$�1�*�\�"��E�4U�t���83{���V�K��Z���O���^>e��밎��d�A:��{�2N8���������}��±qQWpjӲ0��0��s(-�����v��oɶ��X�h�$��Uo%Tf�{�����f�B}��H��c����}�w�).����>�m��v�&�V�{?Σ��5[�=F��ޣP�q�1��+�A	�ъ��BB	��Xw���Wa���x�i��qHU^͜�������Y[	�UҐM�z6�ˬ �%ઠ��~m]�c��s��`�k��5���|����W�y"���_�K-�%4@n��%y��]�졉���>	11���o~=�֮���3V�2��*�4F1�Y�M>ͮVg���<���t�P�ra�?}�<'y���)�)����8_�I��I�Vqh�,�Ai��<Ϙj7I�/����W_�gGz}��Kg�~I�Š�~
��T���������߼�(	mt���ڛ���Ԙ$�����'�o(�]�㍯�}�­�,��dT%����s���"�����ܡP�*X�h�'=����F 47:y6�b�w��zT��ǥ�8����l��&�����7c*��2 ����$h������K�r ��? \���	i��H�r�L�X��r{����:u�����M�� !�V\�1�6'&��m;+�]j����LxiM����"�^���Y��usؕ͝�;k�tG�긁� D��I�w΢r�	�4�}�f��4sue�	N7�����VG'W@�c�9�%���g��P.|}�}�K�n�\4�����|��{!e�Ŝ���/i�����b���z�cv4>�є�ɐ��B)Ӗ�	�����	�[��S�%�'./1S�Qb�-�k�H�/ʲ�#I����ҘD����_���'=���XLȪ�ݷ��&��ar�\�;$��E��e��l@�m����V��<b������Mu=z�vJ���o�Q��pqn��S���������1��ȶj7@���7��V�o�(L�T�%��>�jvjmN:~4��?�8�A���F��������kBX~qض�*s���`n�tI�Qx����(G��z�w:>oW��8W(�����,!�ީ+ ~a8�p�_zZ-ĥr���Pr5xJ��8�7�`�+W1O�a1���~Kn��sA��h�=��y�"�B�ǘ�c_��gQ�Jk��������� �i7}7q[���IT�xL]���)|�!�6���U�F� 
M��s'�s�>����u'�q�y��]�}�~��',#�X�5� ���g�k�Pe)Y����GV� iӾ)T�:���B�F [��@{Ҩ�b��P����p�nH�aO9v՗��{%���i�Tr�b�kk��jKK4��Y��$����9\V�r6� ����ҕ�4��<�&#,�p���<_��a7x�ro��|=��k��1�;�D�P��	��rِ��~���G�]��<B> КY���|"Jbv��D�%g���ˊ3.I>�7����5d{*�rC��KJ�*/r��7hW6��ˌA�'.�Kr!�+��	���H�uu}'��[^��&m����{N*)���V���6��R��	�-��c���m������8\�ODE�S���ف��b;�i2<Zy�KG\�z�h�S���(��1U�@�2S%�*{���c�U�d���«��o���09�c�
�k�:�ު�\-� ��N�6<l�����V��n�{0h~����ӌ���������V����0#��b�J��D�͠�c��in򁑵���/�[5��T2�w�O����SD��]�F 	�����T4���1N����^o$4
$Ҷ��(s<��;ֺ�v�x,W����KМ�{D��˽hi������H��̱w�Z|���c(�@�ٯ�sK)����W.|u���/'�|���Y-cQ�� ���F)�M��&vO�ȸ�:�0>G��%��^'6N+��`1�9UMج��WT�)�E���-Ȑ�7yV�"��R�2۔����#��������	�h��!�.�tG���	�{2/Vmt	M�.�F�n����`9#v�p�)��9�~�7����t�m:�c*G���s|0lr5�ofi�~���C�?�10c�l�&[ uw��e�A������*��a� <�|�e������UF�����2�MA�g�P� ������>��!v)\xMf_+���;=�q�i�zɼ=�����V�g��1�+���	,R2�Kl���h�S�Mj���<�Ū̟Q����x[+�|l��?����J{�/��F�J}���\F��c'7%�엎�Q��v�_�_(>Q�������w���"�q��]�-�T�b�Q��
Yo��R�~��l��z�a9����G����W}���W��on?�lk���_t�6M�!o<����H$��\�����9$�V`�\
�]�S]:��K�{�	U���y�R���w��X-�Au�q�'MeY%���=�X����lV�]�u�!�����'��96+V;|���\Ò��م�4Ҕ���<s^�ʜ��i�>��.�J2��k������/@ ���EZ*�Pg�Q�ki,�&!<�u�NXٌDt��5��O�)m�|3��j����~o�^��C�	��PL.���۪�Y��x�6�RO J�MP�vܬ���s���۝�0��0���[V˗l������La�N�M��`T���ȴ�6�B�����v���&�%3]òơp�K�����o5�?"4f~��w�:�s���%8��?�['��D�G	Q�\�3��Y�k��X����2���!r��M*�p7}D�mo����/�1�')���_���#�I���c���	5�縹�Op#�8�􄻅|y���ef��ğ>����݀X>�l�/p��v��J�!��MI��E�����c���z�a��F���#�j21�%t�|��|����|�k�ۋ�;�	(�f)!�JI8:���!(��>B�ug>�8�%��C�eQ�@,̺��"7_�%ѐw���fr�.�'��ӍH.�G�ݚ^#vy/q=!���J��Xز܍�>o@E_T��r!x�[��k�l�
�q)'�U"=���(w��x��}�������T�E�#�)�̀/^�%�"�Z~<�-�f���Q��b_KV�6޺B1�)Nv?���nL>���;�ޯ>��\,?�'���n��"n��Njo���\�Q[V+��%�v<�=���kۗ.��_� %g��*u�e6�_����0<t *��i;�\��?��l�l[$@�����>�٢شu7��bF��l)�۽v���7�d׫z���,���6�7_d�R��֑׿ǋG�'�Ce�K롱�Y�֑(�x^E���!a��gr�;w@���}r�\���!�=���6S���\q��Np;�X���}���U���gh�\L�|� �<@icy8y���]�Ez\�*�JB��U#�wb��h2>�nf�	H�=]�U�CT�o����lE�l�6k'l�W� b���8��ә����L"��G�{��|�D���&�C�3N�ް�.�0�����
�}�g��k�	ʂ��ۃ�E������4⣣��F��ݕ�>j�/#|���A�	B�{���ғd�u�}�L�Q���׊:�����Q�HDO��4����)��vhk�RT��������+�F\U��t��8k�;�!GY�p��	}�.���GBk�b�0�Oa\�Ξ�8����Ymuצ$�I;�`��fh�X���1ߎP��yDz`؀�,�=U�?r!Ï*�cgjp���j����	�0����^JNϩ!Z�I*Su@�u�C��tXI$�CT{�j�q�E%\��m���z�B�qhF�~�+>��W5�~#�!�  ��XDe�+5
Zz����&/�{K1�><�8�U���cD�8ۼ�{Jj!�F�Dg��[7�dR��	ߚ�����@J�����&*�kso�ID`2�o���^&�3*��,�9���@:��u��� ~�V["d9� ����p-1n��=��4�@X��Yg+B3�m�9.^��|���(@�e�̂�	�D-pfr��6���Ų��3�+�D�����6Ґ����ǊlU�o�Z(\��s��Ջl�m�u��$��K$��{�v����j���64�Q�.�-�]Mx��f"n��1�[�Bš�8T�#�
���k�1$e���B���[�L
+��ޑHR!�h�1�Ѝ>��̛��yЯrj� j*ᛀ
�j��r�Ngf�VL�A�nBb��8x��mH��﹕���b]�q?ZBmS���B���MԲPR��{,�F£�E{�+�e��L^~w��Df����&k����]��_��`$O{[�lo'�+@�B��|Ћ��j�	mS�n!�G����!�ؘUb��N*N�����4O/�w�����93w� ȲGNݫ�^
XJY��1ߵ4,�N>������K������2�Q�w��u��mU�����L�M��6u�>^����Rr>*�7׶D�&r�L �fW��y�$D�)�k��T�݌��b�VU�����,9a3�kG	�	�01�ZB�Tevuנ!�\ �C��{��e��d�y�E��\����9}Ŀ9�cS�ܝ�9D19��s	*�Q���b~���@�r�B>�=�Xӫ^03R*��D��XbyH�7��4��N~H4ɓ��R�'�A-ω��J����-~i?�����y��4?|v�QgMT��m��*�h��=&������|Bp��?��(	�Ĝb/O5��\M�r���e��4٘Wrš�0���9sj�w��H���-O�<��z���ˑD��?�k��텆��©z����*��VKjp��Z,��.i���0�CY�I�(���@�v��ك�o]d9�)�P�9����+@�������������L�vqH|5��1י�8	��l5'v�GZ������J,7��҆��dfC�����ma��ۘ7�Ja~`)$�`%�j�k [Bp{�����v�+(�e�5����Xpk����c`9�n9�v%�1���E2~{���amc�	_��> ��&I���=�bnBc�2�d(�l+��lY���S����<�w:�+�����t��7�}��wI�C���tH�	H��)��� Wd-��[�$�6�n�?�u?���b�,�F�4}����Rh9�N�s���b��y�;!�EQ�7Ndob�D�h)����Y��Ā*�sƆ�����Pb=~��G~Hh�	q��r��y)�eE��2��8�W�D�<J|Ut�41C���0{��u� 2<ʌ��a{��k�=`��ϛ;pg��w�����d�k5�m,\��ҷ��4�2��R�j��~#w~��������b4f��� .�;^��%&#���ά_�-MC�I+̀��祘��D�9��s}����g��� �s�y� k�A$X�����4#yMbz/����o��X���MP� ���&����8�6%x�%�]d��a��X����T��D��_�Ky�۠����*��qz��	�$m��7��aĕ��/1�wP��&f�b]>t��2u��UVAѶ�祹|�u�G�ŀxOe��<]�{�ܡ��Gt0�o�=�A����G~q�" ֳRˈ	;�賥V�CtA0eUlmI����R���{�Q��Cq�x'�}P�p95i�;o���3�����P�`�1��ǖ�|���e�#�JUC��$DS�j�a�������7w��^�e�4/M�'�6�n}��C�	&z�br��\�%�ċ��dܩ#n0����1j��C;��D��M�D�Y�7?���� �޿m����ʣ�E@��/�P����E0_"����k��0}�8��[o�/�����΋��*��IL����M��"؎�ظ}��z����"e�رm;��c���&�V�i���s�s!�wn_SO�1��Λ�%�]��u���3���M|����5���6"HM�����g��T�)v���]nsW"p��X��#1݅���c���]�	(Gdhu"�,a�\�@*�n���w��t��hR�X�m�.��v�G^��sNc�-0W5����dЎl�ei�Q��v��2��7��O:f>��KE�^�i�!�nk���9Saw��Z��`���2·G��gWG��?��>j��m��hp�\�O�t��ׇb�~r������H�����:�chnX�@y�A�x�P�����Kl�_�7Y��⡒�`��b�률�?����P3�o��~�G�˴~	b\�"|�\�}=go�����h����z���.ӵL�V����ć�Ӷ���)�p�SiY�UF#��� ݛ�y#�I�Vz�Т��$ii-ӯ5�62�z�;���v��4�li��D����$�u~H�}���_�����\�֤]Y[W���X�1��Iat:�a��nŖ��u�B�b����y����v�?�%d��anW7Q?�4G{�b�d:�K��-�>o�c�(��Ti��{BA�㼰��0��2�m�1�9�,�����f)@W���<�.��������zce�A#��>�K�����|�Wd"o��3�8oTH1U���x�p� R��ۏۥ����>'p(��-��-�&@>*�:}�$<��W=����F���7�ĵ47\�Ҳ�4��:�ׂ2jH�F��`�-J�����{Ӎ*���L���r���,����'��h&Z��^����93��d���{��������nq���6���ڧ��5�a}}`�fv#��:>��4��1�o�����
��&�V�V�b�f7i�F�E�y�Mz��K�59���Rc�٣
�[�q�zM��s�D�]1=�v?*�U���&����N�y,��;Xs�E�%g��-����b|I����^�#�����ν*+4�+���ZL<he�?<�tA��4�4>BSʮx`�X�k����-3I�D�GG@��g7x���4W���,�l�_�%��K��wO=���K�34�uܽ|[���,i���>ʺ���]�����V���F�e^�z��޶�}V7�^eoR,LC4�������^��Z�U7�$Mq3��p拝�AT��x��y�I��&����-�֋���i��M�0��'M��7����� ��g��Id�:��ݤC_"��|)"�JR�+ed���)��r�p������FHf�V�����ߐ�GL�,x��e���A�ù�ݨ|]���k&�q����N6����&���r�!���b�P�V��+U6�q��b�Ra_ȓf(�$�?'�`tWI�-���������#꘯��)҃�g�\���e��}�|X�g��Jk��Q�s��o�2-���v��Z�i���Qs��W[X6O���+u��x �h+<�Q��zF�9n�5b�o��XO��[�r��Z�n�ߓYfv"���X�h5�Z�Ѝ"K#vd�{����[>����2
�9�w�}�Ar�G����y)lح��ŀ5B�U��f���jZo#�����֫��rԂ��)ߙ�<(#7�إ�x��ކNl�����xM��%���E�.��/<�g8��;C�^u�s�>@-�3ײ\+6b���ϴ5M�7�$}�! ��k��h~qP
��Ϣ��A+Ӱ��,�먅�=�:�þͣ�"�X��c���*����>�t�	7�@̲
(��
����p*��\��dĦAb���Xހ��"\��������\f@A��-p �-i-T*��J�lnb����7s^b�S�8ף&��/'&jaVԭ>��I�ǡj��4gA6X��
��#߯��ƼS���Հ�њ]k�KN���x?��XU�c�4�}I���Ț���w)�¾�/�ă�#y�_�Oy�v�<g6CJq�,e?;s����a���k(��vU�p��QM>Z����9�]���5�y�:&;����DX��1G߁{?�$����������Gl��~��T8��Sv��I�d��x�ß��-pTW�>R�$ZWt��07�'���Z�]u
p����!L>N�⚿���З �S��<[�6�j��v�?�O'�Z	,���m� �����9�*�Ք�[J3�x�Q�_��!<Q��=��{=e�H�����z�/FW�O�>��:��켶/I2��q�PA�C�����)2��
D��7��`�p��j�O�R��-�:Sd�$ŭ�,��ܝ��k� ? Vm��6Y�"V�H�yZ�=Cά����P���U�r�}�Q^?�р�$�a��;I);��[O�I�ߙǟx�(3G-sR�g���z��B>sIu��k�H'�n~bM)k6w�W��HӁO�.����5v���\�n��qC��Jة�`οyJU���*d~�,Kc1ˈ��	��������dQ~ؘf�J�N�H�YĂ�3���ޤja�@L.u4�Y�Z3�&C�ډC���m��Lpϔ]��(�(q�¡�&e��L���PB�J�A�
vz�uS��Zyӱ��b�#$��6�M�lc��[с�6{�
n;Aj���F=רH��yv�㒖�*RϪ���&1������7�w�S��eJ���9�|O � �1*n�$E�/�ϲlYy��0|��e3:��0t�	.�����y�N"n"�U?2}����;p��;y�bJҘ"k���M�be��C�*O1�(�q��0M��i��g�6��b�g�<��-͋��&�X����7�z0��i�{7���T�-�2���6gx@��D�	��,A��c�� ����Iy_�+�?�W�@�����t�9�n�����SM�7S��hWt��� )o��z&4~�-��bWc`-�B�w�����ǌ���f�� SyD�^,�^D��������S\JH/�etB1ꄢ{{w�n-�@π�:�D�������2��o
�=m��-�Z�S�����`��y�u�X<�8���@|a�WZ.����3���Rr�:��!K�Q�l�	�0j)�Vܴ��+F��{�w��;��^u���p���^W��e����Y����o���g� t��|K�=� ﵚ��k��p��(��k�����s�~��H�~�>���&X��))�L��r�+2:�v�{�n7�h�� {v��M8ы�ް���<�B2�g*�R��y�'��q�8���>���v6է��9��P���q��jp|n�~�o��T�`\�|����Λ
m(ON`�I[���'��9�H� ��[g:��?P�C�L\�CRgT=�o+��#��t�[#���E���-���I�y�W�U���A�HVټï&�"]�a
*�����f�߿�[�%����q�K�F�F�W�	�s���Q<�]��/s�2�䴙�EW�����X u�P��$�̨/F[�b�6��T:�`��)��Ŀ�
\a��F
�Y��e��5_�]F�m%N�v��J��5�`�nJ�hg��5���_;.�-�����SQ��-�vM$��W�dKB785�>��:�X�")ꮌe|fi<͇�1\�D�m���+��<�f�PY�A�:�	U�j���[�t�ꂯ`T��*����8�̘K0m�Q��V�s?8��B�1B�=��ܗ��0m�Rv%w<���f����29���:>�#;x��Q�����f���@J%Kڰ_.jk��d�+�>^��tɢ��1�䄚������)
֖�ϟ.�d���>v�0E\r��W�T�-�d
ߍ�Z*�#�� �"��|�g(�U�Ѱ�����T7�ҫ�1���G-�=�3QwVНs &��X�ȹ:6�h�1]�7C���p^���&�9�I�]�� c�L����p�߉2��QW�x�-���Q��<�q��VT�[5��8rs���N���y8�t�"�{�!��]k��ĥ�z�Ϋ^9��硏���P���	ڦM�Y��5�������KC��>.���j+���r��e����UTS$G�=h�4e4OT|�y*�R7�%3LS���X���e��.��9���+�|��}:[C�c��aώ?�ð��I����[)-���D�#��v4�:9Rk�Dw5ԇ������s\ӎ���A���-�ŉ!{��<��">��.�P�<�"H1�$��Z������T�� V�j��}�������Y��% 5�HJS9h~%����ORW��*)��@n��.�%˒�x�"�`���D1�Vik�� 2�qӃ��A��S�����a���#pٌ��Q�=�!T�$��`�j�LGE4��x�͢b��'U�p��Q+.�Ӧ~R��;ז=!t�_�3v.�yyV��N@e�`�B�ݢ4<�)��B��^^(�p�x&��Jc�&����Ԥ\�>�mI��p'3mVl.���\�M���Gz~x�����>ae<�$�j����J��dm�y���i���j3����2�=(>���>��d�:�Ӊ/����vȏ:ء���&I�����Q���i�j$��������AHB��ˠst���t-�ϋ�x�����F�X�C(O��I�M2 ̗�����B���������g�����$L�.�8(s�������YZ�>��Q�����l��glS�^޼�p*��K���}!+K��p}N[;��C�re�R�)����e7׼��l�@8�e��̗���/�ǵ@�7B����� ��&�S�7�~o�o��AO��/ϻ`�7WϺ�IH��^/N=�[����	�2��E��Nܰ�x��������	/#h���Y�Ӱ���Yh�|�Q�����ZbZ�LT��U������=�B8^�3�C���&I���g�7�YR�q��n�N��r8���_�Leܩ����c&E��1+Y3��GC�J�rb\\b�Č��x�#��8l�	�RX��7l���9z�[�D���7������glNos�f�` �^h.�������+����w�J�����ǐ�#���=5t�h;XB쑖�6#dM��s�[�r��'�
Y����)R�?�P)��:Qpt�c��(������S�a��]�/��K��<%�����<��`�������uV���;-��v��s���}�B�&��I�Wk\��#��sy}�Z\L.�1�==����q]��وD/8ZeFw�8*��)S'φ�������O�D��v�h��D~��t����S��@℔�a/�S�Q($���)�X+�Xz~����$��Igq>3��S�K�8��x`e	��Y*ܮ�#+�<X�&����e����*(
�8�U����w_���l9!w?-i�&Km�kF2�0��"r!Q�{:n��f�{xs�"����b9}�ś"��,md&\�}��"��,2�(m��<c`N�����>��k�f3GBQ�e)	�!��i>A�{
�Q�f.����6���5E�}m����d�����r��2�b�X��80X�@�(|h���fQ�I�Ő�p��%|�����B'���5w�g�u�����)��(-���N>�M2�>�)n
��o�ǐr� z�zsEZL�aU`o�"%o����"ܵ`�yo�j�w��! V�Pȣ1_ja���P�5�Ԕ�X�뿘���-��� ��Do��<8S%M;�\$}��T���㓫v�۲�Ȣl��;CQx0t�J0xB��W�{��6�?S|�ƽ/`�3��5��B������1���}�|܍[���g�� (���~��'�i� �8L���=��>�y���{ɯ�5��#��ވ�6;�Fq��d�)L�z]��s�¯���K��T �#j�*bq��[�"G�"����i��	��|6��}U(���F�|���.!6n���XU���@��ꦛ�R���d$B�"A�:iX��������c�=�RႶ5��� -6]Ai7�w�^���`���R������
�h��n/�Y��{�e��r)��4 �!���t0w������L�:��� jG=a>-��U�	��PďN:��/ҥ�"f�* ��e�a�@�=-5$.��Û�ec"0��0���2�^��H����zO���P���#6b�h�g&���@X��TnZ���a��\E��,�Tm�����́�I&�5[��!9o�X �El�ĸ�F���h����|F$�\+��&�zĊn:��A�D�����(�j����#�g%���8�܄�Eh{Ʌ��7���lYч����¦䱧	�467c�7��|X7�!�3&�|�������.� Z>'��8�*�Ww��4nSv� �섿�[��NL7����������o0��l o9} ��]�S�7�eo��ǄPkV4/o�F�Y���=�5�6�=������~�ɣc6��]�ɣȔ'��ϧ�m{Hd�M�_w�R�IY,��.O[�Uc�&�x��N���A����f����+LI��P�$�ևiA��v���]h6*�et�v�B^��~0���8A�|Q�����C_6tZWDGRH�g�v"�|mL�ߗ92@�v셧FU���,Ը��|Lw���T2zk�Kd��b�,!P���b��,F��z�!
����~q�s��Ь�����>dh�9͆��!هb&��1�3�z+Ϭ�@���0����@��� .�w9>+Hq��t8\�YW�N��IIZʂƥ���F:(ԲO�,��z���L�$�/׀�kj�A�!�@�w頗�l[۳�\���z�ށ(�8��?��2V{�0���K����jg*�Ә�N\Qc~,�)X<ZaĀ�'�OUP�Y&Kŗi~۝~��b9�	��y�Z!��u�.\X�(NUS:�D�~!�+�N���"H�ʆ�x�A�UC���DJ���L�y�����l�������zt���}�ڼRz�$e��'���$�_���cH�QK�z��k\۱f<��z��Ѣ��!hH/ʵ�I����+�j���/$1��m��Q�J1yPH�hw���,Bxݾ�u�p7�����bJ���c�:�x5�í[k{�T������"j>������� �SP CB���O�6�|A�4� \J9}�*��L�W�q����sX��Y5�85��H��<I���l��^���a�}���'���ˤ/��㰥$o)�`t�lV~�T���V4��ɧ2��M4<�[�`9{P�~�Us�yA�nک�ch�QO��P��ǑDV�5S��)��4�g�ZrS�JN������� #�x��m��d!�����X%+�p��yݥҸj���}<͹$�3�H�RU�x���c�=7~o���-?E�!����G2@�[�|�
0�Ɖqd�x�$�c�tjl���R"�*;���\�I�C���}X���L����A�U�}�V�w5�ѳ��8D�<%��� �[��X#f�*�"a0Q;�UۯQ	�uB���S��Lt_g�^1�W���������Q�ǒ��VgUZ+d1Gt��	\��gA�'��]6��hv�e7�l�@���3�xQNU�MC��,ފRT4"�I,gr��D��҄ւ8���]%�BM"�'�g�Ǜ���e�Iƫ8�Ƶ���A'_�K�-�6ٺ _�WcH=Y-Coxt�"�@��RfV&��Q�����7j�@�颰��E/I!Z2w�����i�+�O�`j�hVoIZ��R�����]�X~�n�Չ�@�g��:N��٧�����,��~a�u�+A����oYe�(���i�%SJ�YJ" �I�+ȧ�e�]��刢��&�j�k��ę����{1<�e� 1�Q��O��G3U �ח�ΗZ�ڣ��Uz^�����2�>��W�E�����i�X��������+-�r�t���p�¤��	����5��f�h���Or�+�g���d��������0I�������6�;]ȅ�GN�æ�7����dR[[�uo�K�Sh�@^�򘌚���=�D���,�zn�0u`���@3+�Y�-�u��-^�)J%H!���{ȹ�3���6f�WJ�q( DI��]H�o�R�sZ����P��#(}�R	C�k��9��Y�i�a�(հ�U��A�Ӱad�5V�P�24z�2�t��S!
�@�s�e���0gw-�����o��o�x�3���⅐�y$r����Q�I�S��u��@�@$4�)�"#�h�{�ls1��
LJ3H��ϕ��YvJ�f��ޛ�gdmL���_��	p�c��~��o��0>��7��EX��co�K`f>H8\����W����d�%(�j�S"w�ZX�f���wVyCN�*[[���?������\}��\�ʷ�6:_Ҧ��_�Y��ϻ�0����T��V���li�� �e���]�����3���~����:�$�m�D{+�F�z�)���}s��߼&�V� �l�$
q}X�6�L�JMyn�P*�~>ͅg7�1�)�8{Rp��IB.�����Bb�g8�u�FlE���5�D�����-Ce0+��w�/��K��}�A�H{��Ԩ'���b77��xNkjfA�X�x;2LS�A(B��7�:F6:?8�N�H��4\�- �s0X�4�NG���èyQ;V:'���s'�D>K��vY�\А��e�t�T��=p[��V�AA�A<�%����g���]I���jh{� C'��U�x�o�`����cw��p��A�G��_����H�w���w��X-�V'M#�A��5=Vj�i��WP4�_�;�|�ɊKB���yh2��MuG�HM�9��$ q������nMY�K72�j6����G�P"�
�g��,or��8\A�:��PF��=�\mv��q���������g�Qe��0@��2V:�!���Z�#�9Q����
{|��7Y�Nǋlv�3���5q��m��I��moq�|�Z��LH���&�Rqc@"�t��L������ŷ@}Q<�B�ø!�"��鍾�d�E[�|c�*�_��jn��1F��(�:�w��&RE��#Y�Vc��X�r��i\}M|�i�e=-Js7��� Z$l�܀�0��#o�����fݷ� 1.�3B�,�?81}�	��j���1�7L~u���5����ۢ���[a5� ���g�pe�y$�Y�wl��*�k�GQ�Ha���SP"CР!�y�(E@��y���~�;*f�?`��Q[~mc���ʛ���m����k
������=̓ƃ�A�l�=�&��$���S�����A��~.��5��i4��js����w�}�X;[�����
��σ^P��~�}�º$�?$K��D�Mj��ܪK^4�g��E�� �T�)�)\����U���Ow�ý�j�h�uP�`��8TQ�y�vq�[���r�BP��JX!�O�@`F,�v�H�`��C�4�޽�UN
*����X�1�vO�z2�%����B����І,�&��g�7JI����v�&(�T�:�V,jw�Yz�(I��u�44�A����W>B�L�&�0z�d;D���%G/m*��~�h
��a�W�H�4����}����m;�^�X:����9��"���n��J��(�&>��"����W�T������a�Q���j�*�~����q���,{F�1o��*y�sM���J {{��Ȭ�`\T.C��7_���>�녀w`\�Nĭ���hٴFi?pp��T����VfA�[�����.��I��(��EY���q�g9�-f����8S�$���x�F�|�(s��䦕�3���w��k6�7�]������1��jC�x�R5$ŕ�kJ^ �e�[
�S�1Q����|�2��QA�r�כc 8��H�҆+N��«,�-��ϥ�4��4�M�P:��3A�	��_�'k�Cܶ��%�A�j��G��@x������%̜r��]�ᚬ~�d�"=O�[���t� rQ$��G[q�(�^��3#���"s�BX���w4U�D,�VJ��㒠Ċ}7rKx�J�duQ}���%eZ"�J�\G���fX��:����\��Mu����^���+�6��l��j�y=
��鼙�x�xD�	b�͹��G0�`L�Y���J]�5�)�p��Maˈ��M'V���?��t��S.z�8�nu}0wR����#Q3�Y��L����s!�����3�}�`�+p>�&@��Cʲ;��7aG��i��B��$�v��d��	9AxJ}�#����ڱ.��9�oL�
��F�1��亨�~Asy�	�A�-3���*4������	&@ϡ�R��0TG�������Ҵ�#R "w�K���΢  � �I�A�����9N��N����9T�C6iae���'&m��^E�7��w�0E�����c߇����[\�COĵ�xը�s�J��I����M���Q���_C�	u �&�'�^����������@��nV!����J�2������H<�47������`a�l�ء~�?��=�s��,,��Ū[8!��z	�\>g�f�p+��g7���;}�є��� z:YÏ=�[A�G1%��M��P���>����\Ek���i^j��-y��#w$�팙՝;oGa^�;<��sk�h��w���?��Z���n�@�����Cʽ��1�?e���K����\pA�hRR1*d��e�kN�D-�U���W
d����u6�[�SJ��i�fD���5�Hp��S箼��A����\�
侗+w��R�e�!߻��_�#��\�i�2:�a#u��_��兓�|������%�k	�$�<Gءu�
�����D!-5I� zr���rM�Ry�R@�!�o$�>y��Oў��i.ï��$϶��$�e���~��E�"��8�7���sI���
N>4���gZ���V�Ce}�V�&����~w��qAto1h��x\���$�,�zOC-�[-Ӯ F\�+g�I%a!=8��&�6șᯤh_o��D��G�@���om������p@4$6�^�qdaZ`X�u���U%��pJEj�!?E!���Np�����Tl{����yR�������f[�-_ל9��a�Cz��E�3�"	�
'��7��}A�*�؟	"�$q	������1�Te���4n"CN�j_����Ǖ9+���s_ȝ�l�ʁ{meӆ�~�(����h�����؟�
I�4�Q2g¤���V��	��\/��CQ�hr��ͮ��j�����e\�k�)���-�!�Ѯ�`i*�1SX�(Z����sÒ^����#�d�c�kE�H�P�5��:ϝ'%J��3��g� ��kM�IX�+Î�Y�ҳ��
Jtn.���y(Q}WƤC1��2��X9=�kJS�DyJBLn���"�8L�<���������aӽQ����{�6�D\)���P��NtUa�q�)���}�d�<���\rRg{�. R�>(,�e����H�1�����Ÿ]\E��W����������@��gN#�&�'8@"}����<�jP��\�L[v����&/���*�U}���aI��#SX�f��Pq���f`x��a�2����wk � һg��z_�V�xk)T`����$NA�lGN��G�ND�x�+bM�R�_�*]	9��.}V��L!���hW�+�ť"CՏ�.��8��y����_�U��w4���H~�o��
������_�q� �ڂ�^��~���9i���T��"��!�4 8L�)}��w��/Dap��m^�j:�̩�2�U&�:A�=�#}��v5�W���B�{G8t�zl�D�P~�/_g:I�3V-�6z��6Sp����#s�����Y<���Obw\@US�/Y�U�g�h�E?ş�q�	�x��*��������I9�m}Zx�|�u�m�	a��Յہ�mM�L�wŒ��(uR����N{��)$�<s
���9�/d����x4>�� �\�ZFR=�j�π�~[��c~$�*/�-��r��W)E)V6���;C�r��1�.�;���h7hF!C�j:�Iۭh�e���V������5ik�į����3�!�݋�%`LºP��;|Ű)KԷ,.�&�:Ȅy؄������K�;���g���cT�~��l-��Ed�G�:���-%Q��,��l�Wo�҂\����'Ƿ�{�uk��&�}@�jE2!�x|h��X@����B���hzp�j�yx/	�Z���N��n�@"��_�4t3���Y���D��1�����d�ocRҜǛ����9Ƒ[Iiu���ώFY��|�`�ބɱ{c���7���%ᖞǲ��t�"��ZCO��)���z|�.�������I}�	�=��f��LՓ�٭1LV�HR(V�Cr֌�M��r}�4&IٰE�(dż�;��o��d��^���3�S�`�^�S�k62�'��5�����5����Ń��*��r�`��|���C��g�Lu6��K������{��VL�����W��g�%~�p�nW�tLi	�7FNd��?%M�p��K�s���k���Ѐ����(�j6%�g���"hmG:X��'4RC�Q���Y�9�>��Nc�5*� ���Ú���qj�XbR���L_�K��Pe�"����cNv��&�d*�E+ �����T�Z�>���<�רtz&��Hjs�sH�\Bw�J�]��fr	'��)�� �
G����W�n6�G��Sm��^�Q<g�6G�%"�,��&L9��q�'�x@��J��mq�����v�'���A�M5����5�ŶZ��@i�L��Y�67x�9��G�$����#(���%M�	�)#KǲX\OT�f�` ��1c+����A�ǲܘ�L��>i*6V�=Ĭ�͐�paS�'% �3r�O�û�L�x��끟G\���QH�*��@x#���Ӟ���dŪ'��YN�.����t�]f,t@��
 ����u�4�Erί�Qz�n�������2��t�)��c�Q��xQ�hG��eM�+�e9�D��O$��~��C�fu�M��9�ֵ��ag������A�Yi�c�t?�rS����n�<L�R�O�`������ݯ޺��<����**������ȐF��lO+5l���g`\��e�d�b�v��<���>���������_XX�\i0!ӎ<X�!�Ա��k�<��M�#E1J�]Xz977�>�y`���=�3L��3�4�󡘠�����ѱ�b!
C�g^���m���Z��ڙڌ���n���� ��b�ɲ�bv\�	�:�>���Ny�Ť>�a\��h�*�`Me�*��dzSMH�?ֻ�����y�bk������Y�}��_�-��P����=v�D��B$�Śl�Q���WN��oo�T�`Ƈmn�\e4^�egIvȂ|2��(0yf ,k5���nԪ�V��#���gʄ�V��3"u�js�u�HO\�m��-|L5-�Ӄ�m�2f��r��q�=���n�}�b�9����Y�Sc��	�]M�ipkXc<�IF:!˒�1ֶ&Ϲ�:�R�Y��[�h]c����s���- R��� ӛ����Tt���h��Wr�S�^�]{k����2?~�u^��%�M�o�����������ÖR��׮El���7� ��xm��9�!�8{ @#J��E�튘�����y ��l�	��?���]FFf�X�:����nnO�<f���eh����	�]�k�� �����N���$�M�a\��g�04ϑhm�&�xNV�ӵw:�\ִѹ%�Z���"V�������#p�a�C f�~!(�?�A]�KQ�=���S���e�"��.���h#q�8f JzW��uTH��o�v����]~]�����?�mH�:%Xh˧ ���U�:����7y�߀��v'w�	u��.��ˀ����=Ŝ?�y�Ktِø�$�4h�ú��8��K�l�ȱB���\���/`��S5$�B�EE�Ap�Y�ɖ�ܖ �Y�w���g�yt^�g�YiT���]�Q<��. CwUٛQB�ս,mἫ�O�W�W�44��0�.	[���v���:��bSs3�v?�pq���?���5�'pT�����~��MϪg���>ZܙC鴀��{r�=_�v&0�}#�������[�{bh͸y
���I�(m3���kKs����K�b1��]�+�e��[r.���HC9���Bi���Ө��(6"�b�q��1\����<����I!�]�d�eS�@�"D�>�mi�m/IJG��1��f���K��l�N�"zc�8�{�S�c>��I��Da�r��b���m��c&�o}hٺ����Ur-�B��8��q�+��*d�V�ȮEf�Th��j�DP���!��+��ܟp�%uV!]=�����g',5���>�,�G��1c+�;�qOq,�\���[�Cb�p�7o�@�B�EV���@<^����E��~:�7�7���Q��u�рB��%��-�Yrs������`���E�ȅ�~X�WXY�T��~d�Ma�-��85��w��YmkT���:g"����(qd�������<�"�S"nA�+%C�?�쥌�pK�p�`�� �/�Mj&�QۓΧ߽p�6Q�h2~$��L����sy�6��Ȱ}���!��j�}�ǠƾƘ��3MQ6
s&.{���PB�oe%�&x��yk���[R�vǋ�q��Vr��V��ayݸJqrl�_}(�V��+{>=}��eA��5vXԺ$G6�R��1k����B�i+�jm�p{��ȌgH)7
�&�+�%Ȥ 
�0g�&��"�]1�� Z���-6�̩�,�h��d�1A�;�v��?��-�<�J�J��a�C�����>%��Pgu���*�=�ڇI��G-�6��QR�z���Z����?��,pLH�"�+9Je��Nr�f��y����i����Hé���@�ƚ�i��D�4��e�	���(�K��0��n�?�ҋ�y�!��,���B��Q�5�;�:��������'�
��'�@
R�u�$�9c�iŶ�|��(��� ��HhN?���S���:��ҥ =�Rk��zz�.�c�m���B-��^
!7r.�g:��� �E&,�auqW��y����M�uUL��)�^L�i���6��ľ)�wܧ�{o�=Uv�Pi��n�"29�Vq$PR3��Qrf.�8_q�O�s��r����k�,U�6&��ؑ�c�9 �4�xՄԾ��]��~E ;�H0��-b�Cr
H�e^���T"�N��A�bq�T���\��j<�"����� �<^�O�1�j)Ʈ�1Ec�N.�N�ܞ����X�����饏!��0����n4rxNg,��� l�v9�E���Ft�J}�\.|���t���_˅=I@���eeSv��J�-�g����b>�gߧL����z������i0_�bs;+��"�:���"��h��F��o �z�G����`Ъ��j����d��Ei��0��z��h���2��<�����Ҁ�j�σ��{qzUa��Ψ�����U1v�v��@��/G=��V�:�`*�p���W�Ϟn -΄+���F_��w�U���4sa��U��@d��%;�Ȧ�cSJ��WA��+=2{<Ʋ���53fȵ�n%;� R������g��dK{�i��2�5a�=�������o�=��j�ߠ�B���@w
$e68�/SM���'��.a�����O�:P��a�vc��N�_4l�lf�����"������kD8�H##�'�k	YU/���@(�;���G/�G� J2L|&bH��sYCo򈈏�2+o胶���O�������P���_��t����oZe����H�a���"#���:�� �������htR��?�(:�P2te2���N�����eâ���~�B��.����ex8�3�B$���,��թ�F-e���P���)�Tr��{q�w�穔�15iʓ](� �H�uB(+֛�H�AaY��8n�.)�Lg�����S4{荍��%H�u�Q�ϲڑ)�L���%��V˲�����1� �����2��A�CDi0���p]�tei�ev_U^0���~����̯y�X�LT�TFF�M���~�,�(^u#��UI:���>������m�X�'�Z0 ���Φ��� !h�h*��K�r�
�U8r��P�f=�"���_�ぉ4@u�c_���r�N)C�8�(�q9���vt�?�cf��-�4g�?��j�O{t�i?����٬C��C�@GR�Y¢���Dn�V�429G���h�	����b�J5Vx�9[�x�����N���������ޖ�6����-M��-@ʊ�6s�:�U�&���6���5�M*)�N�X���8`\�]�LW9�7_�ڀ��7���}��7{1+�U����ݓg�cQA8��"SA񑀒�Քz>�V���,ɵG����[�]�	s�W3��Q�v�u,��f*������JlI�c���%�(ܨ�������8
�h�ڗ����Tx&x_r/�4�:��(�\���VgKc{|�*%�Aj���9?F�L,��yD�h�����Ne;�l�I3+ �6ŝ���[�-��-[�$��*�������W�Z�$�;�j��d�5Ymn\x�Bj��'��-���

j\Ae�q�j�s�O?�BoV� 4/֮R�\"BLs�Q'�;^�y�|�p��d~���|�Js{r�|�G�`9�Bט��_���������B��<�?�T��!�Y�n�7٨���^ŁW������9$,��������������+��+^2�}{t�Y	�:�;m����w"��7��*ZH,�G�=B���a�MD�L�9Q�i����Ja p.��j��$E�V]c������a�C�W���٠��-0��J�<A�!Ɋe�?�`Zo<�B�%��j?c�����>�����c�������{<�Hpjs6K#Kɿ�q���KՈ�h8 K#y�����?tn�	�8t�g�	���2͉���f�7����i�TW�#sb2�p)F�!���&�X�u�.aGd�� �o���}w��Vy��k(���.��
�!@�*��{ޓ>|I Q�P���q�x��h�˷@��?0OR�ќ������mGtX�	���h��t�1���<l}4r1��%�I�_������u���Y��K��n����Ѫٺg�g�U�e{u�U�$<�%����T�X��q����GWV�!k���X`��S��6k"g*u�����-L��M�Q�F3��%+�GD����R]�b�4L���� �h3�5��e�UJ���S�lR�+h%mȞ_��.���Qў�����0H�#d�|n�����Dj5@�C`O���}������i���pN����'�Y^��;]��f�}���[�;<+�ߠIxbr�u�:KGp���;�d]��0�-�?�ȩPH�ǎ�?OuR�x"x�:�8���I�k��л��6��;l����a��Iu��a������-�wJ��ch�pTaB�Ґ�W�k� ،�9K�ք�c`Q�%���!��֬�-K<�rӧ0?��iC�P�^�ކ�c1�"nW��K��%E���z��!�+�s��G#dp��q�Yz�JS���F����1q���Rp���x�7 ���6�h.YX�0e@]w�y����x�#��������0׻��b �թ2�����h�}��'.c���6Ru�s)@����'� ]�KR�ƫ�y<�T�H��Fˡ*�@����5I0�*�d��x����9�-Y�ڱ8�`���#F]T�#�� 7�ቡF��a�+`�	n��j^���(�q�9¨��������U
k��YP	Fe�8��,��o��� ��Q�8���ᦈ8� ��_���Q�`��ta>��`8�N
x)�@-�L����%�{h��ˬoDQ�� ���<�^J��@`4�^Dg�"V3��G?�녔� ��uUV0� ��Mt��p^�Ɖ�_K������|����f>�L;b�;��Ei㛴>�3����Z�h06 bx�ĕ���0N�M$kK`>_7>��8�(#��R}N�r���Lœ�=�@��&�(bZ}���]�xp@� �\��Ȩ�p�x�*Ж��X��M#q������T��Xrk����*�{��d+���0C�\�٥�@@�N܏�eͨ���q�Y=�g�o��#��)�������f�`�L�vl��ERJÅ决�_PjF�c�����<�9E��L��/+�[%:Tv����DǔU�$�E��ݩ�[�и~=�5�P��Mk(�g<^ɑˢ�O�N�I�^�?*��a��
g$	{��`G�����A$��%�ȔD?'�B��@���$����c���&���3(|M$��#h�zŘ�IF2ma?�`S��g���	x�Y�H�l>	roh@ћ9P���e�¡�sz����6��Gݫ,�?��D�Ս�{��Viu�.�0$7�)V�v�V �œ}���á3��f��x��x@�G�BW���P������o�艹�y��b�I�1�i����Sm����Sa]L�[o۱{v���Vs���V����Y��?��g�v�_?˵��Zg��{��O)�!���aM�� �1j�<V��M�H˫�HYS�%����g0�#�������"Զ\ɾ��d\�Z��"�}F�����2�w��4���q���G�00�9P���r=E�i���T\2�KR���j=��A�u;7�-"ĺZ��?��NVU�!{�y�We���tGe�`��0��z�:�+�m���hOT���ϝ֌$�bl��6ϑ�>��/��CYr�#��V�b�N��Ld��I�kX�V�i������
�T��Ř/$Ґm�'�mOTǠ�Q�"�D4���p�����Z;�mc9;���ʢ/�F�IxpS|���~�P�݃)���LA��(b�5�d���s���2�$Έ��!���Pu�wȖ��^$ѐI)$[��a�a0�u�؎�~8��G�'�uI�
Áˡf: ��&�|Z�;��=�ڷ���B"��z���Fə}��?�=�tS(�L]s�ONm��t+�+�z�N��\�D��۬�r��.k�a��f
~�8�:�?"3�ᴜ��ڀ�ʾ%:�G�{�4n� �<(���x�#9�o5b0F8�#�Ԩܺ��B$B(H�'4rfҼԌ��t ���T]����%Ӻ��T���1
���i�TE���D��}�V�Z�(���`��F�e�`Qү�w%��z�؋(��M���;;Q�9#� \"����H߶x�E�G�Lqb`�0_�gh`b�}��N�A@�G���6�KV�у<��I�qp���p��^L�z��Ţ\�/$��+�������2"���A���U���{,cRFc]'���טSj�%�B÷�OX���hoIN1�ks(��H�W��0��l?m5���q�=A���j��7-��,J!�O��Idb4�gJ�AJ�k���S��2����u,�B��`�:�jm8�Us���mu��@��3-"��/U� �{^�!�&���̚\�?���Eh�g�#���osг�9�	����!�c�����NIqa`�eM�J���m�nO��E�闏;4H�j�rJ��؉����$�s�@҃�JMɪd���V�-M;ɾ�I�av>���N4�G'��cN&<��>F}�3����_E����7��"��|+���U7�7��<��B�+~�3����t �-�d }��+I���ұJ` ��!��U�Ae����6�ؐ�>���SF��1z�<�7n5�R.&6�bRϤĘ'D2l����93.A<ݲ��&вS��������D(E
�r2L1�B�r�1cg�(݁"��(q�f52ܯA�qq0�hE8iPsf��B(�1�~����6?��Mu������OA�Ѣ���Q�]�Fb���+,�Jn)�n��Z��<}{�;naöl���H"<���
��4n�R�����`Yx�Ο�T���
t���ށc<����=�����$����<��Ʃ~��y���S�<�Ę�r9EUZ�V�]g���9��[ ��vN��YgQ69��R༙$M��f��?'"�D⏲ /;��J��(3+*����������x@�OW �(7+m����rt�-�/X�Z�������l���||�&�S�4m{*ܪ�����ѭSΐ��_��\itBJ��j�T���E�P��Hz
)B���JZ8�o�6�#��f������!F�p�6�C�z�=~ ��pq��חX�Ͽ��D଒�Y��� ����LԮwe���d�E��Wo��,��f��8꽧��J���s�r<������F�r<�] V<�����8�7����x*0��~M2[��v��gcb��ç��oHݤɂ <?S�fma������>�R�LK���0$-T�����Y�( ���z����V}��ѦK{r��Kc2s�ʗ��` �¹Bڽ��$��"�4��x�������ą���6�_��_��b�����M�H L�8�wus'���egbe�!'�v��m�k�Y�<*�8�bd�D��\hg�~kL"�W�,�/��}���U�z<�Ot�qD�ۢ/��q�$��|x�D���T�(&(���nj�h�u�h��%-?�5.'��WÞ*�ds�������8 ��Yݗ-~ׇ�|,�X�tC]L��ڧ����v֮Ha�H����\��>c�[*>Z��N����#�M��
�i�<u+p�� ��bx����u�M[�xټ�2��赏^FHT`Gd�mu���*���%^\�_�C�nV���`�BU�[�F�B�� ���z~b�&k�;pSkɡ��{^DҀ7Gj��D��ؓ���.�ſ��ޏ��~��X�%��*mn���%�٨xR1bb��?�;|�h�f�G�A����v�Z�]�e�Wc	\�v�r��%*H�<��/��¥c 	rȋ�7�hY�5�q�mͧ�z�ܪ)eH���Q/Y�S��S��D���]��r�eа����@$���b�^S���<�Z�A��vKT�#(��_�Ӓv�[����V3#"�X�^�)���[�?ƧL���^g�+q�7	�l>~6>��s�����,k^���� �;����3v�u�.�+���)��0�0>oMl�J�����T�x���R�F�V�t��_�>��.�ꨑZ�D�]�1�j,����$ �
=$xb�C�gNN�R���-�굁�5M�������<O�u��(�ܵF�U��u�3J�:uXp% ��z�[�CG�^l[h�� =�b�����k�є:�$�G���W$'˷��Ҡ�x^�)�L1���^�\����:���Ndg��_:!:п�)b��L��I�<��%,�3U�K������3)�����@���:�����倈&��yW���jg֋f�`��y"����ݟʜ��������2K�%F��)G�E����?ލד�i:U�����2�~�[��k�n[M�p�b�޻��}0�Q�!ͷ5k��kȷ���2Q�M�����8 ?`��Ю�Ε����C�r;�w�����΃�MA�L*p�A���x��oэ)��[	^�0�H�/��T^e\d�4DٿQ�����XC6Pe6fmY9h�Mrd;eK��Ȳi�k��N�4!�D�^WW�0B�>��*���EP�yH�w�$mOF7ͩ?6��4�hEb9F����%��ҵ@���&��o����^RB��wsni�J0�Խo��R�;�$���F���XFl�bL2�vj]���l�қ+ޚ	0�TZy�����+��ů`_ߑ�r<?���2A
��X֪Sz�@�c"��c�c6[����PW�-�.��jw71�9n{ˍ3W�;A�04����V�D<@W�|��2u�	��	�@��2X�2X)�C�o��,Ob�N��K��:�R�\� �	�֢���2���^A�o�����F]�8�I�s�Ѥ�_?���칭�W_�|�6Yz,ӣs��g�l�cU�����`;^-/�Ea�����i�'6r��uK:�%��6_��qo\�K��B�Ұf�t�!�^ ����> ��c�$o=���^����m]��[(���~�l�+��N��w����Ta�;2A�^��[�h�oLp�|r9:7f�?m"vh`��z	v4�xF�`���&�R S�AS�YK��/Zי$�X�e���"���"�)���mu�/cb{:�vA��甝����I�*�r��@�~A��!eS��w��2��]R�c���K��;Y�J]k���:�Q�����3=�����+i�x��$_��t���K&����ʖ�)�T���ö9��g,�ge���A��IH��v=�������G�aN\���(��-Z���Be�g��]��na��A��m0��Gwl���QTج*��kcڱ�k��g0=���h��[�9������5�w�����u�ĖJj�o�V��ر��u�>�ǲ�!�e����L����@�lOr�v��,S�����G1�"�^��`�Z.O��K� \�w5!ԟC�q��j��F����}Kh���#`䜻k~�# 
_6~r��$39BQ��e	Ȃ�Zy�|��ҁ�Bh),XB��nW����H���?�u<a��kA�~���n�>�{����Ai���g]���!�N��~�w��)%�y�;>(�__(ve}�{���G��1��������h��p�?��16�#z�� �;�w	%I��q+�����)Kk�3B	���]�ԏn.�s4O۪)��B��F3Aq78"�g1;ŭ���, �dZ�uM���*��V����%��1�W鎲�)�;��M��J��W�ǹ֣C�ߦ
>	�@�#P]�d�O�����3d�K;�$���78����b����த�(��>��j�V��S$�ݳ�V>a/���K/�h<���Ɵ�ѦsR��(��%s�8��(���O:�r1?I�X����;~Oi��oN�P��n�kn�Q�{�z��?b����
��Q5��/���E�����mw��V�C�$��j��=ĦK8k�9�#f�I��J��{����tx��LR�������E����?���-ݒ���)��OD���G�ā&��㎳������& 3m�@SC�B��U�����Hzg��UwE��&�e7L˼}�
��]�6�ه~s�@��'�:��O_��ا%u��}�%@+��Atc��o�щ���۟wF|W��F�hRhfq�T:_��U�j������SE}h�M���S���/<�'8�7�ީ�]��1��}��)�[ӰRG��-r�'㩛��,��Ͻ����~_q \�M3��e�C~���UI��
ȤJ�d:m�~-�L�~K�|��Ԧb0[M�X�\
pi4�z#+"$�`�wpb�|��s��������F�9���Z�NO�Cٗ��ZO-�2K�+7)aa���7�U��)�&ˈ;.�y��,j .L��u���QCn�g2|�⨝�Z�ud����v�t�;�LW���3vNM	J��ZC;d�ǹ~�O[8�Wm�CN�n� ���n4>~�-QLs硅�	���3���N(`��=�G�ւ�\�v���i����e(�Z��CCUji����7�K�&{%�=a��;���Q�5��"�6��Ͷ���m�}r^
<��ڔ쮐e܋`~o&��_���m�{:S�P�x�#pג��`��\�
�a��0��R�-�FΜ���^����0ػOL���S������/G�2��d�A�V�x�ܹ�1u\T��oq�[W���(��5��OL yO{0[��� � ��%�(�f� b��#0���u���8�����҇���exT���c�x�`蓜1��� 
	�:\e�I��s�(ʞԜ����9r藐����ǰ�P��s�_3���mՂ*�r��Y̚�|w��qY%��P�$�@�ev���Q{� �@���8URM�g�<!�"� t�)�BH����Xo�2��#�r��p訍�O�c��H�{;�R���'�ak���¹\J����EX��0;O����3У�4�p�>y�{�~ �+x����{P�i�	-�q�#`�}�5���2/d^,!y7D��V_�`�'��<K�I1@�O˫HU�{�J�$J5Ħv0�hJc=dm��]۷�Q���\�8ȓS�ƽr�a_����#q`X���:[=UWaɱ1�xƎ��P�Zp��n�4�8��~�Mph��Y�T�Sa��4��럃�^�Y9'2�&L�+�zQ�D�������X�xq�c�l��9�i8�� ���f�pug��J�hi�Y)��5<��hA�뎤=����� �Tƨ�_fiʓ$ɝ����h|���߁�2�d�Z�����R��r;fҋ����?��ꢴdC=�rz٭ٰ탮d1��*�v����)8X�(h�u�X���@�.��V^C �gxR�xwi���e�Y�ьG�>��x~R��I�����]�D� ��^�k����y�u[+ �؟��ty־[��@�����9ֶ&`�6�H`��{k�d^o��aKT����*�38o.r�u�0QpN$�x;����s�;��y�Ҧj0J��N����*Q������z]R�h^�������ݪ�љ&o{x*:^aQ�&X��%6�X3�l�-�n� �=��'3�x�����E�۰����e�+0���α���7�$�DSn����-:�׉{�cz����+�%��d����e!%{�����Pq���N�K=���|,{�L����)���;N%6O�#��Ri����G\Z.�� i7������S'x+���u3"C�č�j�*Z�A��`�8�\XJ߇.����x284�M?T_bb���Sp^�O����C; �d4�Pf�DN�����j�0SF������^Q����Qp��>˿{�*Ӳ��/tj�iS|e���Q<�0�$���q��	ɘ�^��F4�s��U��͟l����8�u��~�#��-�6�]zj���އ�L�~�-�i�ǀ7���ú	�Pk��w���	�W�˧��R�C9L%W���y���W�J��vEUBy� ���H�1{�h`��2+6GJ��N"AR�$\�1X7�T�z��^j��@S����w���q<v������0���s{�>��b�^�y����vb�S�r�}ē�O��ᴯ�?n�;�[������H�Z��aD�r](?�<RN����x���])� ��F���&�ŉ~kT�9��O��5��
�#H�"@֖��J�F%�`	��T�������L{Ųzw���1��,�d;��,�#I�N�2����A`���ٻ7=O�5�������W	6�͔u�'���g,_\�0P�#�=����%�IN�i�6��9ʓ���J�p�h,�/a����&#(걸��Sx�w���*�/��f�l/��L@MJ{-`����r�igrM��3�bT����(
O��#G����ڃU�(��7Ia��݅�;+�4�h�l���lN�U�y+#,�;���#>���|�m�����T6М.M�9�iN�1�t������%��}x�0�i6����z�'&c�����4����eGA�݇��RyE���Ь���6(uP������q	?�w�>�S���
�&G�2�����?�}�C����7C�8�.�%jO�[���u(��S�k �h�w
� �F��C%�r�1����'��Kt*G��X���3��a{�6�� xT�($�[�	���	��#�O��KC
t`�TP�x��,i�[��P�!	T�������8�;̵ %b<34�˱��e�����n�f���oh��;�{j̦b�H2���n̐3,Y�G�'W���E��ε�_��N�$�"@B�1�"3e��o�&��O����f��ر3P���}��� �Xh�l�6Y������Q�H��Q���'2��@j,j�憋�4	\�'��j�"#�(0%��Na`�{�9Z�����e����m�C�`��_)S7O���^�mki6�h�-��P�����H���Z�b�Ҝ޺B�4�������k/!��ܱ�m7�����Qh�!K�r� x��<kb?
�#Ħr�N>�i|�ǩ�'=��!��Z؍4�ַ/������u�����9���Ene�#D�-a̙ ���F�M%Dh�+�adBI��	�.U�B�)5E�X������QV��cѲ��p�ê�l��,g���J{/ݚ<���!{�m��x%���R	���2i��EG����;`����N�Ì	�%F��/�G?�H�>��w�L8u�^#7ЂT���\I�ᖜ���xS��C"i����/����|[g��,�Z�ԗ}��{�\_���%�6��k�7Fv�X�XR�����g5����U@ذ���V@b���K^>�#�}$���x�֙o���[֋1��V?�ܔ_M�ș�L�+�*Bu��`StB,!�@I��9��%C̥>"�3����%6�kY�� �N�H[�ǌx�I��n�#I]���Q�U�k���Uu�5��	��Q���F�c�s�CΥ�w
Ox�m2<1n�b#�uj/S����.1�T�!�����G�%;�Rt��؁������)L�	��8��o��S@�i Q&��� a2�2ϝ�=~!3*�vqw ����ZE��B�Z�yFvmԡ�@��2�\���9�u��R��.�tˆ�*8��ة |(A<����c�b1��(KOCV���d�5�u|���9���(�ڎ���g���֭$5b'�7g���\��OI0�8>�A�gH��6P��������3a�20h#Jz�F,[>����+�r�D��:D���%��y�gWM�b�gf��q�A���ŷ��b�L�ua��q*���N�@B��,��>l�y!Q�� ���=����%ȕƠCvX����`W�������0��M�
��X�kљcUїT�Ȣ޾�� �*	���g���������}̈Z�yd��j:��e#?��z:�+����&���!|K0��bxG�=<m�������# ����[��i\ӫ:&�b|��1���`N�z�?|�W�y&!Х�>\2�(*��_�'o���"geX9c�����g6xmh�m�6&�����=ɚ$�oEl�~GV����V���Wn;!i�w�:�hU���7��RhO0��`Fj�fkXa�����#!���)�Ua�PK �z� N�L�5t�Ϸ}�ԩ
Y��˫^Kr�g���<%�3$#�x����Yh�}�
�����r�_e^��C�˩B�s1�L<��7�f�b�ƅ�
���LI��A�P���6><�����!!�"��~;�BE)ϑ&����h���DߚѸN���ztt���V����Jd�Pf��U	����=7SA-p���1/��4���g�ʩ�B4S ����$mbf��́e�O~�/�::
"�e�b�x=�=� a�:�����2A���6�p`h�z��|1��b�� GL\v �
����'~�&M��5$4/�f�/
_��핵�VV���>��q����(h�0N���]⏋\�R�PWG����%�����#���d��U^��-fI���`��u���`��/۬�Y1n�_=���Hj��9� �/+�Q�w�?�u�=*i1vV�Rsu[�Q����Q~H�I]�'������D5�?#�XD̰xrJEmK���%j[_�qL.���|�ׂ��q(g��+����a�3�jބG�. V]X;�C����530m�KJ�QHY�4m�j��b�<�{�{���Җya�W��U���˙�c#�Z쎪T����]��R�~�H���rp�f�/���T��-��+-D���\RRV2�����`�p�x6�=�r�����߻���K�ֹ^��.��I�����X�&���o @�_Q�T��z_��z�nR2/��L����L��>�����*�`�Xm@�N4Zr���J.h��S�t�SM�~�7R{\Xm�8��<ӿ��Y��Ĥ�rs���'����#DG.1�Hs��c��q�17�3�~
2ؽC�X�}�.q�ZZ�O��3[��">d�v��#QRNB߫���%�W:=A��'�Ml�N*���Ō�Ge"t,���u
��=B7A#�=B
6�a�:P�uL� g�=A����� sl�i���5��8��I(C�~1�|�Ƞ�ʐ��� =	r�FD9��b޵nK�V��ʒB����b�\�+�� 
	T�{O;�V�VI��9dB=�L����'��6sU7�^qo���P��:'����K^7��8�{�/�y�s���d�;n?��c�#RKW��z%�L�*����@�Gx�j}�SR�l��@S�!��n��ZZ�Yq��Ӣ�Nv� �c�w�k������ML�f��|�0���xe��g�i!Ŷ��� ����<�@��˕d:�i���m�(�<���cB:���J����Q�T

sn�!,9���3�zz��'�Ł]�%����i
a��J��Ы\N�6�N �/�C�a���6H=��KH#g1�H���C����C��B�1�ۈ��WrlA���[��)�Nn�a�����q9˙��Vj�����ԇ�x��]�*�eL�1��D%��4'�3mY�Tw7�B�?��C�y�ƒ�w���E�&<Ii�Y�MT�	�S�E�;*]m�H� b:rj�:�|��Z)�0�F3Jj��p��f�&D=ڤ_�,�	���-��ڔ�2���.|����xf�uL��/aNP~T�kz���@��-�F�F�Xl�si�>�/E3MĈh�þ�e|C��	�}�
r����(!X˰J�Y���X�0�F��wf�M���-,p���"��T��E�BgDg�-%A��r^WI=ue�"�� ��3�jt����̈���|�8��q�j�$��na�Zjwݡ`�m��W����@�$Zhp�b�:�}⮆HA�5]^ET�qUw~������8Z9g�%t�~T�$�e-�vs&͸:����E}��ʁ(w�fIIt�4�%�n7�$w�u��}��r��(꨿����.�����[�	��7x?�t6ᮻ&.)��^<(udҬ�7�CB���(p�	@p����w�f`DQra���lI��~_!�F�L_g���AW+�s�gNq=��֍���+yyB}/��F
PWv3����+
�gI_�s��`�i�������nI�%މ㞕�*��l��F˴��EJ=�Wtݗ��(�񰒛����<��w�W}��'U�g����[�	����������Y ���VEY-��O̗����4�p�aR�N�܌|ʕ�3�z�����Q-��}�`�S��3�$?�����u�s�(��϶�9bs��� �:�6�%��>쐆�ac�*:;r6Ϸ�����	0�#~���,R(��:�롅P�Л�^G(,t%�䋁6����e�+Ѽʇ�2���
7�">+��`�}a�+l͡'����' u��f�榮 b<@��K	��J��,�&ITT�bk�3�>��Z�FT3ݷ]��H̅׬�$��5IU,z��,�K��fI��P?�ćҊ�D����֜ ��O?$�i_�Zú i�-)��D�����?o�=�;u�.Gs�������?}�"��i�#sAB�[Ғ�5���S(���l�8bd*��`��x�] 
�w�i�p��h��N�����${���=��c��ە�MS��`���H�U��2�rAi����d'�q�o�ן�|je��	���y�
����@���B�;%W��{��l��f���$�'��G�oq'V�B�gW���2N_$�C_ف���N��|i��!�<Pz:(9C�e����"}����s�A/�"��&��g����h�^�=U��G����8|�W2���c�e,�Pz'x�b���:�]_��~���i�/����]�Rk=�:><xC�`��s�f��tU$��㣹�j*ܾ�0h''k��N�����(0g�ƅEC�ӕ7���B�:�����f�ߌb�/�:7�3饭p��)_%yY	w���+B�G��c,�y#��T�L�h321�a�A�XQ��m�
��1iW� r,����N���͉`��4�(/����p�1��(Z�����C5K��0j];-�NĂ���R����&'��5�N��E����|q)�=��zݪ�����9&	!�pYrF0����F�g�,F0r2��}��F�~�2�C!����HN,�87�CӾ#���*Q��Su���*�E'��*�A�ȻZA����<��2��=�l��8�d�T���I<���\���fP���R����u�#@y]��7:��/��J>[Z`E�qcb"m�U��~�����r��^�OLK����~jVvD!V�]���$DL�
�Hn?�T����q�|�������),���)��
[�T�>\M'�h�cW��f{ӰًM�d$���!n�m�R����(�P�O��!emSHۃ{{��o�YU SI��"��/��X "�N:�r0
D���S�b�*��A��cޑR�4ณ����m�tB΁�����=�t:�5ٔ�E(���XE��&7[�T���*׃u�)�´�W��7���؀ˮ&��H�(�,�Յ�߆�h��$��L �h�� C4��]�A���,H�;f)�V�EH'��6ih*Y{X�m�=G#���'e��n7A������@�M���5h��O��Ub@�u;W4�F�CS��X��'�v�
�|��˘+�z �|ҹG�:�.�/̴G[hH�����8]�d�0g��q qh59墒wfL�iǺP�e��|}���c�9LS��p�W�t?�D�C&�a��P��\���:OJ$=fj���|����2�$�} �]C�o�B#�]�8���2��:��ڣZ�b՝�Mtqx-8��l+,�C`�6C)���{�&��gC�j�1���_ct�q�AC����- �����~^�?_Zs��)��O/�4�}NTk-�9&K����t�ԪM��0���|0��Y��)D�+胕W�(2�'�����T�P]~�b��^F�+K��
�=`\/����J^��U	���Q�	�N,���nQ��p�]e��a�0?eǓJ���k�?}`,�8ħ*��� ����C�`~�������[ !�.lH]k�n�M�0�V�.j��`@�b�2�Y�Tc({�`�����8�8p���B�T|Gd.A�'֖�L��PR����[�/`�0��G� ,���$%��@����*��1&��w���N�S1Ax�l-��b�iΡ��=csI%W�Ȟ�L}Ӱ�f�:Ȉ�]&���W0#�-?��?�����CC�7i���2��G�2��Wl-ͩ�΃��	�n&�k�9�/��|_(�=_+I�C������N�/0X=�&�	���&�2��f�oކ�b}��mV��nwॐO<���%F�{H���r����^W"��RtNU�����c���3բ��_���1ϕˣ}��kC���!Ьe�d+��C30�'�<P�ލ�D���Z�^�OO��Ot���� ���P3ٍ�	��т��4K7z���:7�����	��H��/��2r�9OR�[�z㑃ˇ{�*���P�4ђ��:��R{��\,�XۢO�"7�>c��Yਬ� ����+"-�!J"�\L�&����@+����F�@���*�^�2Y1"u��Bޅ&;ko����@Vx:�1g�+u(���P��1�n!�Ez�z��xy�O����D��dÞF��i1�����BڄK?�I�d�dį��gd\��B�#.j�C.��� ��Z��{��=��~��OBdPfY��?μ��G�=,W�	_��p���%|��<rs}�ch-{���������O*~��aGrٽ�4mF��pU�%EqXN��V��d���'\ω��VQKM�D��Nx:&��X��~�1��l��ac��]��Ȏ{5Wq�p���,'8�M��+�+�4�e�-eOz�Q%a��_��b��2
滼�e�QXsX}4�����vQ�x��v�ۓ9qs̮S|y�`=x;���/�K�*���2#H����5�e���cf���Q��~p%��(��#�~��'�z��R/#����4���#!�۷D��+��''n	��A��^0�R��D�2��򡴂Db	�F�'�?x���d,Fk�Y����_7y n)��eC���N��ߝY�kX*v�&uT�Ԣ O�Ȋ)�U���k*h���^�.��Ejs�VU˪a99����4Ϸ��A�x�Rg\O#��@�t�6ԧ{Cn<�u���0�o�$lH�m8�0�xIK�N+#�
�bή�z
�]X�T��9ك�d?t���e� �Qxt�wNP�8���GY��P����S�G4����� &��tG�5��0�mӧdE�^ox���,�?�l�_�=�xTn!�(#J���J0?��߻���C�X��9gZ��'}nb�e�N!�ޯ`�s�x���F!��ߩٖ�2I<�J9؁G�>�+&7�a�yi�2���hnz-yb�������i���t8X�@Mh�«ǉXs ��sE�[!��?�7��V2Sg;nT�����i�1����@Ѽ��aT�G��ţl�<���B�[�u��d�ᧂ�]��l�o�jG�����9=Ws�L�t�v)a#�^�X���_�=�j��6�1Q�}�۩ѝ�/Ohii�q�CA!;��&�7�_ϙ$S�x~3N�M�;o7Nd+ۥ�(a�FC�����CƌP������{:���x�!��V1�����J(~�˿�l#٤{G�Z�ǳp޻�
�]��p	�( ĉrO��<��nj�����Z4�H�١�^Ő)$z[�O��.̮���]�v
3iXQu�G�Q����`�t!��nm,`T�.H���D��.޾7��((���M��uX����]�:K�g
���������R���?Y������D����#����[.=�u��pt����Y����{�ZMf�YC9!�Jh���ā`��7Ȃh��6@C^�G�J:0��z0��|��&�tT�)�_�צ�#OB�8�j�8U�k� ҕ�Ɯ�8�>K�������_�hR���C��b)CYخ�Ly�kc���i��?����]��Jb�FD�����M�5�� �b�J8���}�E�2� ��F��%(l�喛�/G;O����E2
����٫N��� =M^�2��#H�|�T7����sd�[����b����N��,�:HKW��G�lVX]���ُ'F�cl2XA�T����L�ں�xH�*�K�gM��LH1���t�zT
C���p��'��c8�F���n�WZ�MW-m(�\�DP�m�U߽ �������[�������k^D9��`
�290��CRK��rs�I�|<�n�۲��뇄e�+	�ř^��/Nm.fUA���0B���@Or �����*�dh��U凅�@��Zz:�>��HV�Bхg�Q�kAc]^3��+�>7FU-,1#���1����P��n�_֫$d�3pNi����(X��6��t�1j3�saE��*>Q��ݨo!W�sM��S�"T������b��]��J�_��Uѡ(s8ԇk��q�u�.K0O"����5 
N���k��џr+y+����*�o2�BH�^wt����j�:*�>L}$h��
h�����}���D������ݫ.&X��"yZ{��-�?C�[�ޔ�Tj����a�w�T����:�}�|��@��	�ɻ��:oP�AZ��mx=]L�Q�ǂL		����2�U� ��T���S�:w�Fjy`��ܨ�,bB6�g0��v�n������@_o(�l�2�r}"�`�Yo�ƫt��%8���uBr�#F�����x:#�T� �/�vE���Z�B���Gi-ȭ`X��;]���~ۜ��^5n|�I��a���1&�*G���٢���jE�mS��X���:jF4��$ӥT<�%��h�#���x,�J��L�F�궊֏�sU�-�����t:2�W��I����X}ӟ�oQ�[B����ڂ,Дȡ�ۘ\��.Z��<XC�_9�k#&}���]Q��*�|��Y&����&�����%�Z>��]��U�C�s]��SY˺(�H:�=��N/j<��1.e�Wgl�㲵�x��B�qR�h���+�^1,ɻy���-�B�������h�`�cm��w$R�7���s�0΀�=��d�����7]�g0�]ćL��Ӡ���\Z�>��\�w���2����E��Q���׏3a7�@�PhP���/�WD�@�{�K�V8y(��AǦ?��8OD���ww�"��c⍬@�S���	�� �qJύO���� ]��揢z%������4�}K=����)�W|Ől 0�)<�.AH�jw�D,ug���2m^�1��'�k�~R��q���F4.������z�ST���Ì�Ȍ͝w�z��y��/�:&��F*Ƴ�c~��^��?]�i:d��"a�%�n�	04mª�2���Ԅ�WGs[�M3���Y�w)i^����@!��J���Z�o����RG<,����I �i:�CxXB�^��s���h9�0#�ʂ�Y�¥p�R��<�(FS�3���~k�BH�GĤې�I��0����ت��W�|��"�6Yo��tZ&rĕh�;�6i:":+��a��kW�z$���W�d�v����2��-�o��+<��$W�4�W9��Yt�#�7�%�����	X8�<�|}���8�|�b�K4%X
|;�t̻F���j32L��W��态����X)��X�)��*.Db=&#��4"��̚���y7� ͌�
��������RE������ӵVӍ�ͨ_nǍ�����k)(3�7Nقׇ�5P��<�4��ڭ���_R'�TIq�󙒘��lc��R���K	Sj-K�o��cc�o{P*�Y�N�ĤBXˌ��8��{�`ZEȠ�� �u�>H��L�g��0����33�A2�~2��|���r<���g���x�ڑQ�
t���~��-ͪ�8�Ew��ފ���û����{'{o�s��Ń���;�5wH�� �/�.��¬&Ĺ��߹j���
��@�^�+��L4��+��Y����p�B>��J��^�K+$��1&q��2/^rm��B��k�Td���7��9n���u]ƨ!������ʨsD��-}�k8x�������8��%��D��F���N��q'�|d��"�'_�H7�����`}����˦��Zﭾi{��u�|�Y�;��lm��e���dG����R�~��1=�����w�)dpxg�1�.[�٢#�u	��gH���N�<zzVNcVt&�Z�},K�Z����B��+��|�!bI�ޛWhޭq8L���WBK�lihڜl��~K���j"kM@�@�PVn��� A|:��KXD����������E�V2�}q@�Ur���c��V��?��V�S�n�\�7R����W����ٴ�1����R8�.Z.H*je��4��X�w�����Q���v��E5;�xn�Hq{�̿�,�cQ�ñ��q�l�d�����gL
F}�AϢ������i�p?\/"o������T��	��Ţ��B�P���R�Cن��� ����d�$x��,AZ�s�Z������L��;�֬�=��n��_D�6Y��i7[�T������j�g�ĖW"�pp:��Q�}��$y�ޙu<������I� ��&w����Z�k�}�#��o>!EZ�L�{{��.w�j����؁��N�pN�W[?X{g��'�H�!ﰌ�U��㬨�ed'@��F���x����u1@_j��Y�/u�o3��iKy�u��ðU+�_��&O�����߃���!:�w�M^T@>]$��̦۱+��\��B�jg��Vt�L�)�{T��X�Ku�vkl7f�?@@y>� ko�\̓�
������6�]�����|��0Rmy��nd�k�,Ӽy �}¬=z�T��rA�9:��܇2�N=�k����I���)�0)��u�E�D�,�(�0�,�[��_�����X�oJF��M�d�<�'�B�~L����ۯ]���e����,x�dJ�.Ol�kn�
�Uِm���[�i3� ���B�5K)���K���'|;�=���՘�S2���+s��xO����LI����Zi�4����<tbR��L���+<�$�^adZ�GH���_,t��`E-jQ��7:�#F�)]������k�훼���0�o�.5�\������]
�����&�jo�1NL��/�s�[�v��1�wAL�f���{�����Las�<���^�TM�!*�?'Y=���2
�'8=���l�����z��q<u���պ��+s?3�8A�Ư����~G�@���������ۡWe�nb���$Rq���yV(��T�c��_���!<�ʸ�chQ)5����q�T�]���k�W�̨ E�@���E�p��~}P��AuY ��%�_d���AO����}�d�kWlF�����	�o��ǒ��r�ڈ'����AN���]��x�x�)Wq\-��B���'�ѯN�KӟV�BY����J�O�5�/x:ǡ*������54#��'�B�	e�EvB��p)=Բ��fΣ��b��h��HZ!ệ��A �tp��1�b
9����v�ɡF����Wd߆�a%�N#��#�t�Ũ�nD�e�� ��eљ��*YԞ6?��?��+ϕ~�xS��ƣЩ[�#�Q�S	��z�W��ʌ<F��A��A=�8�x�I���Ԕ��h`+«(ߊq;S��L�x���4�� ���,�_( 3I��e�=�v��#+k��j|O�	�4���#'5ђpA�	�{�q.<����'�欿�J?������/;h��{�#���i�nDn���% �8�-�]��-�<'Z*R��t�O1;�^rP��@%}g@�38�R_��ց���>+el��-�h���%#~��ؘ�I�z��D(��+��<n~���>�f�yЎ��CG����n���v���_E�ե����~ ��OW �>����U#	;&�`f̝i��DQ�V$��V����s�˵��%�h<#�Mz>z�y�>e��㊆��E��HN)'6�d�~i���V�	'+X�5Bq��b����'5��9W���jI!�J������mV�b���c��>R���(�r�b�|	`$5���b����Be�jiڈˤ%����4b4f:2��A.N���X�x�6��L���x������7W�T���R�- �<T7�����a*;)3���Ǆ��d���ƚ��y��8�:�T[L��H:d�5���0�KU�qC*I<�IY%�r	�i����Q^�B�\b�C���"���~�!��^a�jw&~��a�-$�g��Dy���?DZ�.*��X������C��꟏�귽��q���NH���o�e�7��;h� ؾ���i��Z��E��kbM)Z�U�~ٗ`�[C���$�����pj�<njH*�e
��n���9�2��'Qޫ��x�>�����r��7bIx���:�f?�my�ƴ�[;,�f"5R�"��c��T�O�l�����Z}��r���v���:�ΐ7PQ��?aK��5?��g�T�>�J��P(մ�Ȏ�ga#s�����E�;��+� ���P��$�.!��!��"z<�7���33�w/��R@��l����2�&zu��ے9���;�wT�20����R�t6� ����&�������_E�x�#s6�Yv�Z-t3u�0�ee�����	�t�o[���}s�׵cS��^d�$-,݅5$��{�ܖ�-V18C9k�8.��z�ͤM���{[b�k;~j�\�?��՟�L�	�w0|Y��0��/3bS��Zj֝^��H[MUϹ9��M~������4^�4ֽ�Y���w�k�Cv�N_�V Fj��u�:,`+�8s7Q�"dC�[3�-��v�ǳ�8��������v�ͦ�����mj�5���s�o݀��q�򣩯-�ms,�Jt�CUs����y���ZU���3J�`K����@��b�uG�A��i1�|�o�@Rl+m�?�|�aVW���R����>�H��'\�� �VA7����@0���Fu��M0�����0���&�/Ny��ί)3?--G�ΧHq��9�4P�1'�@�ˍVs�-���9x�K~���^	�˵� L��<A5lc7��$�oyW¦&8ҟF�"[���n�6a�y��^����]`@j/��*;��NѠ��tY�o#�N+�
e*��%_�~����H�wL��^������nl�!�BqG����6���P��=wHnD2`���؏QM��y���3ҭ�il�v�N�ҹ�����ڿ������Y��Ɠ��Zg库G徖Yݹ�6W�1omQ�����!@�?�;E���g2��c*�A"oB?�a�x%�{�+�!9Vr21�D��W,�-���Jn@/Ϡ���}$ވy!EM��a���g�+0`�E������`B��t��?���G&ZV�h�����V�:�/��6��r(:G�KѤ�Q�f̺*�y1t��h�cN�R����'�F�{�a�]U�kG5x��3��,?!S�?�Be>�ܛ�/mT��b~tR�4�<���I8K�>�k���&�+)%�X�
�%���f(;ֈC�Jǯ���˺�\��T�hZ��<<�(`<�Ns�֐���6�����P���W�u?s٘�sc�N?�^�����t��Q�xօ��w�/�$ ��ԁ҉$]�JW֥s��$��ϟ�},s�w>Lm�������қ@�=����A�=%�p��{oBf��e�m��Я)�e�X��v&�Dz�SݵW@ሞ�
� � �F&Gc���w�J[`�?6uEݨH;��*:I6Gy�K�)#�#L�m�.;ݥ��=�U1	�Pf\�1�r���43iWu��w) �\[����W���G-g+.?E]��G#�0��N�7x9�TZ��TP�i�܆�2s�Ll�T�K`�/H��l/����+(�Q8c;�e��,P�K�1h�#�\�6	�-Al���+�!wg79��w_�J��C)����>�݀	��i�¼r��*�Y$�5�ٓyY��W�/�SJ�1�������$"̰�.��N��@#��]���,����YO6�!=<zy��0oNJ��� �Qʢ��r-re��Q�ô����|�'qtǠ�8�j���7m�P�tZ�� p����
��B$�Mh~��"Ϣ:��m�ׄ��H�!��
ib�)��P"�'G.�zz���u)�KO:���{��P�-����T�jR3���f���D�X�c�*���@����p��Ӯ���#��C���i=��nx�Ab��$֔L�)��k��(Bܴ>�@P:�$_(�E��h���p?��������LA�TT��t -u<~����Uѡ�i}�®>�\B�A⹳]ʒ�C���z�����jb���B��Ĺ��i*�3�v���<��Z��v\!�]�A��ll�U!���8^^��u��(�	��BO�{^����n?��3�·���>6fC,�m�y���Yņ�sph|�g[�?�y�cc^������ļ}�x���!q�2�bo�p�3^�ŧ侅
�@[�����}�bh�9ܓ�~���������Qbd����l7^O��BU��>�������q�Rg�(ܘ�(y9�mQQ���3d�z��Y�N�n���>NZ�"Y��U�t"vxEZAҧ瞉a��?��2םU�Rk�?TĪ?��ꩡ������CF�ߔ�מ!��7�+�'ѥ44�s����Б�m@��R�����&�<�9I�ޢEF�Ḇ;fNE����vQ���S��G��|o�����\*���E��V����۵p8iY	۰��F����Y�����P�,�Bt�ˬ�r�+Ἰ�AO��]2w�v�< |u=�Hg�iH�߈�<��t,���,�)2Ln(�ܰ�<�����O	�`�j�~1Q ֕���^�"��V�W�3��	��?b����L���Y[����D�s�������	���j�$�����6`\�np�}�6�.��H��M�n�Aq{�g̐"2g�ā�����
���m�7Z��u���F�	������pK�*Hh��T�5F��ˎf1�׶[��Ŀ��Z����1��]��3Q/�΂XF*��֨r<�m��83��1�y{�����]�K��@-�6�.��8E7�� ���#wV�)j_H�_��dX">����$^��_�4�k���x�vİ͓��u3s�q�q��&J�8�`��z��܁�L��ܻo7��.zU��n苅��c���aUQ.�#ޱ��?��:�Z�>�ř�1���`�DM�w��yw�ov����zE#¦�8��\�Z%��*͍�������S8$�ˈ�M�:��Y�FS���oڪw�D�be�h��2.�pTP����_�$�	�K)s-�R���(�:2fC�^�ހ���3�SE�����L�+{�&6*+���ڈ��iv�F4�kw=�����L���X���W�H�Fq�]m�:��7��ą���$�t����{Kz�tS�kF��вt������T/�s�n#f>�(�C�.�orr�*�WWbP���o��X��Eذ��I1��H��g�S����ډI9���<4Nz>��'�N��Ĺ��7V��$��K��{u^&��M�&��x���g��*���Dn�́5O�h�����v����f�ݖ��I���\i�p ��[�jV��ᰊ�H��"��&,�̳-(��s�8���ƅc,������-�3�6�\�c␾(�q��}����b�$��s%�x����ST��g�?��k�\H���}�W���Vt��� /[7ܝ��J�l��R�Ĉ�{�N�i�G����X`������aa�q ��8  �?�1�Q:֧r�!�%�S���)����h�vB�P�m��w�h���I���K2BZ*[$1���]�{�Cr"Z�8z(��P>��3��m���k��a����OT@VAA׬�U���&�f�� �����֜>,���x��-e`%݉��3ɣ�_�g=�99&�4���k�0W�M!�SX(���[+������Kԇ)���h�ώQ���Ӡ��xI=eM�#��v�{���k~:�K�
�}��xf����@5�̏����ء+�6��\D5P����Ips����s����?{��Y�,lLةd@1s��M����P#�D��rXp���:g��Uz���W�>�$I�U?[�����ۻ���k� �j$U��y�,�"d�e�:�4���]��nNN���^K�v�99�:��,��_8Ǉ�r��V"��
���/��2���^�7�6|)hlbN>>�mK��� ���y��Ir��ܟՑn��K�΋wzZ�69�z]���^H�Α�{��斕�wv/ӛ�k��Gl�Θ.����E\�Xĺ���{�KS.�k���&�4�!'��@�[�����eK�'��
�D08�����*��9����Y�P\j�^�ǁ6f6��z`�lP*�#�bEp����x����Sz
�uI}x縷��S$\u�1R���]�������Y�H0/�(��Q:�\�sc]�����٥I.�Hߎe���A[C�Gvh��T:���<���n�
jL �'b��`�a0{�,��A�m+�����%��ſ� Df���K���x}p�'�t�����	�v�a�o����x��x�$�I�:MeK���Ԓ��|��p?�n���c+U��؛���
aLU�����8�Õכ>�o(TPY���=Yd��3�q)��!�Y웻�hBM]ӉV����U�o��1Y��h���W�gY�i�]�g�Ϯݧ�v���r�#�X��Qk,��V��7T�����Ҝ���K+��K�c1֨���7�l���}��*�$��I����[��5b���5m~���ܿ3M�Ps_iE�DUm*�,�J׫���D1��T�g�P���!y�d �!hD!���=:=��(�0��1�?���U��hE��ŗ���o���U����$���Z^J�'�����uZ�o�}�[5�z���oBy)��W4�������H ` �����̤yD�P�3B|{�
h��?�ݐ�pgp�W��w�6��D���'�[�X�3Jҡ2��ζ[�t�M��p��%rXmt�Z_?�w:�7�u����ʈ�r���٢��0L�oz��F�Hn��t1Q ��d2va��� �	�b�_�s�=2������aZ`]V�R�p�a�-(������I���=�T1첒��q�S�ģ��.5�{�p�85���w���O�uD��Y��/@,=olr�j�zc:R0+}E�t�WƳQ�P�%���Wc��ш$���s�Щ�ǭȼJK���������i-.r��9h������֬.����*���on�"��[[7�����4�j���}Πޮ�� �-��U�%x���2�r,�fB����A �F��vY�X�j��E6���Si�]�4H��W�<7P���]��3Y����p�wI�ƓƗB ~
SyE�}�~�yJ��P�_���`�����K$喃��g�כ���/�;׬.Y��!�m2�Ɩp�sP���_H��;����}�cϳ�/]X��L���םd+�,�5a�%�o�t(6��/�B�V���M����#H�бBJ �4[��I�_VL-�j6Q�ҝV�Q�V?��C�[LBQ�R�`ẢPjPh)%y~��*mi'2�	�	N�1�"w�z��gE����妜̯j?�]n��R�V�T�봍(x��" �М�-0�"1�^�݊5a�9���RV��M4vˋ+�zhT�6!�{�mJ�h�B�l��#�b�V�J�2q�tN7 p'N��q��uw��?s�ڪl��Hn=�@)��9e�"��XJ'4fv]J�w��U�y��X-q��RDoŉz2�NzF�/���i���\�4��z'��|���H	��I����I��t��j%����X�����a5��k#�܃�찴#�O�������*�h��� [e�C���>�t5�LX�r-����`�=���>mn7��5���p=;S3�s�]��)������7ǖ�%���?���[�h. �DDa\{AQt��������5[�v��(�\(JPR~�Z�.�J�	�v���;:E��ǅ�t���;r���&y`��.��Ѳ�<����w \<�� ##����h�RD�h�^�LN�&��[�@��$�9�[�.tA�e�F么U9o�{I�(���A�XR|��]�����U���T�t��d-��_/�T a05?E�����r5,�{��u��Cl�竺��M�PQ����[t�� �'�'_��8�
���ì��5�,� ��������(2�("J��b�-�I�x>�
�x����$~�E����A*Z��<�����K/ym�n:����ٚ��'ٔ�4ZQ�ؗ>����a��L�)$j����7TeL�?y �)F&��h)0�w��Ej0�\�>�9Q���̡���Hr�0%Ǡ�t�~�ɶ������jM1�ҭ�������;C?z���Y�-�����D"�V�������:�DV;ν���$DXx�x�b^�O�S
&�bޓ��Vㆾݕ�s�{N%��b��Btc���~R\����t���z2̟b~�3g��~,N��x�P�����3g�
隙��m:1�]߭=�Lm��{�����9��8���%�s8ՠj��9����@LF�)�ǉ�\A"�"L3;ϒ5u���+�v���cuziIAwΉ������E�!
L�<g��>b1R��'���zt-��C���Cd����
���i }l� Q�F���'jt�(���S��ID�B��`�5��-�<E��P_�W�.Z5U�3���T��*�Q�߀��&N�7��>�!�Y)��RҰw�-7�"Yx���c��AqW/]|(C�R/\��3§��Qy|<;qNS%�S�f�;2Rkڠ�*�K��Ћ;�uf���,�I�|�J���ĺБ�t#����|5El~ޑ�l�zw��kMY�%	�Aqtr��eKڰ-*_��	�/&��(��
a��� ʞf�i����t���m��]�5]�[�J4�1-�G0�[%Z���jߧV�
?�m����lC[��1x����B�q��<vD��2d{;U�?��>�l��|���_E~c�w픯�A� �RR��0�0�~�7b,���ϥ���b ��G���]���I�_��?q!���,[�?(��ݨč��h�3�QQ"d�������fA��aP�+�A|?��uyy��]�k�:���#�ƞ)��$�P������Vv6��V��Z<A��u�T�����TT�(:�K1����}���Z��:�*�u��4����r�0~�<�ߢ�Ў�/� �\�I��a�}g�π�x�JY�����:l�n~~pPIg	^��;?g�q�yw��>��* @�[��:$G�tΙR�G�v�w#�Z�S#~E�o۝m*�I���ج䋸���
{�0��9	-������"C�8X������'�ړ��k_��@32�fmv�(A�KY	�td�۳�F��ʌ� �V��'_ޗ�DA���uR��lǾC+fC�\���LK��#��n-�v
��3���/���u~pP�N�������q��]�ϝ���ǋ()�F�����Z���Dv���v�E淋�����+�.�o�s��D07�i�<�����Դ<��u��An,��fSh���B�@D ^[ҝ���r�k!�i��(3Og��;Ol<��;Q�iQ�M:$t�Jr�;�U�J�z�Uэ���ȉ��8����c�(�+�[���6QPH,tߑ;���ʪOr	ω��,Q�_��x���+8��T736�E��,,�0��vL%[WP�L�>\�]Ѕ���2׿��R�K�� E�ns��a�NN�Q��1���)����|6L��*�}�x�5*�^Ꝗ�Fl��*��,[{!�H���B��N"�S��������wT��0L�Y�b*�p~6GF�Y�eԽ5�2[���lG{p�lW8�����Eǒ�@���.�g3��B��p���7�?+3�/,��f���z�}��?��C�ňQH�Av���`ﻘW�tf�-Y�O�������k�T���G�����d��F;�w���tЫ8�VB�˷�hō���81�P��VoQtr�a����>D�����m���w��������:��d�rE�N��;���^9u^�)[B5#'��f�o�͞��Uɣ�p��^���W�$}���n�٠E�d͒���y�jZ['��B���l���"�O�X��!h��������S�u,J����1��#��D�U��vi$�I,�!H[�gT������J�sQ��lE ���Ω�z�O�T��	7�pJ��H�U@)l5�����l��,ЉUr�}�v(4��C+F�$߱�������m�0u�_�ac2C�?�����[1$�!k��O������?@�Oi�E�����
h��ֽ���I�P�9�r)wN��д��I:ۆ�T�"?�W�X����oJ�~����k	Cě�>�W����#_�� K:�F}&�R���=��xW�p�U�(>�q�Q��١i�\~\�d��;?1�����<��KI���Xǁ�7<�o�Y��w��.��6G	@�q�,ǲ2m{� �ɢ^W�8��e�G���@���	V�?i�\��"��;���S����Ijt�OiK�O-B{㪞G�n7T��ڸS�IQU��d��e5�]�~rd�;����K��s`�����.�M3aaa�^j�q7�RF����t��
���x˿ۇ����C��-h����\
��r��# � .��ԟ��0�aտQ�T��)D=E|��b�����ף�cg���W]s�d�V��p� �Z��{^��k5,��Yx��˵�S(|kI5�u�m���?��(2�������Bx�j��/�4�3x�l!DhZ�4~h��3BN�8��{Q��խ����i�:�L����1v��jM�c"�~h�"���R��]� my6vi;�6�_7+���l	0&R���]�ߡs ���+��+������~�ju-y�>������Q'~}P��譔Z?C��:]���4A
>(��T�+�L���~�r�V����-���2�� .�=:oH�K� -��Q��>�=�u��)��Y�XH�q�==��w���q\�w�5���3pOO�n�;�	< e?��w-�[r[����"m��� A{�(�=�2� ������K���h��%faTK�@�O��gL`��(��X=�����j �.���r��4�Ks��W�����'^�D�*���T��N�p�qv�5��z��Yg��d�"�R <Y?�H���O_�� "]B���/���/���W�vM�a��a�����7�k���1<E�Pv}g؊n��ˇ�W��~�<�E���%���C��-Y�+��Z?h �sW���	���Ό�����S��e>Q���(,N��nmT^�:��������n��XK�Fc�������-�u�V�a&�ȴ���<�A��!����AhY�7שd`}� ��T����)rBo�/lyhȀH��VI�!T,E�&)�y�����VV���mCHAz��@��6�����1q����n_��&��J��(+��ǖ� E�u�Y 7�e��q<��ә�����"���j���G񒹻!V�����LPYe���2��?��3=R�a�=�G�� (Vk�N�qTx������D[��g����_���M�<��G�a�	'2����L��Zg��vll�W՜���1}W9[����z�L�iӉlДSW4����_���hߺ{8�W������{��X�<�*��T�4�/�_���"5<����.�j֬kuAs|�4h��:��G����_N� �n�#�D0ml�u�Гs̘lrԤ�R+b�@��Г���ف�l.���w%K�,P�Ø����/t�O���h�:�s�9H�Ck�ٙ�e}8yP�C��5�ё�jf��E���U��o�)��<��ϖ(���Ey#Q�x�d�	�P���� �,�N11;D��yQ����w=�\ؿ�-sO���S����o��x$�mVҴ\��@���
�#�)VRG����W#�*88���?��X"|U���֦R�M�B
2?�w�������TX�g6�I�AB���V;� )s\���*}5�(�y�ᤃs@�H�tՎl��4Ϫ�#
9e�;bGZ��������]1�[3�J����g�\��D8m%�,��ҶU.D�����ZXh����(=�Z?W��(�H�=�_&@�����/�ɡ�y�Ao�b<|E/O_e��;#֒��%ʘ% %+v}����
]�6�`��)�0o|BR(�7}�zDG�樑��i�`c�uqx���Q��_p�P��jD�r���]���r֭ۀ�����a5� ��,���*�.J&��K�94�R�z�s�~��<�;�ρ�R����D��p��_-�~���9b8����s?�肁���y���`@��O�����'����xa�'��&R��㮈S&0w�9zw|^rQ�R����+���*U[(`�|� _��Cƕn��2)��QԾ����F��w,�a�ϧV�c���+U��>/��N�/��H��͵&^�O#�; �vʼ������PQ> ���d�ษ�,�\0�#1j�O��^ES3�n{k�����;N�]2�0O]U��s�1ow�����4=���ApD��ﰱy����Q����H�V��z��,d����%�fm?j/�#�{C8ѧ�wE�#����$�S��ud�}��`���Q'"��3�Rj�G���iv�T�r	R���\���^ �ec��� 8�d�5��ed�Q���{��T�XMYg` �{�1���F��z�ޒ�& ��0}��:�B�b ?�4�<I>xf�Q�2ci��<�\��5O�x�������XZ�D?�����`�y�]ny�]ƽ6$Yw�Ԡ��\��A1��^J��m��f��M}~J��eK�8!:}&���&�dH��1&����[lX\�[���?2?��]�vƾУq�$����O�8��
�ow2[�ñZ��@�u\/�ԧGб�㈔� "��e?���o���"���y�w�H����� '��N�`�-���!�Z_�@T�R�]���iR������{���u:���� �VJ�O��87ֵ;��,&�m�f�������Tr����A���$a�������CZ���/Y1!b"__�K�"0��'P?0b<6�-k�v7q��D��1�7Udf3-�����j�I7�*sQi��%p�)��A�)�-�w�df����+��4��r�wY��{r^S�h;Zl�|�	A��RSQ���\�}�k̾7e-���,v�r,O�ݣ H�L/��ܬ)�A���Q��^��,ab���|�q���<����/M_٢�G��Է�!ę��j:��c��R��PtQdыaAE��L('4<7�H�4���IE��J��p)��7�F���Q���?�ۈ�;�tg� �֦��t̢��gʃ��Z�xz<��Z�Ǌ�;�W֞��OP�^�$��w������Z�Yc,,���r�u�4�$	%�w��o��o2�$3�Z�z6/��oi��ôJD�(äcm�x��P�����%/��a[��A�Ap����.�ޛ�؉����CN��{�Wi�>|��(a�U����d�W,U����d�t_zo�f42��D�[YhCbx��R�CO �B�|��T�3ľ$�ݭ$�n�8��ԁ߀�LF�s����^����/��2�!�/Z,��ă�p�`@j�&�q܍�(�ӎR�da�h��
rݨ��[�XyK!�$(Q�NGa��@U��X�;+ȟȱ]�8�7���D�WU�؝��(+�����.����+���[��WLẛ�{�-�pB.�ί�M0=)|RO�'�l8#��#�t~�MJ�8�u��*h%��ڍ2�:os��O��>�O)���ܥ�9���SRt��:�����`Aw-�������8�v]���M�Uw����z̯�v�5_��AA}ޙ�U�=�>\�L�f���!hy���Z�>�r�vV��Z�R�}����=u�!Y_7`��ahD��9� ^����9ga  �K��~������晶E菀X|N�Q)��0=���R���8#��4���ܿ�OgYB�L�����&����^�g��%�`'h_�d/v{t��Л���e ���֐����(p�e���4b��n���<��G'Ѯ�>��'F��MPi\�Q�K�q�C���])�]9��;��r���B�=���%Ү��r(H��d�3t=�?�rAūyp�ǂ�Q'�ֆG��}E��pW�s:&AיF�i�o>�]<ЎҢ-UU��d�ȶ��qW��Ժ�YN*����~�/�B޸�͓���^.Jp�ь��'c�&�8*���.�s23F��)�V��ڞ��:�yvD�<��VP�K��^0��e�l��R���s����ۻ�0���No4��G���/Pe8%G��ެ���A��!��.6b�`��ŷI���0����0�C�V���ۑ���8�-HJX���a�E[��}��e<g"D\yJ�s��l��{�f��өTF+�%�1����VLIS�;��>��y�a<� ����-�BcA)E�q�:m�˕��5��fH��D�|̟���yhB�r�{�?�p�v�8N�6�G,�"�j���<Tu�����2�g��^ߟ;�-&L-:'���0U�[�����5��C�H~��n�a\��8r�9�X��Ë�jj���s�{��P�����B� wd��|c������f|�����*ny�͗y&���' e�U5��7��@��(��U�O>
ꑋ�r�A�&����� �6&�jcfϺ;�� �.]�t*�����d$N���?��_\ikC����:zW�3r���Ky��rj�?�w�9�=�����7�'��8X�#�LZ�:�T"�Z��'�E��,�g��%�0L�c%B5��	�q�m,�YO�l� ��oMC2b�È�S�Ʉ<(� �H�·. 	�$Y�	�j�Lc��^����wj`d�ʜ�<��Z�������X�(�D|E��W_���s����D`l"e�OB`M��wU^@�"j�:�n����%/�i�,݂���/+�-&v�v����C��W�z��h�$�[[�7�4J�qb2��8�������q��Y��E�D����Ҏ���p���:�Z1p�9g�7���@�^�ԪR����T<cYo���T��
 ��^X=�0��S��& IG�X���ir"��lf^$����sf������	��$��M��Q�Ys�@�N�b-	��"?'�����ሼ�ᣘ�]����)��2��¡���|��d��JW�|�p,`]l�P���޶#������v�����Q{�-���0�e�-�G`G����yՖ)�;��O��Z������ӊZ���������f�5�m��%@B��3H}�6<w�"I��w;!L�Iw`�c`�����������8εh��y�6��[RFM����Nq�w��6�cy���P��f鏒���?���y��)�������*���@.D�&�TJ6vDÝ��c,Fp�A"I�q���'�K��$��6�l-���i��MkM)j��?�Q!��<l *Є:P��Z�}�@2��2>���WH��-�D�l���G��Ud�f�o����7��s��S����ז�]Vu��M��pe��y#��V?��hiiud�^Sw���;n7�lcr�'������Sj��?\U^�?!������^Ĝ�b׷s&-9W��n�5�� ^����q�ȁ�I\�d31���n�(CV;����DF����; �X��wM��M"`���I��UBn�E����5�ʗ�w�� ����@ , �z: 8K1A�����6�@�i�h��O3�)*��+(2u�RҮ�����n��~X�P����aM���8TQ����46MD��eZ\(niV���������vܔ�"7r%!C�w|e�]��k]�3��x��C;�!)��ڤ|G�V'����y��n2U� �.U�s���W��vv�I�В�N��z<$�����σ�^�GAhQ���,]��>���i��sj�L�H�$�pn��� �)�8�@�UbT9<��T�u-d;%̮1���2v]xQ�2Ow~p��@!���҆(�I�cc�H��R̩����P�nI��VR��$T%p)���_�g��#;�	�<ɶ8TW��E��	ٟ�M���e �&�޸�4H�嶷r���w��̳E��_���(�.�"�<��#�DRl���픹m�&��x,A���b��ҭ�԰�8�'yܛt�s���\�� �����1$O�Te��P'��K��h�y'��"6�d�.h�;>�����˦�?�3T���hp%�'�g�P�@�o�U>:��a������V��}�^D;T�h�-Mh�P����̾���.��Q�����m.�pn!+�ió���)�P�]�M9q��"޻�F)g$m�ǜ'�Y�:5��lb�9�[WhףG�^��I�v���� a���.�:դ.�����������]kq
��ＶauY��*?�gk��?[�slm.+�l���~�}��E���.�A�
��Uu�q����`�"Oz����b�ɺ<q�׹7�[�4;940��%�b���܌�"XQٺVc8ϰU)�*�o�ښ�fCϷ�Ʉ8�wbj�$?��˓���J��6����նwd�������cm�2K��3��L�<�H�����c�5��t����Þ�d�|��Y�h	�X[��R"�'�� �A�4�_�o6������Z��L!�=ܑOy�WN�yw������I�"m�Ν]"�N�n��i2HÝ�F����F�|86B�UQ��w�����ʝ��5��wrZ1_N��٨�*���)�ϴa��t.��pC�o!�aJ��!H�Y_�5���3��m��0����O�n�H��q���#�t���z���E� ���D���3&r#d�^;��� �7��r,(���A�����$�����&�u��EN�Y0*Ä3������Wa6��Dp=
� e �rTd}*N�=���)�x.���T�e9=���=�:�<�B\�y"��DT�Mhl�(�mnn��4��#R��Md�ae{~�:�r(���o��E��y��"�Cs�P��J�u�����3T�k����z�9+��u3Q7O�Y�ֆ���_��7w��^�
u���I�kqc:��`�=5� �K�����0V���B�as0&�$��*�Η�P�;�$<�0�ܰլ�"_��{��-d��������7�c�����L�둣�e5��N~�����1Z̀��xL��7UJ�>p�;��=�֛U�!�$Q�5�����o�hdF:����P��0��+z�㩯<I����e�q�T�����`�&�]�����f`4��0���ׂ���8BO���v����Q�%kϜ�!_k��k0�K��12<�a��<��`�+�޺�=���no�c��9.9�|`ԡ�h�0�`9T"mc���}W b��52ʀ�_j��P�>&kb�n��|�!��G��c�ƌ�T�CR,����n����.}ޭQ�
�^�UB���
�ő :�4�Zb�k����bǼ��P���º�+�7C����q�Իb'jTOT_*��TҥVu)�.40>��"��6��M�bD��Š��窫��7��ˎH�ܘ�"���b��!Ni��F�#��*.����Uu���E�$�!���C�|���-�VA�sF,�:��1r��/0���°����D.�h,�h���q����,�����He3�d̅��n�P���;*���$�]�L+H-'��6}��w��'�=(�$��ʜ�l���/I�6$�,m8ʄqQFď�� :ضA�B��΀"A;Dv�Q�Yi�z���'
�#ʾ��7�1&8W�n�?R���Z�J�Liuo���99��G��6�Gb�����6,��i�Cn_�!T{�qB�>�-#��P��C�h��[ޡĐ�Ɛ~bF��Z.NkQs��&h<s*Z��F���M�rn�xI��$�&"��g��I]#���1酹~2r�T��0��۟�b`��i 41biZ���i���$׌��Vj�Qt��˽���P�j�8�*o�eA(�_ ���*j�'s\,�V����Z��
C{�W���xd2@��YeA��l��I/ ��x��dR��@lê�%����*!���HF׍xE�C�%W3�.>�Zl���Cf�a�K���-G�C���7����h�=Rɞu0"�M��P�-}��n��� ��	��:�3O;�#��Ƅ�ٽϲs>���҅�����乶Ns81���xE��<4xi�(0�w��z��y���>�"��.ALh��	ynq���
Bɜ�LI�I@1���T�/�7@Ck+���
`|ʷ{�Y�g�,o�J\����c���wn)y8�x^4O�:tsO��Ӽ��%�����Ɗ��z�l���R�ܿm�B�R���h�������{tp�֒�-���k�z3�7�s��ԕ�� �?t�E�Ԉ-�r(�cĭ��
�A�=�`n;A�OL|ϲq3�]��m6�I���6H<���B��&�Ci���(�ӟg�K�!��Oh�C �7b�f?&>����0P�?}��.P����=q[�2�)A�DY����m�F��)Pƶ�mj����roj�l�0Q�P}�|Q��ǀ����-��rv��gSBt�{+����җ;�#f��b��ǔ��w\2�R!'l���?3`����8�����lA3D#9~1ǩ~�Nk�z�"5�����K&9H��25�S�}�^�&"^�;=�!�5kfP��r	$��rX�Ւ��%w�Ua����2ƣ�ai/� H/���.`$ؽN#d0(_��Ɲ\�	��L�E�[x�9�\�̍�!Φ�q/>����Ao�D���'ڮ� �7`b���6�
A��N���_4�c���(���mt"	��e������^��R���pѮ�%�+���ϥ������5/7p,�C�!iN�g� ��2�h�o��M�gЮ��*�p�ˣ�ﲷ�7�FW��L��@Q�����Õ�E��,����몬l�����'A��v��8��,᛽�l%�F�I<�'�3�l{��{��)[�-�8�G#���Z�!�b�^M8�s�E-�z�FY���T`�=O1�%AՅqI��E�J����X�v��*�Ro��X/��fi3(�I�d���-�l���}~w��[є�Ӿ�	�ӫ ꗚ�㿶�_��F ��2R��c7����/�X =r���)DW�R��u��#	��0�ܬ�z�ٝ�zTi���q�fc5zi��D�j?b�/+y���tt&N.�osj��Y�<��B��5�pڽ�U�$����7�-Y�+f=��Z�- �~LkL� ��F��h�c� ��]�����C�`뼫��4�xB�q����v���(-�/x�u�s0�	+(r��xN�P���]����?����'LB��c xs�Z�
p�!�s�^��K�e���Pf�����b��}v�PFF��Vw̤Q�a1��o��D?h�1X��Sx#�|�]�yW�9�)I�q�E��zzpU�wDVJ�>G{����)�+�8\�']b�B�kD'ķr6b�)�lu��kC�Fn�-�9��221U�2�!o�VR��*x8��R�Y3��S *�4����*���6m^9���}���ĥs\��c��_~�oʑhq<Oi�7�ANv��e�Q_���¹!�63����4X��%��^(��t<�^�I�֥=]:.�������U��%R�R���/{��� �A%�	q��`��VP�t�	I݄�|؄��z���T�)R��v�Za��~-8��7|�	P�p��%��ϭY����ު?��5�kU��aW'm(�����UF'.�ksQ6��\���u����*Y���Z�v�ֱ��9W/Y,�R�~P¤��{�s*�J3�R\�Pn����A��#N=�F2'C�B�����m<>��#+!�
o^���^�&	����/�����ډ���F��c�X�)^��Y��Nþ�3)�i��^h�tb�hz]��g���i}i�R2����p��Bf�0�4¢^]�����A�c~�b.�r��4?���$�����f$`W"/F��a��(:E#5�?��^:M���x8�H�З<	�1�.5������4>L,�����'	�)ݵ���*�3�vB������lz<����:su�?bѥG���!��ܿ1=!�`e��H������go�Du���WBӝ�Q�&0lD�	�We� l���A��%ز�խ@��P�:����aNz~���L&�_��꫑���⻧���$������Y@����Φ��hf�RF*�������á���s�!�L��
�:��α
7�k��l�Ӏ����Y�&���<L5���u�+�����W��g�x�&���G�d�I�)�~�~j��JNy�N�k\��X�ͦ� ��q��6t��� =��*�Î��:�;�&҄��;����R9l�+�gL��`X
 �L�\7ؾ{g�A����(��Uæ��$�d	Qq�k��['��h��j�ý�H�K��ܗ�9^��Ǜ�� @}2��@)����b`����'r�.x���^���rS�\��Z�SR?�ik�헽�	�f�=�#�oA[>��'�z����Ӟx�����AAiSp� �|$�!(`����:z����M��[hp]���R�:�J�0�X�_���r]@��g;@�F0��[�c���?r}y+#w�(�9�Q?J��9jk��n�H�a�a{�n	�t^��n���q	2�v�~��Wl&m��ٸ���w_�A���.G��OU�up�sn�
�ڒX<��U��+�IK�c�������(Y�m����@�-j�]�@��VB�y��6Y�
�)q���Zs��tmHW�](߼�O�2�?�ڣ�sr�S�GT�d�|[�����[''���ڽX
�Y઱Ĥ0d�>�L�K��
ׂ�F�7�~=��V�ַ!ģ2����Ts&������N��R`N)0Ǘ#9~�[�%,]��딦Mq5�z霕���W"#"Qn������������H��ml����;��y�rG�O���W�G�t����F���	�MX���7��:t�Pb<Z|���I�D�����JE��	�X��.�����Y��+� �2Zy��[{,������3_Rn��v�U��ܻ��8�u �!2(��.�C�`�	~�oP��,;�p XI��:_W��X�y�`�O��6Y��W+���v �̄p^�*� W��=���4lP�u(1A�u�e>G1݋c.K�,���B��a����4M_�~�W<��4|��Ĉl�6���UI'2�9���6���Rm}�Ԇ�K5�s��5�K��m�d��l�^�4~�"8�����bv�Cd_(��_�Åh���0}I�n�c5?������*|�Aq�Aڇ4zHr����]�fX*O�9	�g�i���p��䓙m�bd�Z���Vp�<���+�æ�3��^*��O8]4�R���"m@TkA�	>�� !�X�B+�$�	��{c�TÌ2���y��� Z���,w4ɬ��@m��.R�ݶΉ���1��e����	����1�^Q��H-٠�F�GCћ�hV-������[�[?��[H�	$ѭ@U>*֪�lz
6�ra��s�3%�VH�p���عP�ޭS�dh�Q���bh\���_�W'��+"�l7.1o��Y�]���@+<��BQ!���Ѥ:t�ŧ����-nY���X\�b\5�Zn��O��ɉ���-��m|$�
��"\b/=ՠq�i;ˣ��ĳ]���N}��0�n�4�L�DT��'�Vp ��x+8�v�B��Y�����o����_b���v������ZOb�EQ�:F�[%�ĸ=qK����P%�dɈ�͕�eL���)ڽ��t_:c���\��	���,��!��Q=4�����~��(ag��:������<��H(s $�()YE9(A�I'lխ�j�<�xE�7���2����S`�-�p��5ڜ�r���~�ˢ�b:��:'�]	9]�%,i���Y�hUGC8�۱����`��t�߬���˫��D}?Z����]���]S:��M�xE#�Ct0ei�O�Ă��%�@"�bȃ�-�OF��'������7S��XT�w�W��ӛip|��W�
SQ|=�
�-;,�oΚ�!��/1A���r�`��n�P�6����p�'���0׬����׃9}�b`f4���W���=J�K�Z��)��(��B[<�/ˊ<��-Ш.����~�P�w�[a��y��y�@z��;��2i�'=ތ�F��q��DPE�\Nb}��i?��Y����l��i5W�8�>og��@���&!R���?��lJ;��u1���̤�	'x�l����U��uw��w�u��ʰ�H�h@6�+y��M��A���QKnU5��'#�
pfK�8��Z��~��uo�s���@���{B�����x2��au�쯺PR�B.��'���-�E�:(\��w�j�<P0T�Z��U���[�
r����Y*Y'�ܫ7�$�୸M����~�rQ�sьa�.���+���8������3-Γt��8ٴ�JI�L�����H��?@�k�AŬ��)�pc�piRn$�65�sEZ�b���r�� ��e@��29)K&c�8#��ø���Y�j�7A�q0��ANXֿ`�'���0H ˱��{xB���n���x�g���"���#�ߨox<�"�Y��x����\�+���`�9��K��ɆI�}Z����Nv��y�p�Z?̞����*J�f����j��F��h��$���613����ow�(#�/@? D��Ԕ�>T[�<8����i�	c(!<��P���"@5����Jb�Tð>�[�`�v[�(HK@7�3@�PhP[-�{����&ڐ"ʃB��P?�~]�2��!�	�H� #^��H�b�J��	aف������,(�Mm���$i�b)+\u�7T�bB�)��8$�ej�q:c��_�
?�?q��А�X�J��Q�K(014������X��F�V%�jr���8=̛;o�V��z8����һ���V&������|����i���$+��2�ݹ��H�ȧ0��c�a�H�C�B��v���|M��~O&���?�	�� Y��N�A��2%Qk�\�'��9�/��l��+$�H�u�i7�mo����rm�}\p}Iz^)�ZTG_������ Vl��y�iӰ	V9{@T4��k��%�o�^��~6��;Cp�.cTL/(x �w;p��=к��rq3Ϩ�UT��,5�!�P�]�.��wJ�ۇNn�e�[��J���PG/렍�%]h�i��\�mH�t��w���]-(��#"2<�`P�,�#����'�ո��x�|5��-���(df@��zN���������$�E7ru����@���!a$	R�6K�U�L� �9,澔Gm�o6Y�����e���$�@1�"��R���h���j�w9�d'���a~��H��l��W���H�_ە_%K5�~��\�L�Xwt}��m�˘w�6�3����i��v^9Դ��Q��+W���	|O����M��u	qpm�o͔��#�Ώ�`�>o����W���9M"��QЖu�?Ua֕G̡b�ՐiPǼ���T��5�Y=|t6}��ѥ�v�U+oa��_'�vh��Y�����'��d��O	���7�/g,Bc��T�.���a�����e�H�d��64k���s��a�ȏ�����Ɂ׵�����͂g�9�Wa�a��D�l�&��!�u�%Q%Bc�''3,��'H��7�ȃv
��/)�XF]/�?Nuq�����
;��w�=J2y�6��W��_�׊��������n%u.y��ށ>��U������"ȸ�h
[�ɿ��_�V���Ǳ�;/�lky���R��f�Ա�	)����`�A�(��/�W�$08�uc�qGV�f����+c<>��?F$������p0��K�,~����5����w�n"J7�G�j�
�G��_?
��iz��A�.����N�$�w��P��LW"d]�>����˹��n��^��nu������TPw��8p���Kb�i�2�]d�Dm��Z��h��i6ay����4Ý$[]CK [KR>��M��
;�GJ ��~ǵ�X�୹g&����fr��I�Z�&��Z�N�k:4��,�p��8������8z1/���;��zp�x۴S�2��`i�g��<*�_fʋȸ=ކ�p�@P�`��E�JA�p�!�6�gx-���o�C�C�aV�\����%�T]�r$�y|����q�o�̍��PU�fb��@��@�ٗ�݄��~�b�y�����"+�ӝ���8E�Q0�R��L����Q�#pBTH{��ʹQ�m��؀إ�
�:�zTSx�q(y/@3mf_��&��_��U?/��
��w�oL�R	�
�����e��v�+��7$�;W��4��=W4 �Gs˚���&��$@bU���]xm�
�3q;�h�
�J�o���G ڌ��Φ1���T�����0��->g�9�̕N�*.A1Ҝ��g�*!�?@~�J�l��p��6,:�/�6�� �Ym�gw�{�slyB�|�2ݲ�5u��XL�¬{��V$w.���+�ȴ��|6!�o�ot�K��x���&6�/���?j}�����Ez�_]�TGV#{������\#�_���=^�4F?�E�f��m$�SQ�b�4�4^Y��T�Ttq`<��k\���o��D6�7LN�S��=�k&�����TU*��U�S�O��Ǯ'��d�����ʯxLqC�i�)�2a�z���<�Wt�ԀC�����ϑo��p7ﴊ�֙�Rq-0&�����K�3�&��-��p�A�h�;��Ii��IK���>O�3��iRv���]��M�ҫ�r��'��H�L�J�{d��Z�Ry�tȴa�>6t��h^������֠��@'��pԬ�H]�,u񘭷�58���M=� +=g��-�@MQy���<X#4�����Qa�83'n#�D�\"������[j,j�pS�Bi�(�)m��_��4�ڲN6	��щ x[��Ӈ�;2�A����Z��T��2ި��jͧ��Z�(H�����L$Lv�ڙU:�ߓ�����"��g�i:ѱBm�s��%[g��dh�4@�6�%�M��S=b<�{�X6�'Vd֚����������1?!��
w�E>eԒ�nY3r�h�k>��ܽ�/�糅�`���������Ua'�*ZZ_�����B1��^.ٍ6D�6�f���9��#_�}����u��Cp�;Tz9�}���r��	��A���M� Ǎ����ַ�D!��h=�� �>R�q��Gߪ"X�	�h���rH���^8@��)&��� ��?.Q~ŧ��R��^9By�X�Hp�]���4�bP�]�Z�**�v�u�>�h�����23��h��M1�q6��f<8�$'j���/*K8FaZ�`�ك���Nn�v��!.�s��7�r�6��0ˍ�["��P�N�r���^��"Z�~qX�e�D�d"���w�.?��q����|ҭLd�l��4b9��g%o)��OI�@5���R� �P��-�#�� �����}L�-Z;e����aC����p��/(Nv�Id�"��U�ҁ�N�Y��?z�o퐦�RH�����.aб1��p��|���������ˆ��l0+@<F怱�(Ѹ��"�f0�K��'�v����м�&Y��ףS�����ꮤl����Aq�u��@>{6z��1Ge�e��khҿ�E���3J-��F�����Bo�Ќ!�K��X�V`����FeH>�*q�~�x���������+�;����D��ʫk���"Q]Sj�_a"v��{(	��^�r1��s�d�z��0����,`��W�xL��B>�����⺣�U[�m	QԠ�hO|= 5���;��Q��W#��r��J1�v23��^�&d�a}5|=��"�����8Q�ơ�'Xd�VBYt���F�حnu��B���w@^ƾ���w�]��؛��<m�|y<��.٘�ۭ�8�>
z�@���"�F�aу��� �ο^Z�&q(2i����h� u�Jy�.�YҮS�,�n�'����{N�ȣB�V�W��0�>, �ObO��������wm���N���tQ~V�g���joĢ���K��14P 2Eff�U/�9��&U�E_�槎'��b�d\�>[�_��=�0 W��I�G��'>W9��c����Q� ]`R=�Z��Ϊ��Ahկv/Ȏ�0���\r�IRS�~S_J�%�4��9�&�eSl�9����-f<"����%E�Q 5�����Qf�}�?
���.-��O�,�MJ�d���	H����`���x]�[?N�������� A��*C���q�����)|��t{$ӎ=F�C6q}	�[��~҃�p� j�9j���&��^���"��_%R��f�"?��>�E��7�P�v�=F�2����.�3dkL䭴��,�g�������ۮ����W�$/���ߏ �J�iƓ6�9��.�b�ny�;�3���9�}�ܷ8�� ю�
�x1�[�Yy��i%U�աN�Ds�~5ݶ�tb�Vek4�`�`�+��d��b=��z�O<�픒��#A7����'��96ݱ&�+{����7��@��6���z�"�oJ�5�-h�\Am���|GL`usrQ�rk[���E@���S�"y���/[�5����I��}q(������\
�>o}���b����$��%଑Lk��m���-���26��uS�;�K��9�S��{dOG������� l%n�ϭ�=�����)�E���TЍA�4Z���f�lŶ��͔����k�f��=���'ns�ynV���5�h�8�U��b�M/X6��!�Q��zx2Og1���z�X����A��9��`���uְ��c�J�_0%�TR�����6%)�F��U]�����U����?�)��Ұˍҫ��I�"�E)��I�Fi>�t�/�8���>�:8�E�u��!��#N��*��Н���QPf��j"��_�I24�����V4n��h�Nw?0�<F�(P	��Unm�7�������o"3'�H���2l����d�n$s�]��[ �q������2��[�P��r�؍X_�܎���4�vF�#���**��?�����(x7�SJo�����1��if���Z-�`�4Ae*�c��T�V�����ٰ���������v](���+)�W����$ѩ�����:a�3<zt����],C�J2�֩�Tb���kS�6:�U#X1̍q�j�x���l���E� 7�.|���j��Lֱ�4��1u�	S�B��j4�~ڢ�S�N�=����
�����L���T�v�	,�9?����]=$J��N\��ћ�y�C�QoL�e�c���$��ڑ��rFf�×�����������<�J!W&����E��"���InѼ��Ԅ'��)��>�J��~'�/�v����!y<'t�Z!lt��H\���7�'\��O����%̥z9���� ���x�Y�snn���B<�w*~�h�Y�`����u�r�6(�\���T9n���uˣ�)J���ĺ��P�a�}G�� r��0�?�����x T�f��c�dR��-�h<n��@(��^�=�^����u���u�L-'�R�#A���'�`WR
�����������
�N��i-L����ba2���7��h�&��km笳�\� <	Y�%���̕�|���zE
C�x�g��N�k*
:�}	�4�����@�y�0�X������W$�9QK�/�TH��=J��~�"لtO�&<��W�d�;�@�8M�� %.���R���ϭ���B!��V~��:
�O/������ �d�mD��K{�9x�k3an�m|Į�E�8Z�V�Wa{i���,&0��;�R<	.5�63����i�:�(\O�	�5x��rz�*�^�8�V�a���v�r&��E�Y��xo�(��'|�A/?a�{�e�pC�Y�����0(H��Ӫ��	�+�S&R�u��	-d��ȕ:� Q���q�G�e����JKν� 4�n5�t���p��yt&tG�y��t�U{�A�w��	��;(@�}�H��6�7t�E��>�~N�;�I��e�4Sx:QN�bk�����S�p;��0W�R	2���ԉ�׳�Y�R�V`��v��KΛ�����P( ̂U�\��݅����[a��h�\	�AxDm_<�d�l�O.ha5�W�^ 9A,��'H�T�y:c���w�L�˝i!��w���rZ
�K�B]}�ˀ��hC�i�(����gFFJ���"�y�eiw\E�Z׼�"����c1l����p���}C<�_v�v�x1��|��0ߣ��l���n�C�ņ򊂞�5�����7�(:im�a��[ �&�׾�5i�E|�[� ������q�T\M�L5{���7�Υ����.!��CN�r��E2H1[N-V��n�z�2L8���`�V�R�d)��p���.��A[����*��[�T��e�����r�M�=B�M��>g�n��8���_+|ӡ@%�iҮ1#�������On�z�JQ$�Pwr4��XX���K�4�I�\�=�
/�ι������rn���:�zF{$�M�MȺ&�����)�ǒ�SB����gk�U_=dN��m�.9W�W�AI�SWG-H���N�C�Tq��Cr���'�~�[ʴ�]0p=��X� >'���kR���bd�J_2����*[t"�++��)�<�Әd@�����Bb�cqX,b�E�����i��i�?�L���(�s�߯1WJ��Uy��Ռ�I��4Z�nq@7����Ս4��W�"N<i\�V�<�[�@C��&*c&�������3�L��:�-&����׬�K�+{���m�Z�_O���S;������a �'�"��3��ѵ� t5�F ����3b2׈c뗔&S����w���'s�w2*����[f_!�0�������P��\vQ�5;��_+�6�-�L�3#ܻ�$��:i���	����uU����3��٤��	���-�nGH�.��S+�J�V�:��~0-�
�Y*C���Z�п��(8�\��G�4�LK�|f�����G�od@�}�8�`�����(r�QW����a����m����c��f5��J�~��U�p�f4��Hi6r���,�%�-Mk��7N�7����,�S�P�>/-恫۔*�N&��(7,�����`΂t��� �أ}á��$mGX��iA:Vw�
�� �)X�l�Эk/!��C�IG�S�W��J�[�P��Q��G�i�ް��Ġ:��^�ݰK����/=�D��|���bpTDǫv�kì�U����A�����0�� �����������щ?mt��_K<��0������N�;L)}ϰ�Q-B����PQNwv���:�j*�.�9s8n�n�t��2����)r�y��#Hθ�95|�>$�!��ٜ��	(�Z�c.���<��"S�9o��������AX���~�y�;".���(�n�m�`�yi��h�6��7�(��@�Es}]]�s$|r�M	�	���|�����e3)#qPeL�
<�;�D�S�$H�ǽ���1=�:#w���:�rN�̻D(C�$�ܪ\�Қ��Q�r�����e z&�$ml���E�{��1Kz���l_	W�D��� ��Ѝ ��Y8[w=8y�GIPz����jWy1�}��$��ԫ�b��j_�g���AH5����2���ʊЮݾ�	�$���!Ѡ~Y�l���.�F���!|�J��&��:���O�R���Vs��(+=��8^�,&��EG�6@���ڛ��3�5A�����v�o����|�A'����m۳��7���}�JY풕;��x��̨�[y�Ϙ�m�\�y�|�x��
�
|��L�ƴ�|"��!�����),�o8l�֟ԅ��sX������c������zjںa��r/��=^V��rUǶ`S�0ګ��3J|���x��$������u���	һۜVȋn�)�]]Q�HR���j��=<*d���-e=P� �?�c� ��	���5D�U4d-�v�<�	�r�l��0&��Yr�v�P�y)����<�d�������K	�)��+Y��`z�����yIPD
�t��|�I��q�k�\+s��OMXԒ�D\���u���+������|���Y���%�M��Ȣ�˻UZ6T�s��P��� ��m÷�Xt��K�P����n�9: �x���.*P��a�.��!��Z��'c*(U������X3��E��@;U��֩ǰa�U]U�M�n:�6�]���ZǁOp���������<�G_Ο]C@���lE?�K��KWn"y�į�{��xr��+�w��W�+T�v�?�����9E�����i2��8w�p_��65~�΁�B�ap�v���&}�ܯ��1,��ů8-�L�`��ڲ���oc_�i���z3[U����b�ktG����5|{V0��+;��#"p��]a�Ta��}���e,MV�oK�+KpԳ�����~w�`Xfi�=62�`���Lz���u��v����э��U�� Di���������G2@�El���b��<uHI ߀�Mժ!��a-: baMC��2��X0��p.sP���EкE<��K"����P�Bx���M�Ǳ�v���d�%q�$�[��}��(��N��][-�)�СN�)݌�(R��h�ɫ9��wv�v��y�Y��CN�NY�	�� )U?i���ll#������Kǣ�2��8KS��Uj0��7<Y�G���GI����j��k߸�����K��E�zĸ��z��#�1^>�n^
y�\8B�U%���WF���I˖q�Oӛ�%��Z���R�y<Z�����C)��ci;�P�4�������V?��v]4{�v��aC�^#cc�T���A�����S�v/��!AD�y�Y�/t�ߠ*-����|���	 �&���,��\ⳢFt%5����������v�݄TL\/���ppT�����S0X�Hg�-�Ҕ�g������c��m����4�2�%����d[*�#^5"{�0�0B#��Vl������%赿�/��w�����(ޓ����;Gɞġ��+$���<��
�uT� �L>�m��:<nB���lH��/�q>_~���l��/�8�"��>B��$].B-uU����яz�,~DQ����S���o�D�$�7lsւ���V�t(]6�"�{פ���G\�����%�_�Ћ،���Ƶ�qӆ����c$�b��J��X9b��C�Җ?����9�~���u%6B��(u���W��z��z[�����v���]�������R���<�$��ؼ��DzB"�Y���P���Q��k@kle��j6��B(�q������.����.0� (W�x�;��k��[�0)���Ҁ���G#�vm���X�5�Nx{b�X���JSVRX�U7����sa������k�y��Ԙ�_�����I/�V���K�M/���;h�����9l`���ߑ��>0ڞ�����o�ev#~HW�U)k�k�'�|m���О�=Y���B��EL�n�N�XU�wl��7l@x(�۷�Y��Ja������aJ�?s@_���D���!eh���,ߔ�����a��Q�����M�3� �T�t��?�9b��K�H֪���]qIv�Rݽ[r3��e�
�m�V���/_N�I���usņ�8��Y䤁m1Me-r�Ϭ�i@p�`��$L��!��t��*�b[�A��
e�^k�˵�����hG��HoTu#��� B�F�
'Z��<&6'�#R���bV�e�p0��ǐj'�R��^��cg{��in,j%?\.	���I�!�������xIv���)�@��٬`F�!E��_�3��������e��j��@��` kWu� ���y��}��Ё�{�?;�r M�X�*o��,� ,�	nC�тz�rl�J=*��h�]��Q���IٵX����o�Dy������M�!�P�{�j޾D�-��c�������K�A��m��f=�Pb�3���
�r%$��hE*�*`��x���D
�N:Z���^*N�;�)��!��"����9�t��������J����}����Z�Bb�U}S��n\�Jh���iV������)(���h��������S��A(�%G�T����ց�dE"�޳����l��p�)W�ɠ9�H��W����V�Vv ���#4�Zh����ߝy�00�`��tz(�*�dudwᨓSq~p�_�7^���u��/���R𢡄l�-j<TSj���Zev/ҵ�l�h��oYK�f*R,���� c>�΃E�t*V7�(���XG.f_��x+���1%Ui�TL+UN�y-��Ӊzo�n��Rv%�|fCC4~Ͱ��۔L[l���@C�<ԅ�)�_Ucl���V��l<r�浽��)��ܭ���=���\�.�-3t�����]CUf����.S�'>*f�+횊lH�f���Ưӂp���q�sL���ya�`�y����!�ۆ:��=��9$U-� ����9!�Dӓ�A�^�;��t�&Z~�����d=�}/	�$�?;=�S�����p�.��^�c�_Pz��&��M�=%��Ժ>gW"6��؇�'g��p��B��02����.�wq.ΙW�K�������^�c����g%Ix	�צ��Iי�:���f�03z�0JF_b��q�n򋅔�P[Oz���Ɵq�v���sx`5re�������KzD��n:�ӎ �$}�&���V͕I�˝B�ӟ�|�ZAc6�P��X�?�m�!�kp��Wu��B����+�|!�@�Q;�i�C-1�`�|�n&!�k���n4(��4�v��'���(9�eKqc+�4(`�m���k��ԩ��Z�O��2���&&WV���]>"_���l�w	�=���Q�4B UP��B��~oO���C]�iΌ3���]���Z�<�l�26����^،ˠ)�4��1�� s�[ܘ��Ϳ�fz�����׸�wϕ7�n$�мϚ�bҮi�\�6��d2=���ׄ�v��R���MD��ŭL�ƗQ� LdK��*/ `ݠ��B�c}l~�����ΜИ�ǙȦʣ!�w��e�2�[m���6�)��S9�r��2B�]K�>C�яe��:�<�p��<����k]x��F�K��YR����@�=Xܹd;/Sa����S<�
����Dp��V�^
Cg5��v�3.cu\z���Dsk��l�A��j�Y�OO�o�ŸL0a�9�5��j���8}�4�8��6,�ڪb/�w!J7�q�^ǋҙ:J������,ģ�yR� ,?]����8P��o%�D���O�i! Zp|���u�~�.�)D
�?�bn�ɔ��LRu]��d��K�(���O��1;�F��������:���{�6�-&Ψ�Olo�aMؗeؔu�I��l��M�Z�_�'p���3}��^4&h�G�#Vf[���p�/���h��C�Hg��+���}�pT5�A�;�v*��g�JJ���`���Y^�}(+����]O��SE���[����:��"��� �g����'F�Op��n$���U�T��$�O�Ff����h�u���X��KW/R0 �����ɶq�53�^.V��yt/r�
]?�zB�@�4t����e���}�u?��߬��w��4����G���s�*R퇨Vfʯ�/�5�c��u3y�%�]�&kÀQ�oZ��r?�R��+���g0*{���� �i&�m)�3�o��,x��^�އv9:@���V�RhQ�	�`ݑ҈������![Rᓨe�/�&�B�`xt�&]*Yf���:U|��-�ف���%|r��7�"k�rfx���P����O��б�,'O\^�v2<w4ƌ9]ׇΔx�ן�r��?PŸ�`;��^o٬��?x��ߑ=�	���&�
���e��p]�;4ES�~F�|kϛ�����I����>�-?YbL��G��������!\�C~��˺�>dK�5�I�Rv���?e��|�����1}�6}���"�ޑ��{&:�M�8�0�ٹ��9�i���9�!� �9RR�/��2�q��x�uw�/�M��#���)�)�?ϡ�iJ�:���d����+v<0�y��"���g�/:�V��;K��F@^��#��_�f�sPֈK1D��<�p�ppvX�VB۸%a�K���.�AP�s�g���E�>�@ei�N����JԌ���{@l4�W��FHi��/�U�C˭�F�Դ/��s�0�#��+gٿmM&�6���
�'�s�y���H{[d��=O�r���p������/�Z�j�K��L.�A����46��@��K)�~�g-?ƛ��e\���,�{)j�^��8*����?Z�YjR]R~�_��V5�Mh+ھ�M��3BP��x��L?����dϠ���"=5���V`C���c�����l8^ k(��z�s��qeV�ª[I��̘"�l�&�r�AE�`Ȥ>�[+�8#*r���ezaP�x$�d&ƺ���RY�tIP���k��
�h��fK�
�7
N���0�V�/v8:������gr����ODΠ�0Ep�Y���к��U�GOUjnߢ�y�@ݥ@�%�pβ������W ��D�H.��8�_��r #&O���H�d<�]�TT��K�ƀ�P��H��!nL�ڌ��y^O3@ܨ/�5A�F��?]��lcVǤ)�����ϲ�@[b����;$9�({��k��w���Q�����_��K�:G ����0X�"�r�\��(���*,w��m�[�:W�y��@'��0�>"<�)��St�jSwT�j�*X��~߻�%���&�f���(����;�׵��!	3մx��s�cdO���� �S��M6�L1�k��&�ew	���1���T��vi�bl���^�5)E���e!��$h�g��;Em��N�e��l�P�l?H�H� ��E��M������>б�N�%�s���a�-t��֗=�>��a��8v���/
8�=��$���RM�$S���&l��b�U�7���h�[���?�B��Nf�4h�z?
�����&�fu�`�xܑ�/�\A]S�gYr�ȥ��h�Y!�hK[����Bo~���P�.����Ջ�K���ĭ�$�$�Ll_�_J�D(���>z)��3Pʝ7Ƈ���;(���N,����qtd> ���ť�����;+�2�Y��F����aT��<T�T��4�}c�*ѕȖL��NJB�\,!��3��@:m4*;�	�]��g�<���:����_{½��I���]a��\�f��v2�b���ϰ�c�5�$֐�>�%���#O���.��ӑ�� ��EY�͖-�G'�;��+i�ٷaP@A����I�(8��W���v�&h�������� ��W��{·�*+��Ø֌9�ȇ4��Z!�T&JF�2����񟭶�(w�"��+�`yV�CZ#f!I ��L��Ԏ ���F�&�{�My�d���=���-5\�k���^���w�N\aN������ũ;'I�f�E�\	V�O7I.�\jT�K�(��Bz1���h�<��,��@�F��M�z[EJ8�" C^�qL(�t\OS���x��9%{��v��b���᳑�2Q�����D��k�L�8�d�A2O<Y籙� ��֧��p��QL���H��z�$%q-� �n��^e�(�+��T=Î��ݻ �q.�e�츗����/J+ �ˮ9�+�$�<�	����?^���E�E'�]1T
�_kUU���W��Z=0��f˻/q�*�m���Ǜ�F2��������e$CN\:�!*� �;D�ge��<&���z\a�jp�K'ƭ�^�vl����� "U��t��ue�o�'��r�s����`��q$Έ������<;
���6�Zl�J�q�w
��s#u2�=0�l�Ɨ�#�0D�����m�6cȋ���*�1��jD�{�?ՙ=#��%+���|g0���x�R�>��hGI�v�����؜�x8:�3�������؈�W����"9�8yMK�S�כ�x��G^rM����O-�`7�ҙ��\�ov$9�j���U��Aj�a]]9t>q��|K�j	���0�/��/+oi��(��W�<��N��j&�����a{�9���O�0'.��['��ş.�T�|�ʃ�mQĞ&1��6�������R�B������(���6�:���M3N7�zE$vij�:�D�|���4@!x�B��1LZ+���6&8�\'�w2���x��� |���y?䨛��V�	��o4궞���?��Id��c��Ym՜P��z��d��_A_4(?1��
im�5�p1�{��,���z���\���J~>m\�)𷮪��H��G7�l+���c��USB�i?^�
����{Q���
2�M%Ξ���2����['	��Sl�m)����<1�����4\����g��fk�����J�V�b,�^2
���QV�>N�"\������1���QYt���tH���J�G�ib�C4(���IBX'9fr�~�e�E��1|��No�Zu������1��;]��a�/��N�E����i���v[�w�?9�����'�� �V�-������$��rbbǂ��h��i�)	/X:��=�6!��Lg\�5���φ[�a1F�)��՞f �X����"��ih����j辒�~N�}����Y��<x�3�W9X̸�*;�����Gb�$�o|� �,Q)�7Ы�6�CN|ۀ����ʽ��g�Y�?��������䒴��>�|]Lu^���h�F=;!K4��I�&G�lG
�����:�9�4#�	p�<�o��ޞ�-�k���E�߆�L�`n���=��j|sxc���Ϟ�3���f�]` ̻C���-�k�ܻ1Ns^�g	�#~�yp��M|��q�S���|fs%<s7~h�PO9�i�B��}K�*4�S��)�0�eY?���k��J�������'&�����;��>����0�Ga�����	��(�8j�|QI����8?ӏ�e�U��k�E\�t�R�/���@)����Du΅K�2�VM�K)����e����)JH��#%C����+��O�Y�#�FCN�^̆W�w�VRS�?�Hk�@#�2��W5��զ��UI��#9�U��x�(���/�2�X�vn�J�8��쿽~$=͕�����h�+�Y���P�R��MS��5�UWow��R��L)/dO�����#v�9n j zSH��[}.Y���y�GÙ^:�-�i��t�[��um
����rdK]�� �VKĞ��?`�A{e�mb<!
E�p�W����o������<�F)��Իn0�\�)�N����PI��G�=@W
�t�Y�l���NF�
���Af���)ԙa�8�h���qn,\��Æ��-S��B�<�T�2�y�d���2�+`�K�8kMXc�8���f�-f����[My����dm��QİA4Y��I�b#�}a��ĭ�F4��	�.!ʎ��k��˶YXq6�o�F�16N��MW<�|��:J:y2�{�x�7&�j�>`�V�d��%�@���I��l\̐�]ls����RM���T$�s?��Gس�5M����1O�$�57���A�e�K7㏅P�~�i����h��1�=�-���o��������ɤ�o��j�;�5��"�M���'�Nhҙ>??9Ox�+���d�����}FZ�l�ob�f^���p3��R�j�S*�:G&Ơ��P�=�B�Zq�������쓦2k�x��CLf�W�!q[0%"��d:�a	7Hg�M��q�G���_T�t_�7:ўW�|����VP��B��T���j�"��4��c]����<�8Ά:A�j�� &3C�S0.�/��TнOmJV�v�	zJ@�;�v��b*}ߙ�nr��AX�ہ� Soj�a��������!�S$�t4�K�Ԙ!\�F��s���x���]���q桇�������BG�������2LS�=�s_�&}�+��o��~BcC��u�d���|̧P*Ru�H;�{���-���=����.Gv2t�2�ڐq�H���D�3���y��]l������|rot���TC?�W[��Y�b�Yu��.�50�-���|�	Fƀ7Ƣ��k~��2y�?�S�C[C�e��B���d���,���U�*�ba<�4��4+��}���q�b��ʷ�F������W�����u{	`�R���#�Lr��M������������v��;��h�@,�z{yi�&�n�T̞�0���֜a(i�6�\�1�v��;,����]p�?�fi�Nf��$H+&w�	Ǣ��&��~�|2��$R^��{b����:���B���9S6e >��13fk.DM"��דd�PWz��@>��}��r�`8G���;��܆��R@��5��(�5
�r��. sA�ez�E}b��'�I�8ٗ��\1}��E�U.��e^�s�qWJ]'���f\1���9m:_�9J�����C��������
SF���2���378�R_k7�)x��:_�'�^��x��#�uA��l�(��N�\�˙�v1�?n�5u�4S���z�6>�u�T�}���ZT���N!MGGdy�����߮��з�q����@P.O�kl�vjd�#�`p˙`v��\�,H;❵��R���C��0j�Ʒ�ӢY,��X�v�
�׳s`���I!�ؠ�������
v��'�R׫p�������É^6�]��-�rh�z�E�"��EڠJZ�閹�q�P�X�JյtBU�r��|��16�:�u����pc�b���hr�C)���m���ҙ�'[~�W����v^5�`&2f�G3��d^����7���xĂn�8���7\�tl�D��b�q��Ĕ<�gXjikޑ�g�4z��Y:�3Wb� ���ي�yF�:Bm���i�7nw5-�%(S*UG�NRn3�����%�c�Y�M�K�-p#ݟrD�G�Ud�#.F�O_5�!�=)�p���~�w!�k�V��x3df�5�=l�ŋ�B �	1���׌V��r>�.���ۨ�I� ���D�d���^������u��'4?q����:c�l}�A������!�X��-C�t�.(>F_�Y�:���~����/�Њ9G��C�0o�z�	��B����	��c�CZ�-a�9�!i�-�ќ�;�;\6�X�;��𵻭$"m徽
��h�`'fN\�~�]� H��\��t��
����[�t|��pHg�t�u�m����
��� ?6<��U�ڧB���oJ�tWpp6Ԛ�k|K�U���]�ʯ�Dc��~9���p��0|��ǭ�4����pp�c/�ш]���׶��3�勤��Qt\=�(�l�F$'�H1�$M��Ia�k�P�����A��7�gv�Q�gX��{�M������(nH2��O�>�jڸ?���=�h^%BĘFt��e4��"xs�CnMh�=�9��>�fzrS2$��*�J
�l�f9�K/%�a}DꬕC�"N������vHEM%����Ӎiȇ�V�`4��:�Eb� P�G&�'es�zz*Y��=MwE�`4���Y��e��S�Q0��#�|C\�C���KJv���������ӎ�|�<vɫB�U�o�Mn��eGy�K���7-��z�	:8�M���b�M�܂Ra��k�8No�Y�UA/7��eme}���u�M�4��$�]k3/�6]�S�8�N���e���"��0��#���$n�s;V9^��6P��4�#�j��^�r��#9���E�a�6�Wi���S����F�����죸	�w��K��M�dn�>$_gL`��gE^�w�_6�lO}�G�W�E��FP���� �C\���uk9��-�j�T(���RWM��Z���V���[�������b�[������ɫ��.�*�!���s�,�2���\C<n�̩��Qcqd����=���Pٴ�-6G��;��%f�^�Gg��l��ڼ��z� �̖���~8haF�M����^�_�p��+��~��Ԙ���;�� �PO�B�sq�E@� /j�Q]/ʖr[s��e��®!?Y*/�DK`z��
*WEߞ#u������3�U��P�?�U`\��o{��R��eO�7~������$���[�ŕY��X��d��)wUB|EEh�ͻ�_�_��MR�b��~�/��+ު��p �p��@��+�d�b��qs��{pBL1�:P��U2�;�*�N@�u���p�tv�V8���+�\_���+������s��3��H8RA���E�=�GR����) �-�Ku�����ȥ�.Dp�u����y���A�� /��~�_��b�%�,��4eZE��cY�A���?���&&8&B�+M�>�Ф�fݩ�AIS������ �?�	7��g��ڂ�����k�c�Od�{n-�)m �+��J�V����-ZGE9I{p�|�Lz�0Nl�q���=�A�y �CL���e�d��/��$��P~O�b���G�o���m�����נ��4o9¥�ௌ	mF�?�,��V�F�ݑ����P����$L���L����p�����Z�y��m��*_�K)��gD#S���?��O~H#���­˚�d��f6Lp��^��{<��ÆR� �|��]䝓�qyS;PnH�oN�zi��	��<{�f�v��Ǭ9���-=C�a!��W�t��^�����g��'��iMTsZ��r��FLxy?�n�[H�m̓ �ؚHE��5�}��@&��{ �j=�g7M�H�:OI3���K!;.�[��h�`K�Oݮ�D�Y��;T��� �& A�_ ��ɭ亪R�\4��Y��H��	�RV��0bB��Zth龱�䪡�o��MP�9�Ԋ����b�p.n��X6Z������\D�&1V#L����Ni���&�����Iam�{en�R���~�u���\������Bi����r_t��)���ހ��E`�EưQ+W������q�r�`��'4���P�i���q ^�����9i����M��^��uc��=�K�E�[�j���=�7m�!�P��V?ώ��c�U1���2ƹ�
+�A,C?�}B�K���E�?r������0C����B,r����+N����uʋ�U��Tl�lKA���ޔ�~������X��ֵ ��C <1��St����,?���
��,s\�@�v�>  o1I�|ǲt�M� �VB�%��=!�⸼v���ر�����-|�L-��\����]i����WB��u*�OHٍ��]���[ia��T���y�_ -�Mɑ�/	��;oY��i���L��E6N��G�}�L _����t�='��!+�׸C����7�d�4;3�j�%��HXQcr��{�1m�y�((elo�9.W�i�K�_
p��$�b��@��U;���@������^�ԗ�y�񚒲 ��Q�3̵�T�w�tO64�j�V0��~���k���Me�?E�
DN,�>���M�;�;��뎘pY�fA��b�pP���� `��S�V��Ng�L�t��p�f/��;X�;ʰ����*��4��{�V��g�%���7������뫔"�v��P9�Vi�G�27s��Nbx�@<T�����Z�S�>�&��S/֧�]�ӖP����LF<9�/��;ЭP�vE����>�ǽ��� X�����&S���P�u�m���&��4���2k�4aיG��E�:M4�.�� #=L�h�aC�H���d�'s	��,c�G��F���G�fl�H��w�z�?���*��
n�Ti���NIk��8�Tx,���j��.m��6�+��3����^t=�&�*��Xܸ&ٖ�́{
�Я�~��
3�N3�gǒD�A������>o��"�kh/�؏7�����"�1��S��'��P�ӮMo9_+�s�����础BE�:��-D�՘_iw��7UU�]d'T��¢툾��U�h�����k��5�4�%��՟��|��J�Z��I���.�g=����M��c�x������K���&�4Y�����s�!X�X�$Ǐl���MB�|̸9�:V�{�q��Ljsvc��n�C�����zz_sR�rn����4�N]�x��G�Q��6�38��߲�*v5��(uL���uU�y��� Z���z>����{l�lϤ��>��M��[)$�ށr�/Y[�\�P�+���Պ��#��~{�g�۵ep���1�\I�ڍR	�����K	�^�'���k	��v�~^�HU<Y�����<K�t�pCc��@�q��8����7�Wԍ����N؝�hX$�`p.�����\�Srm�a36`� �<�X4���]c�ip�s�y~�)�Q�S�f���CЕ�_��sPD�q��D�a��C�&�xe�w��SN��:f_���A�`|������;+���
�[��!|��Z�̴�F�~��K�2��s�!��*�p�
E��pXV�c�ǖA�m���{�d\��)�?A�]�I��Ì���s���[A��f��������x�mbWcE�N���������g̽������-5r�7o	��δ<�ԭ�;�i�	Ht�C��	N�=��!'��L�X�,�w������,B��/�О��P�~ aϋ�a��V�,3����Y;�F�
z��Sq��wG��M�v70��k�oܳ�����O۬�D6)���M��� �U��&8C�&�Vj��
E���E t�%��6�%���_��#���K���̾�T6�K��q\�KZ{�k@óc�a/Ziv���ÚV�͚`�,�@\R$֦x�U���BT��^�Cd'b_=zvM���v�.�]�k8�L,�H��l�&����q��<Z"�� �aۂhD�{E�
�«��\IҤQ�ч�Xp��׆Z7 �ZK#�m�~d�3�;4��0��U���|�jD9�m[���.ڸ�U�:M�Q�o'�."�-�S�NE��wT� ����y���0�@�<�h�����}��e�d�]=u�I'њ'��j�4Q>E��܌y��d�@a@
�� ~� ��a�Lqe���Y~��\a�����yJt����
#��cI��ӚˑW�4n�Ї��]�&�W�oG��4"H[M�P�K���L.�_���N.��e��BSZ��Eçgy$)�Y�<���z8e�F�u0�q�b������Y��8cp=6���	�w6�n����a�ta�2�p��<Yuⷔ��[���7�,s�1I�޼�K�?l�M�柼Kt�~ ȥ�ٞ�0�L��' W��_m9U�c{MdB��N��a�0�����W-e{Y����{��c�d�˄=�4M���V4=PU	J�w�Uj2"�-c�
��������22�A�E/[%�:���
./��R��o��C�h�7�pƐJ���ͯ+�cB��Pl
7�Y������6E��v'�GЍ�:�ѻ�ey�.�8��d�w�W���ށ,(��#��ՙ�]�Rk����[9���9� ��q��cZ��#PP(��߻E�{�C�_���_O����� Gp����N_r���G1�΋:R�tm�T�K���K�F^���(�&=�&r��2�}Ӱ@�M�n�0>Z{�'";m^��K�_��~ ���ٹiTB���+[�ĦsJ���t��5�7p�MWXJ��B�̌���Ka�I�z�bcvt� �Ӂ�T��G�s�QK�L������y5�QW|�G�!����Jޔ:N��%b�����֔���^$��N3LV�`���G��0ϕ�%g �a�L���9 ����.?%6�5��7z���H�nc��Y��.%�v�w�v����~�!0ů=���vW�-1�C-���V!�o�����UCi���	����g$��l��mBq��3-������7 $��EGBZ��4��uQ�8�����V��?�,Z������ j�A��[�,v������+�q_�AGT����zEw^y�_�_�S�ʪ��஭8R(��"L0�Y���ׂM��
�舂�89l2_l=�"�U���SoMpО���|�1�|���j�)5b��J�.�'��p� ڽH.D�bqw�ـ�ud�h�{~���' ?��Bf�$ |)�X} �(
�!9�.d�[�o2)���M��b+�9�*(HzXN����F�2���jل)+�r��)x}�	n�l鸼D�P��ި�&�x����X�gFQXB9�@s��*��b؟�e���X=D� �	$�o9i)��ʔGELZ��?ơU	$��3��u�g�Q�����&�{el�Աs�
KR?��r?�ޚ�g1T�tN�HJ�9�>��~��%�����h�Ok�6:�]4������ۿ�J�E6Y:֛U�3;ʽ��z����W�ʌ��-�=rr�V5ڰA�․����\�]�G������ %��U܎���7W��wd���R{��]���J:���3�!}���a$�Nݹя��q�O�Ŗɺ��8m��Ǎ̚! �v�� ݽ��F�~:�n��Z�6��v�{5�x$�G��F��S2�z����X2;��lxݨ|�F���B�@ě��^fAi}H0��-j��Oe-��f�'<���G�B>�c$�M����s��9贾�A
�Km5�@
s,� #c����$1"`T��y��jr�.����Z����-ȩ�0'�V�ӎ����������|I���d���c�쓏L
���d���e�!Eu���`���T�/m���`�Za��	�p�ЉC�����XE5�C���X�q�����9q�LZ�	Y5g$c��W �UV��R��o�Er�
�������펤49�7{Cb�@��8,��wT |^ñ����T+1�����B�a��UQ�i���lu<��\��M�,���`j0:�ۋ�S�B��1��Q�Ϩ!��2	�>�1N���_$����|��d��G��L��f��7�����x��&�oL���Y�Ow���R�~4�9�[cN����W=�,!��W��$�@��c	�D\��#`֯͂Gx9 K ����z����}��=�CwǼk���:T�Ĉ:�W�ߓ���=�/tI��U/CJ����c|�@S�1][���t,��8R��ט�䏐E-糂}@Y�j�;�Mup+�.7�xe�Ǽ��0��緇�#bs�x� ��6�k�����$ߵ$�,CI�����5L��*��n{Y7�|T��j��(g�3T)ٻm(LrԄ�'�Fh��[֩��n�{z�o�ŊYd���앪׋i�Ո�(��3�]��`�*#�� 
Ƹm8'����t#h.Q��~�XVs� g �,�j���4�*�چu�F4W}s��>b���`XC!o�m��M�IT�3�{� ����_����i��Y9��T_%�^|����lwe!���S�d`W�p��.uW����aI�I��eN'�KXE�M��e�*��oQN���2j+�ϧpj���}B���p{�=M��<̪v��V�k�H9�'�~Ϻ�7����f|�W�dX+��O�����'�:�Av�!�9��t>�_��"-�ϝ�jKnu'%���י�6h\Dy�R����w��F��+"T8���7�㠑0�g�����C�\�A���K��>���I둯5;�쵏���1�b��ݹ�V�]ݗ}�?�`��
�
.�!%][v��^쵁��SY�>&Ġ�<R��n�w�T�H떳a^���i�I=�=ET�e��|Y#j܋��M��Ş�APcx��5
�}!	��Ĝu�1��שlY�|ɉW>7�6o/<WtI��H��h��] �b�LB���!s{Gt!�ފhL�~U�EvP�.I������:�-�
����dq?�?X\�%nZ��b8`�z�qxkg<V���$�a����E��ŝ�X\�'0��ׇ���|g़�,����V;ߗc��0"����+.Y�9kJ+��E cР��*3/��+�G���hKJ���E\��f�m�5XrP�D��]�r�ֈ��5�8vb�@��'
`G����Y������A!�P!�>¨��As��
�W�7�U�a�C�K���W�&=*`þ�B�Ml��}�U�B���f��8�9���%���g��!"(NI�������O`�u�l�;V����{�f�r�vz.��G�̙c��}���f����*,�8Т��������S�C�0��Ż1��s� ^���f�(�N�3�f�C��쨮�[�}�6�1���� ��&���&�ɵ�>)��c90�E\sg�����]�Bd��$.�G�a4uq;9��p���F���\U�d�/�`��J�a��Vz�m}in�T��h���>H.�N|��huڐ���]�<�����H�U��j����I��or+�c�*��9I� �.��8N�ȿ�y���,V@�{'+#6D�zUi���J�%x�5�V2'ۧR��r0����ZT�5����@��m�knۃ�G��^���'yճ�E��+��Й?BA�]��~����?a�h�N?�ڧ�L���V���._wq�(2��D�@�~7gz�����`�Y�<(�X|��+���g���^�}�t!C�HM�8 ��$u���?I���{
ق�n�����.�ZӋ6�G��W�!�bm�`�v��b�������<��+�t�@�Ѱ��-V/M�Q��V��:ǮkX�8�"v�_h^lLL��Ex��w9�h��?"�)c������~�j�+�9u�L]1��V9!{_,K���-���0����M���l�.F��P,���]�P���`�@��|>{qx��Mдz6�x2�QX���9�����4su��Eյ�[GJ�L�B���8�0%�Oo[dp��-:��-i����J�GoD]�oag��N���V������ڬ�K, ����2�';.�\<�͔�5c�8m�/���'֤�ȭhک����xO�h�u�>�!�dk;��m�RAH���x��������5y|� ~M����$���2�߿8+~���1lA?$?,=y�E8��6��)����rH�c	x*��2�VqA��C������BV�����;�y�uZ� Jy��Ѩ�#�����C�Ǣ�R�բ�����M�BK: �c�HJ���g�7���j|#�l�O(�A��1�۪�z��4����w|BF"�f���4���/���\L/:�.]\�$���3���6�0�:��m�N�բ
��`K�Í���54%Ь���k�<2���Ĺ*���~}��,�H[w���b��(xzB�<V��XoY=aЀ#�^���_"��f�3�,�U7�@+qP~�rq`M����
�H.g.���	'?Z���)O� ��^���gߕ�7����脏�=?C��/�?�(��q���~$s�qė�U��y���NK�>B�ȑ�wSp��ƿ6�$j��4����<����X��)&�

J���[y�A�&^W���XUOޤ�ITs���b��~h�6��p�M�ND����J�a��$����l�6#����"��+ô�d����-L���YWg���@ݍ^�SB[�|hDB���WP����P��e��W�~���z	ߗ�p5	�TMx��2C�m5�Ď�R�^�@��dR?����s���'iY�
(�p�Q�p�N�$ҙmJQբA�����,D��s񞈁�m��m�E9�@�33)6�Y�F�"c٣�)����`�F�r�`��+������%J"�	 އ�[�3��3�\S��CnK�v�E�2[����Zg��}PKVP]�� ]t��͓�$����X���s��Zv[b��u����RB	G�]G��D}x�3JW/uz9�+m&���H��?���E�yc}^#�7r� ��ѱU4Mg�
��~f��U�oJVaӂ��Ψ��մQ2t�<��V�?с
��v%�)w�8�~V< C龻Fq.-`��N�l�8!�hX�\|�Nd�!�B���]�h���32�����\�����f��]h�:�eq��GDj��e�S]j�V�EX�|�QOLXYծ�Aнh�⊭]!Q�e���}��-X��(����)���dN�'����Y_�	��/ö&�U�V㙼mK�/�1誧���,�<A@Wx�d@�c��p|�z�������k6��w�s��
K�iqZ[�o�qh��}U�[Ð�*2K��6
̥2?�G�}r ����
+�v*E��m�+|�{w*;ӵ��<)4v�II�ۀ�RqM�J�l��X� ��|�ӿ���iY]J�F�Ȃ{cr$uk�D@��}�іS��	L*!t4� ķrE���{�w��IN�[���{�"T:��oSܣD��yا������&oZb�͆sSg^K�UV_N��h-+~���쟳+�o~L��"������:I�ɶ=@�Y G�̡�#6�����纃?��4���1�-`���e!o`J�.n�#�HO
"�w�,(��M�k�b�
��7�\�41�oz�>�'5tj{t��y��m+��9�t���K��K~��
Vٻ6Qi�3e�̿?޻[�YY��j�hB|�����
�L[O[�*R'~���!�k�)�A��M�&ѩ�|����g�G�w�̈
�b��m)N�ȁ�QhK�k;r׼�A��&��@�Ϡ�J���R����n����⍞:\v�0Z�5w������}r���Դ�<2����C/�}Sϙ�kJ�Qk�<�K ݁���ٙ��=,�K�9�"��CD��-y��i�( >�n��������g�7b�'W�<�G'���C�����T�n������L��v�v�zA7O⭇��'p����~ �ǘm�ڬ2��`��.1�o"�.��B�h�g�m<f�X�� s�t�}�RR�@�|S̒�UGg��&�@g=,/3t�݄����L�6Ǵ��:�OQ�"d= ���C������n.���A��L��8�`��3�'��c�xt����)�mN��?�Z�tF�Q��؋��������IY�k��h'�;S���w&A�%2��~9L��	���<�s5/b Y:�S�`�������)I�#^`y��"	&�$r�[<R��;&���Y��l���l� ���\j�H�LLe{g�1j6w���lR���(�q���h�2pw�'0@�f�8���n��*>e�8«�?Hx�R�g%c9<��ȕ�vf�_�C���|���km!�����JF�i�>�#��0��ү�s�.��9�HZ|�F3"�5E��gi��AuSF�m�."�H�K��W��lAّ,��W(@d��~�ݢO`/���¬��@!�Ĵ%�D��K au�)�?�m@�c^�s4f�oDx!N��A�n�z�$��s�#�O "�SA����~)u�8��v����+J@s>��P�"ִ�T�j)��˱'�.^p��T�e|�V��ٻ���M2�����PK?��nV��IlB���:ͺ��+��1�Mu��΀d"ʹ�~̩���ӠfLQ��n7ۨ�g^P���=W��B�BO���z60��Q�����B�n]�����U	~
+�:Y|W6�:�c�s{Vv�o�eԒ8l�&ANgkt���#r�� �F��'3��@��O~XT���3	��q,���m�2L�k^	�`?��E��u7�+���ym���8gS�)S���kL5|��d5����b=hL�=��i�3��bЍ��_}��BXH�Yv@t��R�ph7�c��{�ڀq��Tn�+do��kB/�5���I�g��j`�D����mc���.g�Eڶ�M�N�##D�m@�<jx�v�!O&�鬻��׌ړ���Z�օʡ?z�y�A�]?�4�(���jv����RC3O8لgCHġ�W+&�`?q
�A��M�	�ˀ;�Ɣx�8���{�8��5D$qj���v�It��G�|y����U0�eTDB@�5��޶	����n�H+D�����J
l��b_�^��7� �eޅB)z�I��y�G�9N�uyA$я�_k�z��XC��
�C ؖf1=��"n�9�}��I��s�(^��D�B�y�_�Af��v��
c�H��K�C��ԯ�#��%zҖ���?O�~~�ա�B�l� ���9�
Ⰿ-'�1��R�fn?:L���#��	�{���r�y���W&U@&zXi�xB'p��V��#"�򘚽����7�����b㢱pD�)��wm�=�(LM��N��QZ��-�x���bI����/يUt����)�O������S���9����y�̛X��j�0{�=����Se�[��G z�G���[h�HZ����*���i�D �=T?x�'������M�O�KTA�F}��al#t��*� �X� Re�>���'p��R�!�%��D�d�:�45�Ǆ� ����[�l��U��A>ܱ����y�5G�� �ɻ�#��(�f�'�}z�>�z^H����^R:���Y���� ���G����Q� ?�}�,Y'5��MSJ-:pU���шĽ�}5��L6/B�@U��	c���̝ ��/l倒��i����wѬ���0������1t���X����~�;rm�>�U�mV-����s��t������g�_
r����%��*,� 1�f���f���޺CH��i�|eV�&��m?a@��;[��a��Z'J�o��[��g�N 7��2L�"+!�a�*;��9ZCi���eS	e6"�}�Y�$q��#�%H��.���~#��R��̑*x1ޏh3�.�uS�P]�0�Y���s�9�4)�Zk2v������+�;���Q������;��*�z�-�t
l�Z�7��߯� �lk%���p��ܧ�"�dJ���H����P=*��򓡳�?���W@��IQ\���(J��I��jշ�Q�l"�"vS4��M,��a�@���^�V�W����^~�4}�S�k�����p]/�B�n�$˿d����%T.5� R�̥�Q�͉����`���$�v��Ѓ�E=�����;�cP6QAn#�F5@�yF�ڀ�k��?�q�����	MM������]a�;4�� *3����8?d�G&)�I�z7m����/��+q��I���ySC:�X�N��
�M�]t����^��@����^r	$����l���e1�j�,�4o �|�M��������x������ �X���$?��ۅ0^� �_{ ڙ�ӳ!;e�C'�6�`�Ǒ�Nz���!�C	`�4*b�wBF�(&$c�⃓,pJ�^����DǞ�^���X�XF.'� �c� ���)g�4sH�BW��l��ba84I���a��"��zCwȢʩ;m�һ���0g��8�P���=kL?h7��͒%P��[�"尰i־PG#��uT�`˿������+m�K�D����<U�5N)��<�(���7z�����*´WG�������d�a���&u�U�Hy�J��%r��^��ϧB�E��헠�_e�	�L�ٚ\c�^�(\���0�9Bo���L����sx��>�ֵ1ߏ��&��e3�q�ϒQ�%W��0K�t�]�0����PT�6_�u���޺��(Kxa�� �2`,�唨��{�@x���-:A��1U)=��2v�bw�� �V֊j-l��訲l>��W�zѹ��6DWd<�˚��(OZ�0���s���<����kh�{��SM_�SvJ�d�5�����j\現il �꧞�]�7>�I"�:i���50���d�Af*�/#�4�v��P�b�Yd�������#�*��*�z'�����w� �%�M�����8)�Դ
X�#��D�~�X�'o�����uKSF�3�|�%.�A*/�&�Ԥ�H���Ƒ��M+>.|ⷼ?�Hi��܆��E�A���#��$1�_el��L��G�z�"$��*#h���O�GS�>f\[$��8�G"zZ<�-.b��B�f���܇q�D*�l� �.�h�z�7�X��ʲ�#
�w9�����Z��fY
f����u�@����l��39�L�}Y�b8���������J&��ظ����X����á��j�ōw�g�#�J�e�ϰ��F/U�>v�rk@2�Y۝oE����j��F���;��6K�۪`u���'��q"<)�Pb�f����IU����:���jϡlq/qjs�cx+��̳t��B@\�%}U��yk7�H �:�V�%����3���$�kk�b������\�f���q���X���>���S�E|^�Y��U�G�"O�c��/d?QgM�|gΛ�/21��a��C�amʕ���n��w�-�/�!����<�d�+�+��<+�}Ԭ4L}r{G���l_M'�z��f��PU/�=�aע�W"�[՞�ዥ�%�>�U��%ϗpb��	��!B�`v���@F̮j�o
���i����%��K�Qh&�A﷞��"qDW�uC�����ę�h+qԢ�_-qԷ�0��9�RZ;j8�/��@�%���M�� �}���b�G9z����vI.[���v��ɻ�_h�p���"C������.�P��>������6P�8_fS�U8��ۃ�4s3߇�ϩ�|���㯙�sz9(jd`�(��� �êE)� #y~8�e����*�����OpYFұ�ɽ�B��:���Ct�N��Qٔ&���ܬ.��-B�3u;VF���0AXe|��ô�jj���J�S���l�=By sS��R�������gV��$�5�'3�"��Ti`�����a��j+D�{,pd��Zd�YG�
B�����撮;t
��L`�P��g�~u�4����Vj��˓# ��~+��%2�FrJ��)�~u���;_x&�Y�!�js+����ӳ��jg7���p1C(��XP6*#�a��{�U�57�Q���N�_-���,���I3�-�/9f�� �#��t����Trr���L�����\Gڶ6=r�u����ɥ6r�� ���5�4�U=t[�L��#qBy�+/�UMhi$�:9Sh�J�\U�K��h�E#�������MlDy �#�!0_�/�:�9�~-��R��Q�c�U�ɭ��=�YABZ�+2�Cs�{ٲ���D�a5�.����B��#��P�:h^W�{�/&Jy�S�1����R(����j
�_�0͐fUM�������˝*-��:�M�z!�ͩT��S�K~��]���;�'���KZ�1_}IH�	�Ev`�#�H؋ؖ^-0�����%_��b��h�-�8x�ҍ\���I�]�������P�D���[�,O4V�Y5�H����"5�Ɖ����m�b�WS�Lp���W���o�7`����)J1�����o-�p��5%��d���8�A�$Ceg��n���g�;R4�4����a�G�ސ��:?�����1ܼ?����]ݑH���x#��5�n��VW��&���Kv�$͋���j�5aFO�(^�Ӎj����S�Ra0�:�'Ёrq��ƑBc�e�NS�>�Jÿ��I	�J���E_k����G��9O%LN�ؼ<��kʈ	�܌(Wn�����g�Y0Upy�1+еiO��v���ֹɍt�i�m���ʄDDd*%����?7b�3��8�՟�(';�3I��7�A��R���"���-��'ӭ�B��u>sm7�$w�f��Cwy��W�<b�ɂ�c�a8�kC%O8��R�����ŕ��|�&��"�,d�c�2U��c�au�>���;�.#4�����!6+�oкC�������3`�R]uL�G��������|B� 7'�6.��R�Kzځ��G�T<
�!�z�$h_��C�}�N�9�^���	�&�&��"�P3@ڷY���Ù�����֊�=�X�U��~��W�e*����j�V:�!�T��ԥ�f����fY��[��Ғ�^���zw��z8wy�3��[���0�R꽨y�S���D
�`�­@����}��x��F}M�6K+(����3�H2K�Q�}���4��a'^����a���K)��'� G�=�HF����}0���CXI�(:�myi�+jE
^����mol��D�6gArOޑ"�4%h���sI�.�M��	&�D-tgv���*�M@�!.�ʡ�R���|H�gY�w ?�G"T�T��Mm�z���p���ɋb�������׾���J� ���\l�vp��5��eԤh��p<�4��ӌ�^�ӴK�|����u3(e�ᒳ�wT�u�G���;�_)}�Dͣsݧ^�<=Rq���g��_�Y߱��W֒�f��K�  ���v9V��(�YF
6����7t�9<�7�����0f<+�j�� ��qPI�; �D�%2$����vmdi��v�)��J���w�\v��6�g�a���)����Ѣٳy[.�Qr5�I.�ř�󹏠&�ؽ���f7%�0�r\��0�Xۑ{ 5/����-�������Lǝ�5�T}���i�����>��w3?�����xC�_z,IzE�H�R��|����S��7Wd_N\@~���q��Q05@�!�V� �*��]W�w�6��,TE0v�͙'���RĪ�N�n8��NE��(���ۉ�X�?�6̞�kDQ���at��9��^�Z�؀毺p�[��2:���$5࿞�Vv<=������	J=t̔�]�sN�9����L�Z�Ʃ�����uWi�wr~Wͤf�t�~v�f�h���'_6YV:d����>&W$�d�pZ�;'k���Q(6��k	*��\�]8x��[��bfZE�۠#�]��u���$1��c��$��63��8T�#̓��I�~+������3�*��đ��ȋ�
�X澶��J����0�_2�U���#���lr�����f:gE!Y=^�iw
v@pD��G*D���{�;#k��`{k�!��<���|�h����T0���������g�I<N6<�b�� �ij	�&!l[v��@%����a�2<��`�Q����Q9W�c�[�/���n��fʾ�8�H0$��ݡ�?�_����;�w洊�7�����Y%?�l�i5x�#�n�F b�[�<G����1A�V�F-���������eA�l�:�7aŦTX����s�w���׹�~*6u ������j��؞�@oU�D((���d�8<,+��By�1�[&�]N(�[�CK��mVI��Zk.�VV������Ţ����%�Y��ƀ���<�&��L?�(���^ҥG�7D��?2��@F\�(���,�ZNg�a�F`.�A*66�٦����;�L���d�*�:��I�������g�+�w	n�PƲ5SB���@�����O���֓���p������:�|`'�d���Z��,;�[H�'^C?^?g��9�8���#�m-�6��x��H�����'����
�^��@xX�����l�*�h��z���eaAq�/�]@	�������9�NAO�<9M�&oE�OkTY��� j�oJ?�H�Uh�}P2�&cy��bEA&��X=\����8�4&<ċn�I�6��<��%a��{�|h&Z��{Fe鍋�JnL�W���Ռ�q;s�k�Ȭg�K�w�S)�i�<���q^o�����/�!{��]b8D�V+4�����@i���б�3<�h��Hа����X���qx�K�K�K5�b�R�'R1�����mϋ���cya��ǜ����f ����{ַ�"4+�_W:p�@�p+�,׆H����2=J1Q�}�j}�ɂ���p��G'���Vn��x0ӄ[�ra�R�E(	��b��
����Ȭ���~��'400N�oS`�=��d�����C��j%�h��}'�^�[�r/-��s�y�B�3Xu�zc b� ��p�,'4�JMK��Q�ӎJ�u��1��dװ�z%�w�Uz��3���(�*�S�0�l[9!�r_�m�x�E���%q�ޥ1����+�89�%�.�YU�R���!�$��)&%G"׮�s�2�@�Z�i�(� "����ao�jN�j%>{ UN�gA��0�`�`%ိ�-
9���F"d��0���#���"�*���b�kb�D�� ����m�]4��k��ħ%V�P��V&FQh\�/z{%�hz���ޣ4�C���@2�2�GM
��@(���\8 }� ��������z����� *S(j;���4ȵJ��|XB44H����4��ᓰm�d�ӷrȣ���²���$6m&"�p��ΰ��#����|��_-�l0?Ѷ�&���ß�bZ�-�;5��9�2���X����R�&U��F�sz?�ai�}��I��J�S6��k1�8 �:��z�����r��=�BhPrm��Dّ��?�ZO��`�&�zr�}���03WQ�I���ܟ��I��A[���*\��R1�p��h��.e5�����o�FKl���$��d���*�,����eIB�cg\����؛�?q ��d�n愙�1�/P�\Ӄ�yX_�X��؞������B쭉�NCԮ���&�$�(܁�W��x8�*F\iYCp ��#f��4-xwW���K2*����Q����FB�n�������é�b�w��9�t�{�V�&FH���siށ�X�#�����]B�.�85�� ������!P���/�AEO�[�,���"ߋ�ܢ�KK5r��g�^�'/pY�?e�$ �1�% �͚j��[rSQ)��K1h������b�+:d�����@3HHg+w/�v�F��qΣ��Ky���q���u�8���N��9�d ׃�2L׆~c�"Qho��ׅ�/�U{3F�>��g=�z�o� �:T�|���sa�?��2I��3�1ݸ��uشN<�]z܃�L�S F����ʢ�ҫ+=}�)�:ks��c���rc�Ca��/��k$����HfDI�+� �?%cۦ�1��y`�3K5k6����6�S���;P��>�'��yC�;tIQџ�'��uh�NiJZH�����D�R�	 )�?�q�6F:Q2�9���.�Խ���C��@�������BB�>�42��.�Y��� ���1�t�T�y��T�ڤ���@Xy�ۿC2�l$=�h�����z�.��g�Kv��-��q��pdj�v�{=E�b����T��&�Ɍ��N���࠭PL�W�ytn~��V��}<���0��gNףT>�e	��3���C�2�Z�����<j�XK����F��@�P$BN!O(	�?lt-3���Yaai'���P�`��Sb5YZ�̵�w�pl��?�Dl L%U|)�Ѥ�F?νS�Kr�	$�l�������Y�UN��5�g�B���Y�zհblJ�H�����2�r��拾�����z�x9�Wfy���$�ӥ�	x`�VNpBWYH;x���<�=(Q���GG�B���c���Km�v2yOv�ߔƮ�Fi�~;��md�ϕ�$�B�G��c��<�Ȕ$�X��<��t���ZP<,�k���l�p�}��i��i��?{�2dI����#p	�%YSx�9ҋ��gG-�\�8 S��g�,� �Վ8��e��o�(6F��5�����`����p�7@���C@��wuy4�v�[sB����v_�S����Ȭ����b]!z̽��l)P�<&���`~N�Ky#��E�=��*[�Zގ2��͉2� �Q4��L�����\�n��g��m���i0�E�M�_�*�p�T�h���a��hnm��j�P�tQ����	�vǚ]� �ۀ�jqZ�8`]i�PGEk�@}�zǟ2�O�,a.0!j�>�Q�?6'S�?G��S��\*��3 ��y[�;�Q`����@S�FO�h؁�oufx� X�yD����R���WD��T�WoW�{���-^0r��c�o��ޑ"ym8䚀 �PsɎ;1�<PG��A=e��rL��KվnZl�{�����W
��	�W�˳gW�ן�j�ʠ9-���n���2%�TOP��u��¸3鼡yK�sR�9�Ò�{j�R�}ȶ��Տ���`�24[
���'jw [����!���D.�A�:SE98NP
Q@���G�ygS�h��5�z��5|�R�Jh��n+�ӋKnj�-w�etinq��V3ׂ��uHR�t�Y���s���U��2�-_1Wy����B��N��@�a�q���=��QV ����X��Jo�x�q-ɼ({-vk��u�Q'`��{i3 C?
���s��F-v�T��n���� �>�mwh�<�:�Z,�����j�����ۦ��q�-=g)&Z��b�rٵ�"l=K��������A��̸s;;�}EŞ�v�:�n:��!Na�YS�/��?l ���bG_�dd��W�v�x�I���cc�e�k��5	���Ϲ[rި�����C�!K����H�a,5�������b��k䑎����9�'�	�M�PA��ę�%�+�w�}�$B<��<�Q��p�_b��b�Yg���?�&i@�(��QPH�1pl��7�/ј� 4Ү��R���[~�I7O�n;�i3x=k���,�����w����B��<5n���1��C�!q`A����>ݗi��)K��\]��E��j�}�V�)p�;X�B$�#+�^�>��BBn�Bi�ʻv��d��m�g/�'����5aK����l5�	'B�آ��>#JvqE�j�`_WDFr����X�'�~��?"}/󣉸F�[L����MPHKN��G|p��}�]lT����L^x��9�X%z/�B\]���ZtJǛݘ�!3s�ar܊��{� X H�j�N��m��� �BIW֞��K���n�,��ӌ�H{WT�(�
ŗ���/S���v�]�n���h^��E͝��&v��?��s=��Q�,�ǖP�����5�{�;�yi�tc��E�������(f��A�H�!��i�FL��\n|m��р��D=R�I�툱|~�wN⿓n�'��s����������	���G��k$\KD��XHN89 �:eىJ�?�Tt��Zg��M<���y��xTg�>j��7��pM�ƘЯ���$�JcyS�j��]��uk`Q����Ȳ�C0Y�������<݀0�+��ʚpӡc���JXD[dOOm�� kY�Ώ�lƬ�MfN-��m��/2�>��= zS�<���!�M���|�5w��k/�ZDH��M�9)���b*P����Yأ��ˡ�ɷ���ӊt��� �Ř�H�b)���&��";'qE��h��.��5��?��vxK6"*ONP��6yW��+��nx5Rްڹ�=�8��8Q�Ed !f��<�+lqPG�A7��p���桪�g�+J�-��R��Ә!H�x�f摿����A���0�Ɇ�����A M�^��H����'��7��H����bN{����3�*�$��,�����ʷ�&�ݛX���[!�L���J�c�.���m��PG��%���{��>���e�q&R�K������#�V"Yi��Yg;��P�s[�L��G�Ü`�Y��7�
�"�U��i�#��|��\�B�'��]����^��߳6q���vc�^f[E��.��Wǐ���?n"]�-w�QG\�Ȥ�B���#��T��c�@���m��b�Lq��ƈgck8��tz5��/�U#���Y��A�b��=�� |*�-�o=8u�D�i]���立d�.�˓�⑺Z����e��"u�)���=>�p��3�Hds�Pv:��A�m:Q+�ٛ���s�^[�a^T�%��^�p
kԁ�8O泮Meu����6��_ 8�Q�\^�t	�d�e�\��D׆�tN�U��3yq��P�A���J�*�-� R�<�݄�����R8�	w�`�/�ඎd1Ic� ��s�i�]�~ѳ_o�g� @��o��}-��{E��=bQN�����H^��pp���4 ��}m���$��W�k_���W��	���]>o�Z���hO�3+��i��{�j�P+�%�uRo����e���b����6Xq��៓E/!�Γ�y�ݸr��rf=7&�\Cf)�l`�`pvɗ1ie�!� �� �
��#r����Ћ��'��|�����ӥJ@�"��MLVsj�'�  \̑B�z�!�x��~�i@�6+Zf��?j�I�df<��$�`nQR�x�"�!��hF
W1�K)p��F�h;f��񐡏;��|)#xPv͒c88��.��m����/%u�Ghk@����V9���G�]	���~���k��=�sS� <4�n��m���gs�uÆS	�cn�pm���"pÞ�6�)��a�:��� :�A�ҠI�7�o:��6MJ���LMkݛMrZtH��Z�"3r�M�a�ꎾg��|+�K�/oq^#�c6E�|�@�F^�	sMEh�(� �k�,�%Aa�̨��Rg����d��Zi-�Tܻ�o���T;�*���#҈S����c_?c�昢?�j�T�ޓ�^���WWvf�
��Bʮ�����-�~�l����񀕪P�$��(n?����a(��-M8��T�>���L�xZ�ā:<Q��2��ǰL�S�.V�M�ᅾl�@{�,��cs9+hjc�b��BF����M�ܷPBA�M��~n�?��C����L�-�r����m�>��[K�6t��o�ٹok��B(lup`������Gz�m�^��o��db�3�j���C�%�A=t�/��%�=U��:�ۛ&0&SO@��;�.�QL[�3J�ߙ�\**R��n� 5���n��6Y{�x�=��O:+�Q#z�սŃ�9&X��!T���r�[֡K��B�/��;+��ٺ>·�i�]���������zr�=N�^�@]��L8Sq�������@�xط�X�0iX��JY�nQ��l�� {��	��"�;e�6D�X:*��u�ц:�nf�68�&
m�S���ڱ�,���-�{�2ޝm��`�hf��V�`��x�j�
��I��{�Gx3Y,?Q��e�Z��@m��ǻ0ʨg5�nQ��uV��2*`)(+��&ʲȀ)����#�ʰJ��aA�0�}|R'c��e���X\�u��{b��z�;*��6"ʻ�s��𚷜�Dڿ��Ce��������;o����խ�;eG_BpK�X~�����i&&�=�_�}�Ř��+vN��U����^�,Ŗ��/��y��=4	] W���o����n�Z����Q�
�C$�	�⭼�+3�-��+A�4}��9�	�����I#1�7r���PF�PV�_t@" c�R$Q��b�2M�!aG�8�;jTy�j�����N��}IҒWղ�����//F���K� ��Ti���Qs��ߎ��I�����g�&�a|�a���Emf&C��S�3/C
C�j�h����*�y]!u��HNE���0�d�y���`Gu���fji�7-���낺��C��d|*�����P�����r&^F��RC��^ Y�y��ԋ�Oh���ES�ܒ��v����>���+D�>��.p� d��y������[.�D���^��g@���]���>� ���������9�EUy�t�e��L�=޺�?l��#O�K�q�Y��(�h�4E�D�#FX�˻��<! �Ĺ���̓m��gA�?�W����{��`jTG��.�m�Ngj�K��/MlE�镫<�`��g�.�2o��ԧ1�:,f�o42X6s�<ߴ�ҙX�|�Z�eί�~�����v�ٚ�Ci=�֕���/�X�]b�Dͼ�lQ�l�>�I�bw��<�-�߸��{dk?��٭w�+(1�5k>N��{�j���R���N!m�O}|�t��L�/٩�WV~nc�ww�P��7k�����ό���k9�e�� =�� ó�T�a���_�%|�f��[�ǹ��A=vM�(zly4 0��)�g��n���Q{S�|��gc{`J��|����I��C��
.��#�8,��kѫ���ŗ�Sy悹ev�{�}�0�.M�	qw�Yw�ג����+�b���[m`��PTL}��|-�������n�?��)�Vp��%�ߗ�"H�c=�?S��!"5�+���%w!��d���t���ؔ�0}yHQ#f�����:IHLn��nD�:���G�Z♨)�ס�����[��kf�� ;�SN%�����{���޲��K�����N$�_�a[s|��F�����$�0`&�w{ʼM��2\'���d�響�QO<!�:KWa�N7���^�z,/c�e1=v��I�	2���n,�Ү\���9%b�7��E�������-\�m�ˈ ?$4�9���d�;o`��x�;]O���5>_� ��9C��j�r�*� �1����1��ٜ��k�L������!�L�4���90�C���k�_�K?�g~r����w����pL���U���*-14B����E=��/����x�#F��{� �2�|�~�� Iʶ�J���K$a��cj����	 ��z��&�h���+x�1G��
z�K@��+$z����W~��*��G�%�֦�lgCҲ?�ǘZ�|S�ďSy�E���l��-}�g�'�� V!���'�0�>is� F��bG�.*ٜd��F�W�x� uT/�x���;�h"=�A�,]�d/<H|��ʹ#�Rm�ɦ��q
#�=������q	�g�BF�J,�1��?�AΆ2`�5�i�ɡ�lzDz(�DX�=���.c3t�)�s�����o����g�'��O\�c�\���.݄��K8�z�N��!sw1:՞�ƭ�&���bXu�C��!��Ӏ��B[NPb=2��>�Y<$�%+�M�X��|Ǖ���/Y������f���4a�@�3�H싱�2 �����h���S�X���o|�'�q������_5e��C�G���%��;��􇀥q��� ��ϯ�%���-�2f���tEv����N���@��9k�olH1	��hIJӌEa�P?1ș:n�!��j-���:@I���,S���X[�ˆXF���������$�W{���~�k'���i��RUB��K�ϗql����@�\=� t�����ŢDK�B�~���H'�m���$�#�L�D/�8��͔���73Y#f\��5
�9aC�Kp��opOi$v�;�[qy���L�,a��������1�!E��_���~�I=E:��}w��*t�t�j�)��c���)���ϼvH��?���� MOd���N �x2L��I���0O���i
�Qj��j��ݴ������;��D�B�c��
"�ܧ�e7�~`�[�/�RFK@6z����J(l���O{E�ΤB�R�(H51=�8�qˑ�����In9�����:���.��X�u�"B�{�)�a�Uϋ�����Aghȿzw�s��Q=c�JsD���[�VM
E�>�]
m�XI4�7ܒW�#`5�U�k3W�NH�S
��r�mݚ�ʀ0���2�.tG��&>[�H+�67��J�_.�tI��'8��5�u�NO��:7��,���G(��lQ�}2�@h)���uN�n6߁�?f�<�]6��~�9@f��,8Q��0b�Y�(]_�] ���TS=z�9�K��:�~��ώ{���[���n�e��6�����D?�\��ˑJ^ᆪ@p"F3��w���؟R]
EB��ZP.b����0!l�k34Om���v��*�O45��s"�04��_��#ꅵ:�"&4"����[��>vV���yX����]}8~+~�Q"䝦�,��]�Q��]����#\��?7����r���9��u�L�;S֒��g��RK\*���7��O|� ��ֹ��D㌄�eG���m���.YՋ�m�:��Ps��T�6��%�Ȁ��&�N�N��G�"����!����t6�����S�ނIYd4c��gĿ�fΣ���pT���`�i����{�p4�Q\��K�c�6�8K��~�"� C��Ҷ��Xc�N�4Y�J]+Ɏ�I�ZM�[$����H�0��Q�]�R(:����;-֋�����2�G+Q\��UD��DSf��5�h�TƀI�˾u�A���>�3k�Emps�N7��e���ک�p�}�
ډ����LϪؔ��S��]�޴AԎj)� nKt�P�����3�E!i,�q��� >�����uT�O��H���N���a�#j\^3��R���BN�Dz�*��{��{�u��M�����F��a��;�F��8�i��8O}�8���,v����U���`��z�q��Zqߟ�C�ٖIL���8pQ���x��k����C�uK"��/�9�kq��7��G?כ������<"��z�n�V�D��vvd�!�5�Tjt���U=7Li�A���^/���ь"wP�uDF�5-%��
���<�w0�����A�L���z�MfC)���!L�����ȌfF�ز��\N{��T����U��8����p.�,�X�t�ۓ��U��~��5���}H�����EdKc��Z��
���ddˏ�������N�˲�L9�z<ڻ��ݧR�TÃ�Ey���OM�w�n�Ia�����L9�U��g8��������ٜ{��Q��@ �������� �ڡn��ՑK�ql�31���l�\rr@�E��X��w��N	RϟUz�|\q�V�Dd"'��\��9ꦩ$��6�S@����6-O��Z>]�pu��OEi .�h�)).R
�l^C[�I�l�� f#�#�ф-���^ ���k\#�9^�K�Fd�!���&i�b��C�̭�ߢ;�#rdt�l���8��-@�r�9��ѭ�{���˷@m�F5?� Q��LBD*Dd=3�0A=�8P��色θ6�@'��A��>e����l{J��mT��
�)ۙn[/+����q�'�זv��5�X]e�i�2�6�5��㲬��v�-4��}+����5�]�"���%���nT!�p�?������m��fU�8q��5	�Ψ 0�)zs�˜5�3�l`�lw᱿�b,m����@O�������ZE΢�g���;d����xoFc�N2F'��FѬ��� ��Q��B�2�p��Ǫ
\�`���\��[�I�i�7�m0�rq��fG�M�'��jp�B=�����/��u$���3Y�Cj5τ"t���F�D2Uθ䈵M�誺�I�r�����P\�v�*J �����[�;Du�1݄~
�u@@čg��2j�Ϯ}3�K�-(�͕����m,��f=��RF$Be?i��/q��Yy׊�F�sNE�r+�Z3ԇBP��*:���}����=4����n�҈F{���\X!��V�H��\R3������J��>���OP�@�v�$p���b<�'I�ѳ������x�rf0��e�C�斃�U�����7��	���!ʸ�b�Un��~4����?�V���ս��3�Y�g�
t���ץbz�E�:-qq���{�a�h[��=]	d��u�����7g�+b!���u{eC�T��:�U�Ƈ�re�S��mu�w�h���~��:�o�m�b��~X����nm����K �m,�n����������̾/p&_ܞg9m�í�������+�_I�bJ�d��%j3�~�I~�a�:B4'������(`� ��F'3�P�ƒa��S)G20��ZۮGC��t)�+��ThRcL_��c�r��-�Q�J��kp)+��)���c��h��IXabBEȉKJk��'�k$}_�˖8f�4'��p'���c��[�%�[�%�V���D��L��1=(�e7f�J�ǂ���I��2�8KN���[�K������$gӻ�т��Og���+��׀%?���B`̑R���P}�sQZ�'Md�����x �������Sq�s��t�a�#؞��ڜ�T��$@�)�ޟ�5����q�'
��{�N��(����_&]�KW�Hˇ���lb1r��!	S/#y������S��̨]�m�s�p9@WM��2e`?/*a��%��?����
�pilZAk��v��W�H�'a�3;A@�a�Fo��GDxՑz�I�c���7)ۜ�M���Dc��Q0�:���VC��m�Z��FJV_�f��f��x����6��l'
���״������fZ+(!�\R�ǫ ��<,z?>������_��+��ֲMK2{��;�s�����Mt����5g���Q���hy�e*��`W�:�not$�T��9��|	ЎFbb��ƹ����Zk���jZ��[y)ѣ���,^P'ma�g�I�u:�6�o$3���B��O$4��٘<��:�3*��1 �" Oc�ʜ��`Ze�Ї�D�#��AIx��a�\Վ���~� %��'�a�"M�9��K��gJh̽�²*��c6Y$�%`L �5��>�MQ "߁B#���z�ϣ�V?8���56��Y�����T�{��������A�|#�3�E����#�N�\s)"Hg-M�_~�p2��UI�ұ�YY^�l�����
�,,Y.
@g�Ϻ�vĨ=�8}�R[�h�p�z��z���� �}�,t�I��T�VR�Z���g�OH���q> ����Ǩvq7?�L��Uޛ�Y��Gl�S���'p�;z��w�9�Oi@��6l�h�mo���ѠD �6%��C��Be]�ˤ�R�f۬�FX�]�4��6ÿ�q9�Q���D�'�{ԜCI��Ad�l�l���CK�k��M����������N��rX��H�v�����a��l 
��[X�ǁ;⏦������EO���:�>g�>%�u~�.?��Y�_�ZMX+��^Dc�e^�5.���1�r9�ǆR���>0��Bړ��pGH�� Y�h��e�T�>������۰RѪג|`�BEh�0߭%UCrP�#E",���*p�u	��>:۴����9�J+XԊ��E�7���8NF�K�$�y(�2ll�펅��o�������u�(�U��Ų��!7�⢝k$�`��YDb|Q@kD!��grWT�L�$�X��U|���({Y͕�lQߜ��!��޴�+�k�Ʒ��)����[N(x���NQ9����m�v�k�l�4؊��l�0i��8�;>��"?8b6���1�����Y��]�#-G^�z*��|��R9��&V�:��S�}�0����e#����a�<�|�3z��[��.q�o�D�/�]�J3_,�(z��|��t�b��u�Y�W/Ɍ����X����Yn�[�����AIbN�=�]�;���꨼���Z����>�Ef ;%��W�80��(v�1��+i��`zU�b����/z�8��u��K��b�h���GUɽ���Ң�����:M_n�|'�o��3�zvD��i%f���^�*�L�8|ɟ^mY:�@�5�կ�����l�vz:87a�8��x"�8�2�Y0)5Ȩ����-�R�?sgI�|��:[����)ÿ���U�V�.�"-���Ҋ�y
ƺiy�� ����i9;=�N��l�ǗB^d?��nޖ�b���9�T�Q[z����6KȨ�����?������'%�%�5��^+���Z#2��T���W��v�l첚�<�N}VdJ@0����Q��׉��Q
6F؂T�[��c��8��`�n)o	�������m��������O�Yc�W�����FԈ�����_��Z����Q�ǡ�UZvb�~]v�������¹{Q����^!�y��ګ���~�1�|P/�`���ܴsסǓ>�ҡ�iȾe֥�� ���&�sa��[?y�[c�$P�?�V:�'k2�hp���"�НO����c�S��̄�2J	.������44]WVBs�a��泷ܚ�,7+�1�ʦ����d3=hx�FS���j������'[̃��휕O4�����vOJ+��ߜG+���N�yQ>#_̋�����M����i�Å��qj�7�`��Mfz6�&�M`�+h��~�}�]c��SeK&�ۙõ��3��=�-�U1�sbT�����$^���,���~ui��"�'�3C�2�5D�M�|� Ǭ�r���.��m/C+�ĭF��P�,�&%a6u�-�
���6-�ԫґ�b�P#�^�J��yzF�_I�)NT@��x�[�e����l	�:��r�,�/�3�e_3�Ku&�7NE?~ D�	S&����p}��Z�yz �[��_�@:�=!��-.�Q�J�'��/��d�{w��}ʙ7�lBx>�-���\����-(f�o�+(��XM���������(B�𞝓���3x瑊_�����ϊ����,Z�k�C�]�~)%Y��
�/�~�I5#/�m���y.�5�r�t�z��8�� n���E����JHu7|m2bN�${&�%?1����[\ـ�C�9M=ɎQQ��+r@{��}Jh�8�
���~��A�d���!�1��ۇ�|ځ��ϛ���#��T깱�\��[N"b������߀�.x�D���˟����
MnR1&�� ��Z�3U��P�r�X��|\��/��3!����3rFa���}A�~c�^1Q�q4�="�K�*۬�?!�C��Ӈ~}�-���R�FN���*=�� ��Q��ز�$�u�I)k���v���Xo p���:	R�=���f�����Y��ܚE�59�P �?:���%O��M����������^7��_B���B2E
����-K�T����*�hMP!��5��{˜�."#$'�O]`�ki��b��`��ⶬu�������UB��r��g�d��J�����~d~\۶q�Բ/�{C�J6��5�L%�d���m��ثʼ�K�m�������&��|&]��p�~o���pV"� s����V �9�J֍O��gohkxR� �?8j4�?weJ�7���!�x�E	�����ۧ�8lB���n�F�cˇ������V��	��7��֐%���g��U����T*N�aٕѝ�(
�c&s��j!P��#���uC��O����3�@���ћHo�;ta�)��J �`5k�J�5�.o2Mju#�=$�<��Λ�$����Ч-�U�9>͕^ⵖ����l��aJҞ���zt�"7\b�q%$�D;�ܠ���ZV'�ޡ�.A�z���z���d �U�����*7�Md����oh�W���O#�#��_���k�ȍ A�����W�($)��'P�������H��B��/ٱ��k���#_���f2:����K�;��/͌�=�E(�j�g�+�Q�bD��}^Y�r/E¸E}]��բC���L�f^&n1uJ�	*u�(k��Vl��B�Giꉚ}X䌬�˝]Z�-2��D�Zr�92V�mݹ h��O?8:���BB���Q'l}�THWZd���SJ��Īrc�5c�o�ޏL�h�_����V���]���_h�t�$+'�Ժ�=L�ټ�)���8�cwl&}[O�T\?;�v�݃��kl�z�c)p5�)k˧14�Ō����O1ck��8�*�M%�o�jn%�1%�b+���ܯYUb�}�U}?!@�j��~Ւi;!˵��W��RM�u���#�K�<�U�xOG��7���h�Ut�!]�4x
_A�3��&��)�O'y�E!�c".���r~��a��94�?!��t���U�X=
�~ sid��,\�l�ck�ߋ�9��[\x,��,���u3���Z�ĀO�=j��j&�S����G���nv�O�u��%`���P�ibw+��k�S�����'�z�蝊��������u�xE�����VQYd�����iˏ��z+��Ms��(G��0C����}�y�u�Xg�[�N/҆��[aKɉxSG�U�`���E��=*Aw1�����Ϊp!H��������%y5=�:�4��6Vrݹy��&���N�[���Ͻ����,'Qգ&
WO� ~�7����Vh�v����5�KS9�>Y}��I��J���,?`eY!m�#�uc�X�/���o��%�D��v莭�ѱYVɁ�n��V�Q�ς��q�1s�1Ͻw�<�Oł�VT�)�u���Wm�����f�������U}���Ѕ��e�3�i�o�o�!�i�}��|�I��q�7u�%��{���wN����4-`{BW�4W�-.!E�o�gf=*�_����<%{a��� 簻�g<(=Ě��18K���au�iG0��
��+��� �N�R�}^Д³aC��S=���̻�T�gU#��;^�j֍r�\��L�����.�ρO8܆�S%g���/b�?^��T����@hT��<�a�R��u�SD��_��?R>j�Y=^���P�@��z/5�*4��Ήk(x
e7��g�c'�^��ɃY
{��(�H��.����->��X�d��<1>p��\�G�ܮօn|�:�ysCWI�0ݚ�I����[��E����9;� "ʯ�՝N)Rqf���,h��uM� ���X��zcŵF�Y�I���k��a�ۭ�b+&V9I�rќ�L��~2����!��7�+]8�0=�ǲ70���=�J��.��0����_�i�>v]+�hR�v��#��(���VvGt����?l���:Wo��MMQ��pQuz\���	(��B&�!ƝQn��*�w�?2p '^_�59�a����� ��1۷A X^�.�$�f�j��x�00��.7��L�0���~���z��ܙ�92Ai�wYL�V����~��1Y��r3�T���6�.�ߜ�,D�2������}\��U����{�4�	v{�7��5z��]"�˕�H�Z�tƱH3�؁��$�`�p˅a����*�	
�y��g?�zf�/ִc:K���+WO��a�����du�7��W�#-<�] {��x�(��;悈�<fs�'�b�x����r/߁�=o56�q͚\W��'7�I�+�3C$����K�1�b&��+]��}Cs��J��C��wAu?�+L{+����q,��EAov���(R�S��,-���~ےҩ�앜|_~%K�{h���џ�3�>r����q�%�!�s�tQ���
,[�u�`����4��B��d��%I�/���z��zz�5:%�ȗsã�Ov��>U0��j�_y��|���|�)���7n*�5᧊�;��ߔ���`�F�81*ͦ�0���tɍ�\J,��ޣà�1�C[H�̊�n6��zX��j�q��JI#s��3A��m���� koW!�kp��njn��J�煑)f0��������j�X�=/
7��F�$mc�O���c"r��Mh9�U��G B]���u;Es_Z�=
36�%]�bUM0%��8��F���(���8���Aq���!�b�C�$-�B���p��:����r�9�c�H�"B?�/Z�q��y�L�����.���p����E[D��Bת�r��t�Z�r;�:|�::gs��f�u�*����r'x��\3/�*�b�ݒkm,=�A���R�#���2�5a�c�K~$u�'�Z�����#3�˷��f�!.��*�Y���L?#w98T�V��%�]<R��й838Q��e�
��1�����
�������I�M�� <���I`B�����6�����w���)�hxxs�y����Ƥd��X3-E����،����`��9?��~�	)8%�����f"� 8H�����D�DƦ������7���ʪ��ͷ�BƋ��E���Ut$ ��CF��p&�z�[k��{��]Ocw`�.��2�4$���ddFų��!�X��t�rv �0�,���m�$=�n�w��1��A��O�;`���<
�Š�j�y��aD�EK �k��j�3�.�5q�y�p,D�g	s3�3��]+3ӯ�ie�0�E� ���kce�������S�s�%���r�F�}��	�O0�2��VN��8�?����S{���~1�Iу��t4��o�A��v}�0���D�U��:(���G�T��M�T�S?��e<H�ŀ����ӡP�vW��.Q��.y�����_r������я(T�	�A��Y�JR�s�VJ�H`�h9�k�2#'k�8U�#sLX�\�6�=h�Nd��x�i�����^���*$`$��s<���οH<%��Rn��H�xr�R����663����d��������L����}��g���6�e�[YI����	�@�R��2��G����[��=�^V𕜼�v�67ROr�����'�[������n�{V�!����'hv�U
����0�	Tyt���Ӫ+ ���
�4�kZ��j<�c��_��N����v2�΢9�*.>�c>T�5 .]��h >?�z0q)��,�Бq͕��l��"�taxM�O[G��Hq����I�V/Y�=���K�^@^Q��V$�$A�c
��J���sY�#,�2 �����g��zR �]�W�1��r��R��q��N5ݧ\G�e-�>A�̿�[� ��0*����i���46��M���#�*�����4�6�d�j�&4T���e��Ezv���O�K��Q��<��	�zx��T�;�it��c��Au�����P�z�2W��r`8B��J��|�Y$��4��J����*��9� ��P���o�x��j�5N(�Z�i]��X27lIv�j:YZ�o3������>��O��yܕ��U����2����b��K�uB6َpa)�gt��������p/,`���?�B�:c�u�}��z��)%SJ�	�I�ͮr��i��G;C���܁(2�q�Db��zT�r����[oO�c�p��#6�CU?1&�gR]�>�w$�Nd�dnTb�4��:�	�+�D
d�����q�����b����J8o :�L��Z>p���r�`}w�l٬�(720�<��f���L^�z��"osƩ�Lޓ8�rH�F0l�s� FP�M�k���;ΆC��
|��3�d��^.�,�G�M>���1��`@o���>pV���%a����[�S�[h�AԊ���_':+��AӼ��� ����e�/�`]�^���N�\.���r;M�L��[J�֦���������h��kj���]m��tS`,W��������3
G�1�/�Z�{�)��挙�t���o-N���)���ac(�YB�1\�F�ns�t�<R}�1o����kG5ݤ�`y�����fR��j��L�������#���
Zڧ��\h��J�̍��(�I��V�5������4�V(~�^S�����l�&_r@�V�w����� Yy!���%Ei��FS,A���G��
�œ��L�*��n�FS7�PF�p���g����l�d�S@����~��W���G
tE��&�i:�<^e�J�?��f�/a�����a�ZQi|�s���0�>��E>�h�F�%]�Av�%�o �e��z��6�@�m��L6/�����_9�r��'�́{�^�fS����3�)�S���*ܥr���.�X.m�#����<៥�:��Y�;;�6�铖=�P��ֿ���L}���یڍ���8�
�|����������%�ªP47�;����s#��KeS���SHkܗt�C)��	�J�LVUZ���,�2�t
*;��l�`E7�II��Y��G�g����|����ֲ�I��M���n���U�d���:�X�/ t�߅ۊ#f�l|b|k/�j�ߍ���ECQ�4��\�s�<d��Ky�:2o������k@��Q����-���/�U���=g:X����Ё���V
,��zy���
+4��"�?d�R�a�%���4�=ڢ��e7�X}8Ƽj�Ea���:���)]eЅ%��_�eY	��|��3]D�[����x<�3m%�?�����1�,_�8=8�q�s�VCؑUg��F�u[Db���W:2}�EEoX��[-6�3����!�䖀ڈ��}�.��-Y �l�6V{�+@4?��ZE��\����g�C��d���3�&�(��4g�(0"�.;V/<W/�ى�s�e�Q]F*�a9�nơ��׀�
���'koGpY�;�?�<��C>4�sS�B���6	SD�����<5�A�Z�E�ϓ���3g�p�FjLUE��I������-���Kҵ� ��
���%-�Nn��4����\�=͖�[v#����CF�|90θ;��sr��=]���P���vh+��{)���z6V���i[��#t��i��G�V��VE�\9���Ls'�v����~���� R�_n�LlN*������]�@��1W�>��EM�(i�Zv��>�k����� 7��*Ne��z��tI0Lڷ�4�w�מ�`���Zr���uS�e��*�A�d]�Cd:�xX2��q<�&R�@��������S_�
/�/�$%/+/����i�\����^������	8�T67����;�e�_�k`-����*�3�h	�������Ta�ת�p���H�+���$�3��&t-%ZK]9�~�ߏ��Sѝ�5���vC����Ae��İ����hj4/�4��`P*j	�&1�c��T%�H�W��N�����$!�7�??�)��f�P���H]��1G�SL���R �s��_���-?���&k��2:P����e�c|ڜ��@��sa{)D�8H�W!�M0���Ϊ��w�/�m�+��cf&�3`+@~"�Ы�=�7�a*�����HyBR�m�?JB����}AM�V�݄�0~�E6\�!sN�Qv�kɭXNv���#�������(�aF!U��<pa���i�O������.i�n���-P��} 3g у~�#N��+���ni�1b=�����C�����&]�J��9hUK%V�LsЌ,��Z�(��A��P���E�3H���w �!v��y�*��a�&���grk�1�LY��7�%��e=���A��Ҫ�ڂ2�c�}�c�k�g�a�����\TH<r�\b��כg�n�z�w�_��w�9�"B��4`���6#�J�l��s��a�b9Y]��m��^�;Oly���Y�󤸷"w��#�ϥ&�֍�w �uZ4��7C�0DA��1���:]�od>�T8�>�NoE���\S��X����l:S	�&Z�v�����&1zƕ(j�/��/A��.-~U�s��6A��rkT���8�k�.M�4z�;`�S��R� ��dևWB����&O;ⶸ
��(���drG9� �S����2�Ff���l�8w~����T'm\��z�~-�F�~�G"����CB�|Gw��/�y������at'>��G��̊4u@�#d���%o��&�U���7���N8��� ��yr��	�o�)
��%WLn��}�wKQ��LW{�ci��OR��,]v�i`��&yV�Cd���2�Ң�2d�o�D�x�:1�r;�7
�U@b*���F���r��]���5�o\��oN\;��]���%�Y�]>ݼX��К����]��wO �2�uz�/S��F��D�00f� X� ��%���DJ@����Q���-�yA~h�H�=i;�aJ���TNC&�S1G@O1���2OK�H4��,c\�L!���a�=�������y�X��³Y�n��x�Y�|H��˔���"* 7y=
�߻��������_a���t���f?�̊�aue*��.DF�( �y��[f��u�͔*�mU:MV4���-�S4so�Ţ�8����߅���T� ]�~�E�Ӷ�+��;�!���-C�&$13�*<˗����ȟ3ӟ�X-Uү�j�G� ϒ�dᯐS��M���� ʹz�՞]ٯ�l@���Y2%����TL$�YRz/7_ 'ߧ��C��U����_/�SՃ��}��s*~6Y���#;�1u������#������*t��#�⭫�>����1��%�C��������e����#{�J;\��tY G��g�/�a�Ұ�����1G�,o��!b
'o	tZY�U��� ų6�	��k���*�c�ϸ���؝����yO3�b���*u�=�DIh���kT��+I��:Hl��TB�-	Bz��~�Y��A9l0�����y�)�	���y8��."��[pr�L��`��������W�A�O�1��kl�d��2I��A�g�S����Rΐ�����ٴ��n���O��J�Ʀ�u3i�5X���L����O6`p�1%�����7��CǨ�=8\u/��$,Azb{�(�d	�#�ԋ5q=u1Z%?��~�'s��@ ����%��.,�n�[������t�!Բ��0�r��fa�y�$����@��ܢ����Fk�'/D�[��$�u*|x�,�7��
/T�9�D��R�*�Fv�"F��j��a�hS.���z��T��g�GgQr�zX��HK����#2�m���$�9��։��o��A�(0g�Rb*:��Yk�)ٚ��X�:?+A~�VG�&nw��5s�a�1�첩I��|�Sբ�b�Dg��"�4��8����Z����o�en�y?o�����N�g����-�b��Ӱp#Bnj(
Q �G���%-r	�gdW�Y�]�$�*��0��qsnB��1�I��r�"f\�~��&�
-��욗�i���D�ņ;e�Y�udL��zVh�U�8B�6����|�c���`�K	�1M(
� ��J�m냋|4h@�;�!y�K��(X ˤ���� �>�iatA���U��q�͵���~W�|L���̓ty��o>nw��<�s�_�"�����U@����<�����-���rC�˱�Lf�G�XW�[1�:�a�����y�8�1=�ԅ���-uh�B��l%'S��Ct����D�rq��3�^Ł�ֹ�����uPk��7_�7�ؑ,�6���/y���ŭ�Wk��G��9��rz8rq109|U�^It���b�g�t �*=�@I~ԞgPO�&;����	���=�Z�~iW�'~E�����_,���`[ku��1 /ُ�+��zk�,�$�mG��H�m��!z���2%�l6;l��;�q�#�Z:"�\�O�&,�N�	#A�I�'V�wI�ox�����\���^�ݷ�%��=r˾\�?�%�#�e�h�L��"RZ\��[�I@�jE�]j6!)ٛ�-��-bX "��ul��[�L�Z��Q���v���� &�~s��9���f�h�L�1�b'���L�b��+������7:�Shlu�f.��IR�q:N�L@���{Dr4�l��)��)~<��@��޿*��ӒX&֋+�I���0c�fm�p;����Ng��X���x��t���^?6���geӁ���/yVA��=/pGg��������&CZD�6N��/�������G��18(�/�Z?G)�*�N(ʕ^���ņ��v�]�9�W�;�=]$���߶�^Ҿ����k��.�|���CN�φ�5>�7�0�1̦���+������k����)���]��˖� Z�V'T�J��n&�S�0	��E����W�L�j1��O0�~��f�_�&1ʿB�*��mzP����j����\g`q_�j?����;4�,+��[��T�ӅbKT���ܞ��� 1Q��-6s��I�4|�l;#T�M��i���'��ьzazVI��U�J��2U��8ɕ�Kr@�\��X+8��C���`]/��3�}9CE�"�������Z�
oF�S�=vSQ��3.����超#�KJ��5�n��#��%���O����r����l'kHIF�4a_�D<����&�Ix�4%o}t���m~#���#�T��Tdp.T���J[,d�\�'�jC19��l(z�ǘ�R
��8�$ϳ��77�l�˫�n��Ѣ�>��-Lʫ(��N���Ȭ�����7�7�V+�1
1��,��}�#�D���½U�Zl1n���ߔ !c|C|�m _�S|H�w�_M��I����3��w|�ԟ����T��q!t������\q�2��J�+��Jg��'�D}Hѳ���q�p�*@J xn�=�BU���l7TȞ���Rb��b�P}��9!��E�5���cf�xNa�oo����F���MW'O2(,�e��`����.�Jci�q"%��;V:�>�8Tb�Ԣ��(Z��2�e6=	,���ț&;��9
����R�f^\��^�zRtF%�����L�b�Rs%��:�]�?؟Z>>j�u�@c�����d��G;)_|�$���"���Չ�2?�y���S�0&�B�c��Γ��zK���m�oyVj���}������'��Zlgţl���Li�C.�
��w��T,�#�ѭF
��|�[CS�c<*�jbN".��^�����@��xe�1xK�S܋LŰBa�=�2M�w}|����o�'��.8��q��j�D�4�c.��F�0�x/�/��!
J�dT��0�d��:�[�)��D��g�]��]��[��J����C-�P9"�k3Z�I�'� ��f�;Ӕ}�ʎ���V��q	��^��c3�8��ʉ4�#��@��.�L 0����G�Dzρ�P�<�ά@r���vz������˗�����qF�}��2\�j��;��mQ��,ٞlW�E����}��"8L�yn_��u��01|ƔC�О
_# ���1�K�$ॉ�p-K�m�*��s��[�YC9媖�/����ʣ�)l۠�x��_��A5�w	��
�7˗݀ы~@�
_�Pa�{N��S�b���V��m�̩�V��T(�4�e|��\�|�Q,�X��5���� x���]�,�w������&m첵�N
P�9<�F��vL�>Uw��1V�y��>lQ��C����Q��L��8gWV_�cRVL���2�\�ܨ�!?(�{:A���I)���f8ܤ?��!$MfL��o���Xо54%-�:Wj�%h�ͶE-`�)(��1߄��s�E'�,Ƃ}2^Q�ts���~�/��E������"H튗�K�P�"�'~/�����_M��p*��;+�?	������.C��ciqǘ$��w��H�����i��9����Mj��8�Z?�i�;�寨
8/�Z��ޱÛ|��q 0YN	,��hU#k�zs�����X�]�j���Lb)�' xeU+�-e�v�i�D�%�6��nM��f6d�0�D�|'�k�p�L׷h_��<�}S���UY&?#~E��L�2­���Y7�`,3�9/N�fK:�T���ޜ�-
�*]���j9�YK��[hw�t��PϢ�t��G��o������*���K�mE�%�V���<�'N�����v�=9���9��r�a�0�8HgÄ���,���R� �>�������[�� M�n������M� �Q�K���g�����/I��C�!�$���U0,B
�$^�������Y��ΥyDi&��r�>��
�]6��2ˇ`4��	wæ�IQ�{��5��3�yI��?y=�����>��_BL�?bE�.
�SOz��z4|�j�i�FL�?�$�:��� ��|���^9��Et��~���d0Ǥ�lk��N�]w��,���w��b�sU��m�ta��!�.��"sr6�Ī4%=wtAqr�E���qBl����T���G��s��g֊�k����YAOf�~��L|������|�p1WX�N7�f��S���I^�u��<\L��Iag�y�������y3p3���0�$�vׂŕ�š����aLRWm���D�.�s�lKד�l�V!�{���8J�-+͊�/J���6!��J0��Q }�5���xc0sq���"����^d��s�-��	4� F[ �ĥ=j�3��-��yX�%$���x<�@�=3b���j�b�k,-M�\}�s��(A�{�a�Wbj(���l���-�+��WG
?�*�2�"�f:ޙK���I"�����:���%0?i[Ĉ���Z&a���=&����,+������N�9�mTDߒ
٧f��$��Y{9V�$
��G^!��1��#z�A,�uǻw��`s�qF~pN�
Y�x�������'��U��l�%{E�J�H�^-u�D]���!To�H搸C��(B�=��(��2$�>���_�8��,�-��VW�b�?���nc�_U��5��I�c�0�dsO�~@U�� W}�eQ8����KG�������k�Q`����d����]jD]��T����n��7��:��Y���ac��V�0OFl���	֊8sb!���N��B�\���*��\:su�˺���sH߭����2[K�Z\q�����nD���{��c�+��J�)�� Be(q��f��B���Y�M�<���]��-�&��{�� 
;歌C��8�J��T>[t�+Gc����!��&\�9������N��ot4ҿ��A�f��g�!_H��EKC��P��N���Xp<)�����C?/\;Z��\�ĕ���2�42�Lx�b��l��P�cyr8S_��׿7�tV��6���E��� �T5<.�ge��%}W(*�����e.Q�'���N���6�_
~=6уfy�i���P�,��&�� ]���������hZ��]�N��xu/{1?Hk��P�Z���Ǧ�gj���W�(���#��T���w����ư����/�n�RŃ��#G-�R��ڟ��c�PWא|4�y���#>`~�ݝD�K��;^p'�~���c�Ho뷲�ӑ�N'� 3����9�p�<��ԫ�۪�'��@ؠ�����gc���,R�a�M�_�S�+�cȫS�������a\�y��,Xm��D���gc����0�5錴(���f��h��D�v.�Ba��R���>����������5�$�.�r���#�R��r6����.XQ���"�;��2؊���Wyn棡kp~����,Kes�#Ch�@L�?`������22;1����z��x|`OE�W&�e�W���-���A���=��NsfB���x��$�66B���&dh� �ojj1�'*$�J܃|�t�Z:�(�g�j �$PW+��A�.E&K��{�Ca�C_sf���t�~��AA��K4�[R�vF8����L��� �f�6a;��č��L����1��ϙ�����ב��s|�P #�݋;l�ZL���xl��t �c(+֝�CATІ���m~��5T`�[ῐ>M]y�W3�|�A|M5o�	i)����v�a�%�Rʡ�;A�9�+˸���;�����j7�^�}��SA�q�Ϛ+���_�-�8�x���=e�ch���$�~|v,tG����v- ��"e�6m�gX�B��Yqߪ��D<������\�b�`hYg�LyTz�j�8_�A����P ��E�/b��$ /ؠ~ {�
��V4���L�V[�ICl�G�7d�DD�4��C�� ���ID�b���i���)�j�9-�(�[���-
9M���)^��{L>h�l5��C��K!���c����0y~k���a�ў�C���؀�a����f�[C�y��s��p%����;j�9�x��
���F�oB]!�!�F۫��4�0tq:ϭ��4;�!�?/Cd�w�v�c`�Z�r�jp�n� Tr�5)}[�&ﶒ^��^ȸn3"�� ����C����ak%]�a":��I��� �:�E|�ˑBP�y)����r~���T�M��>�Op���u:w�Y�[̫=t��+PM��d�m��3��P���rQ#q���Վ��@ǬL��o� �S"C�3�8o�����w?c����Z�a��2(���H �褟\�����L2&Ȅ;2̈����Qf�$�?����A_�޿��d���r�"��F�SI��+9;F�"��i�g�kmʹz,�sdP#5d]�_WPH��{�p����*�h�S �'�2���1�_����w��� R)ze�L�G��dV��\&#�\��pS�*߱���%�X�r)�`���}?T~/Z�� {@�\�ر1C48�f�S�4J������jg�ʬ�2�����[��?���[��_�?�p�v.����}�Ґe�Q�)�����gw#B͐�3�_B�0E��fzA�fAQ�A�{"i���S��-:ԓz[����I�;ƕ�8H���6}��j��9�*���=�H	L�dB�VK���~��x����/�e�so23��y��͂�3�$DNڞ�f�Zz�7�T�	K�mƯX�R.�b�����Ir��];g2�8μb�m�?�z+g�Y�x��同� x0�}�2�d$p�F,A4UϬ1���u}�HUx,,竒r��N�~��1��(��w��NPB�T��dK�2�4��P3{<�͘��>R����o�w��.�$�e�'�TRG넭��E~A�Ą�����w�S����B�5��ϟ����敵���.��ֱ�=δ�q~#����[�P��Gyb�4T�������sچ�^b�&��7�+��#��7}��-C��h��xc��*k&i�A�;�R�3���I�ث�1�ʩ?�C]�j�x�ϼs�MW�3��{a�:S*2�	�݌0l ��iK�/�b1;2m9�氬[.@7�lbD�|�.�k�m��
z�3��e��5��-6d��_+����A��<���{V��Zd���dx�g���R�<3��t���}�Ygi����eF��ʾ��gco7Swߩ�8o���9��2��l��y��:R ��y��V��0wpO�V���e�0j�A[B�4c�"o^o��q�s��Tx6u
�d���k���}�"�udΠ0<���иTw0[�i2�mp�I	�0.��%�(�����m[�D =%��>7>��x���Ƙj"LL��E������;)�]�%'��#j��p6�]:zV���\ܡnf���}��P���p�l3Z�ܙ#���n��[���B��̓ˍ��b�z�_:͈D'�g�L)vO�-�FT�@1��.c�/\9��Af��f�ɨ�N"N���S��Gj����ѷ��%�a�49�މP��B�ȵx���=���*W^^FA���JY�4�d5J�~@2�x<�:�k:m/�[�$�q�z��h�����"�#���Nr��i�
��v�&��Q���1kA]T���\���I�WOլ��7"I�QN+ O����}��B!;w�oYYq=�wwP`�o��$�e�����W��d2(1�^��*�9s�9�G�6�=�w���a������j�ǜB�i�vt��$��=������# >W�pݛ�&!
�v��װ��/��C�7*�d.�=��=�~1%i?��m��(�}g�L�Ų!+N��cq���؋�YO��'F�\��sS^t�5��ɀ<~�`S�g|DOmo:b���{�C*'ߐ(]WQpn�$��L��b0[.8N̈�'�*k� ��ɰ�n��mM�<���~��h8���/�йr�OphS������/S�ȩ�w�r.�E�FQ+	�B�C��}ll���5��2a��Q��
W�b7�O:��:*@�\��T���2{aϴ�!��C�C��R�L&W
�����F�Y+�SH�JWa�ا��>#��t쌼��5n��U���@��gT������\]���8�u\N@H�@��W4��@j �BΠ����{�NwA�%��vB)~j��J�5%{->��#<�H��uv�1���Q�6�c��]��Q(V��do���P�������)�8�R�-O�e����rG��h<�3��[Fb�w_F�V�j�hz�:-��ޕ��h&Y�6���d]���rh�2wN�׭ƥ�zAo�O�kW���|Em9�7sw����3���?Q��-|*;H�}�*�����BO1�X��D����Z�M��'��-�� -ȁ2[8�x��P�ٛ�Wf� ���tNz]V�\�7 m�c�ߤz%܉Yq�6#��n83�7L�\�T
hl'E�V^�Ǡ��8�G�s�'�\�����n)��Eτ��g@h�]�������)_e���dj�z�2���D�Y�n�����u8��(�W%���d��6p.�#�,hrڿ�<'���Iɑ��I��V�M�aSHMOK˕f��ܜW�=
�;n��_�Ƣф���4���ވ�1�j���%�f;dϤ��q�EM�$�R;rK�!������&~��D( e¶T��yt��!g_���Z�h��Y����CH3ħs~���}%6�D&��,��p`�RnT�[��P1Z=����)���s�������l<�(��"!�ŜTd3o�(��XN�;N����]R��`��:� �K�v��������7ٴ.=Ek���o��cң|ޒ�:!t�v$Ih��[�S�M���F���#�3�Yh��������0��6���_���D��^{��9QW�K�	Q8��ؖi�A���\���1:�J�DX�B&�:�09r[{�q$��R�\7��g6�2�M��nT�@���m��A��x����v�E9d�4htY�,O��9��;��]v��rD���~8������-����4
a�W�k֢�O�7�Q��D�3m�xq���m+}&R��z��3v]S`V<�Ѳ�Ր�t	�}㏥�9�sɛ��OF%*?9�m�k����:w0��w�[d�n�������6]hr��<Յ<-��`BT
��+.t2�\�7<x�F50�q�u2jE�J���"ɩS�zT"c-UB�tI��:���_sG�Z�e�'�Ig������F�3E�FN�+M�vn�%�g��%~�SUQ ֌��6���T5BN�)��$-_2������b��;�t��7�q �{�Y�t��g���
ϾEj�0���h��|��Gw�TM7~D3)���2�k���l���}��udeT�)�-�@��ԧ&�f�R����B����+|�@W��8x5�3�8�վC���#N���_�oY�e3Q�F�r�9�sWc�Η�?�}�4��������",#ڿQ���Gw����P�h M���'z�'E�����̀��E�ҕ�G��C���8��9��Q�L����8�����*��d=�h+���dE�G|V}��(�dq�	ƹ�*�_ع����zM�_h������Z+�Gt�E�p����M����e��5>Z��t�WV�# �&{đ�s��/k)Z��K��d��_�M�`�q��r(�dM����~D�����hd0z�*�s{����@���9�oh>g��=������(�1�Z]�m��	�׆T�"	�6���Agc��efm���7��-�8[׬��R)(��9�ľ!���U���������S��ґ��Z��/~��������?�ż�HT�:��H����4:��}���D%���N�?��K�?�k�	���6+)\�I��9HO�a��u6ߵ��u4�=I!ZA�do�ar[��kkd�L/��px�\z���Q�Y2=^��%S�ؚ3�����$��X������Q�s�.1�1�w0h�-Z���L����6w�X��aڥ�~�����C$d򾋿Hc¢4��R!<vm�r��0����qև\��<�9�/2K��LXBr�DP���0�odw@S���ؠ,iOZx�"��p~M��������\�a�|�K߳��%yP�+	*B��(���ܚy���		�U�lj}�!<:�遍��Uãu.��XJ>R>�0�1k����d��F.��l@�%�~�1p
��0��`>ƒ:'��y� �K^O�69-Q~�VX�d7��.Ѿ�o Lg%,`�c���L<�Q��oH��xVC����|l
��0����L	���nd}�K�ƍ��	[V�¢�G��^�QG,��8��k_!s��O�N����Zq,����:� h�ŧA�F������}YR׌27������z_���F g1��>���h훑�	C.������A��-q�`g|�W��I�$���A�Y~t{��6W��92����hU���?&o3�M�{��\�R��\b����bn���-l��CB��H�{�*�a�~���~����^��*qR�����!/�l�wwa�!���2(/\��N�e�G>��S����G�=ښ����<+��5N0iu��x�#w�y���џ���P�����j1�Q��-+��Z�qJ�p� /��TQ������m�Җ�h 1#f��#A�9#�/�K���*_N��
��W�w����@V����<�=$Z�%�b�+<�:�F�Ֆ�X�D�M5��$MS��a1�5@���Wʉ�]
]�P���Y�9��FT4�^,�(�٬��������!1�p=VO2�H�;p�l�`톒E+cb?2��[�h$*#��֕܄�Q��!�G54]�>J`_�1 >��.�Ri�.�Y� "s����T8<v�F�;���=a�BgF����DQ��-�*/�����#3����I���U���R�K�o��d�Q}Z��E#��Bf*��ZY�r�F�t4�����0�k��K�������u�)h�8-[&j����@	8�6�cg��0D�ED#�?��2au���"����9\�;��K���$��[p�)֍ʮ�����M�G�;�+�q7��w�Xm�.Yу6�"W��3�9�o��M�%�Y�*��Ҧ�*��L�9��(|=4K�O�8@��S"���}5%@b�slJS?�p�HQ3V�ՙ�[�0�#�#��M�-f�8��+Ye��G	\1�L�t��N6��S��o����\��؞@�\�Ԓ�L9��/A�Ga
˨@e�	����s�8�K-�
�;1��B%���Ϭʔ����G͹IƓ>i2����B^(����&��tk��[h*g�8Y�E���.�J@��F\x�3��ЅIs ���U����5���iIz�:!���0F;��55'�h*����D1cA\�v��׫[��݈�rܡ�G�0��M�/wi!6�!i�ڿM�$j����8���ۤi	K��,�-c6�W�i�V3�Gh@��9��4ٽ�lu�����F�P/�>W}�������K|s�����
��X�2��ˋG&~:�+:�@�c���0�F�H���؛�mf�on��tnO=�Q��?ϛ�b���3@t�^:��/�C�
�g6W�ұ��B!�L�.X�:.I�� �X���L�v�ǹJ��Y���0_Ϯ�Щ�Qh�6�w�s3%3RE�[�1�(=��g9����e��o@�{�P?�Q%�}��U_	�mF�����X�i���/����I��祊�V^��zs��~|��Z���v�奙��&û&2aw�"�@οo�P�e���ӞrP�Tj�Z9_�-c$bט#ֺ�$S���N\���$|��6:Χ^n���H'_H�3M��.W�YG���`�h�#��_-��+Q�.����}���p�Dn'ت���%
V�_��i��ݨ�ES�f�G��+�� ](I"�ĸH��I�]�W���!��q���k��l��V����"��8!��	5r�7�.h�0��2q�1w7�q��9��V:6l��:�ʃ�K0���21��k:=�hS���mp� l��2�� 6Uh� _h��G��^��o����e0YR�HM��5fl�a�2DzCT���4�+�*C�+Ƥ&n!�az�V�j"�	i�s#x� �]�	^S�m���_��hB��`u߸!���P�7>���(X8?�8�8�z�M3塠(�>��侃G��8DjB�Ŀ��h���>�����V)?^�G��~����VK������-@�ѓ������x�Gk���)㑙��x7W�8fX�TfBSr�|d��Nk����$��$��řc.�������秫����7��܏�������@��d%�J���u����FekIG�h���� ��R�|/�{F!T�_m�I
���QY�d.��q��yJa�bЎ��\,�����
R~��\4I��`f4��wr�p�Z,`ϩ�b}q�JI��� �Y�g���ӀgK,p��Y�\$��dey�+ڕ��>���
.���� ��[��~?\o!&�'�m^�r�Q�R���T���*�kz���o�B<x�Cj�_��da��{�� ���Q颐1DF�S��}�����e˟_�[��J�TY�͔Ҏ���7n6��ˮ����	����5�|9�®��P/՞ZyJ���,��t�ʨ$�W�ڜg�(��ΡyzbA��-���mv�n�%W���
"U`��-Tl�����r���oN'r�ĺ��p�Y�(��D�ة����O�-z-VaI���7\����V��К��D�|��E:��*�#
g�n���Ws�R��Q�	������g�7��B89	p���P�S��ᆌ����jt؜���~�&����z̢	G��:�K�����h{��	�LB�|j�ڠ�Ȋ��K�<F|�_��y��2L��~󶯄��j?�9l,�m�Z�TƵR�a�@-.>lv���;
-[AW��`� ^��_�0
Si���	x� �u��l����։\�n��T%���>�E�]4��^�'h&m�w�>D���W�u/�nو������G�S3��f*�=�E�.�܀�^���W����N�$5Pԇ>Bm�]��ӕ0�½�/�߉��������ߐ���⬳������̆�J#�cK��o�� '�r�{jN �r�Qи�41�m�j5���G��p��z���=pC&P�&e)P�° ���w�*�����c��I��K����7���N��p��mm|SifI�r&��c@Y8��yjY־���_$�%r�Π�؇ZS��}T�{6+M}�6��,� �*J�Ԧ:�/�������+����ǂH��f+�aj�"���țlk���K�w�_!Zn"������ ��N�\�v��{�v�4�&�w׊WE�V�ؼ��}(t�<�ߝl�UOX6���r P��kT*�b8�$Uz�m�T���h��<޺#��'�;����P�m���C�J"q�����C`Hi�J�ͧ`Дc����x�6�m�T��)���a�=���$Egٓ_=8�uS���"���{�7�^�!���B.���#Vk9��e����$8%3��ѵRJ�*��D����o�(ǭ��n�\�%w(!i��rf�y�Ք�iL�F�iջ���^ۆ�o7@�^����5�\'�Q�����J�r����J�j#�,��������^�O'EC%5��*���.m�T�(J)uk>#�R֧紞i���v����$�H�j�����q�zA�1�������%�ʠ���uf`�	kV��L��c��߯&�X� @�?�	���,>��#t;�P�bX-EV'�[��S�'�g'�0Q��ZK��i���[ykB�tq���)5�6�(F�'����7�l%bQ�C�]��.���Eq0�9D��j(�bNCҟ�?������3�&����O��xo����*V����p�i�<����"~j��Ra�������Ӡ͈4'k3VR��Т*m�r��?�.�V�Op�-��Q������H��&8s"{��v�bt�/�{�xH`X�6%p%�t��eU��O{�{����_M���wT�r��^�Apa���cU;u�^���ᱜ�j���.��^�L��Я�q d��n�s$"�@���j��lؐ-���V�����Es۬Dh5-��δ�!3R���Q������E�Or����ܻ�� =���{�@�̟D�M�v��J&$�� N��!���\�Ȍ����������9d�޷�3�Z��$�Cǳer&k�o�u����� ��f�CGR��7,p��e���l���W��߫!W�!1(P�̱�	E�ә���XX?o��ń5���s�����y�AX����es0�N�v�)Z����[ǿ�����ڨbg?Ԇ��J�U��/�)W�� 2�M�W�=�Rm}( ~��G��O�C�;K+���v�H���7'�ߩlh��U��,���)ɩ��F���~ se��*]CSY�[�ቋz���I�MTq_�~+8�[WI�?��.
c��sx�x��;@�F/��3/)� Df����{%*�?E�e
����S܀���q��s"P�6����k�J��A����)���@�(4���B�a����S�T��@�tx�Z�S��OG��R��$h�kD۝c}�{��NUϧ��kf�#�^I�[�q��z~/,-t�:��L��G�Q�Kx�n�B0� =��tb�-3�M7)�B��G�2���M'��>�j�7�k�Cj�+Ƙ�D��~"���}�_-̈-R���l7�B�7+��X=�2mҊ��+3g縋r�ژ�[�����_d5��*�� G���
�S���e��f���~ȯ52j���q̄�\�.�Mm��U������a��E�[��df?�5Ow(�P�m���㼧�J ��ޚRj�Zhy���s��.��TGG��W+2̏Msz�Ɏ6�F��s�i�>#Su\J���!�w��oӰ�L� <ш99�kn�3��q�$�P��7:ޜA=5-�jπ��� �~Y�d��{�m��q���A*D58�xQ��J�)Q�C4�L3�y��1��Y�ܭD�Q=tTX ������/���D���?-����Ԝ�t+8U���a;OecH�x���H�Q�-vxBQ1���~E�s�����FX�={VW���jrd^6R�zA��pK!BHK�%�#T��}����1�0��&����|���i�=狊����v���8ȹ�L�s�Ƌ���x��C����Kw5"�Ѭ+��g]K�����K4[x��)-��B��q��rE�����L�\`��rM��^�����:�j�Ey(��Q��f���(~�/�\�B�İ�6ԕ��H��)�wk'�����ew���B�����lײ�W�B�z��b��pO?B�.G���t�\� `S�1�}}���P�Z&�)�˘����aU��B��{�>�l�O����נ���~��b�zE���d��w
��B#u�l\	�Vpi�0&�P�GG=�'�t�?i$%t���'y���7��vQ`�=P�� ���	3�@nU�	A:.2���u;tX���n���r:��a>H��[�ܽ$���\ ���S���Nwf�i0).��,��#6������u���!:q��qp�:2k���tL�N3{k�;�DM��C	}'U�ט%��] ���N��������)��c��ZM��e�I��et�e��=�{�Xz��H�5�<o��/8E2b���U消��%���	B���D�?8�X��X�.��W^��<U^�*��RRw�	���[,_�1�5��2��)D
E.>�}c�p]_Û�vgǡ�E������wabJ*Ց������Ư2
$��+��\'J��@��]�[�-n�N$�"�ga�VE��L����_�ؾ.�I����Om�;�pD�������T+����%.�.�heڅ΢P�c�8 DB��R��0�����`b� K�F�����'U~):�\��M~�;6�o/��=k�!<����u�D5"�Ձ{���x�=t:�ۗh����D�6us|@=��MKRM0��35܄�Y�a����R��!��a�Ȇd�k?*U�?9ﬨ!�Y�%�AK稿��[�6��^�hm#:H�aI�y��D�8��63�����_M��T)�`���5���x]%�ڮ���U�?޶��B�(��͑9����Q3��S�,��D�8	��):R��)�R��_c
ꑀQ穨�� �/	�M,%&�Ƙ�S%b�8Z^k�|�/��QN��
�eT��6�?+�E��4�C5%�߱eX��v�M4Q�6`���SC�N�y�aХ��~a�"|��Vx��.��f��^��N��~����ge��߄�)�����D~����}�N��5�1�aH&xK;/I<��SՓ0ʵ���-����N�����;�R)0
+��$�4�C��F�Rx�w,���_��Q���H`1�k$U*�)mf�s���5k�����(��d��f����4E!���/R淫�I5'g*����/��3��j͜�@�ikT�nmu)2@]��=������6v�������vD�{>�}��f2�n�T����6qAkK)��S5�@æٗ�
r+�P+���Is�ΐ&l��{5�@��z��챮�>�7lA {�kk�9�R����4Y�V�Cr�ڟ(��ꋡ
��[�r���kˑ�,����@�wĠ��ĴjT�-~�2�x����0����T՗t�'�n ���[o(�����b�.��dl��eG*�(o��g#�~|ځ���±�ĉ�vz|jy��w�5� C�P�_JKXL����U�9*ve������o��3�WfP��Z�Y�K���Hj1�x�u�o�/7/M��6��FdkR��|Lڠ��7�b?1����MO��*�#������O�#��%&�E��LB��w�lق����ʎ��`x녈�ɠ(2J�O��(d�3A��B{�B%�)2��t�ဪ��$U�)j�؞0��6c+{�m�7;��ے�`FcM~��P�
k�O_��O^��HP'Fs���?�!��\$-{3}!�-����ipaf�C_�e�<G�-2ٌ�$����K��D��:`�l,ѽ��ۡYd�S���:ҙ���nw����dY����,��-3�{GbLQú����!��[��ӟ.I>�[r�?pk��~X����Lio;��O�L)���}8\D�=N����rQz����V�<Д�v���f�F4���f�Qj��5����U�Y�K�}N�'W�k��k�
�Ùs�;�`Z��Q@o������;a�}&�J5�$]1SU�_��S1Z�^f�E�|��6���t��?���TNf��s���tE��!���~�;6)QI42:x*W�D�@&��a�? ���Z�n�h���l81��k2ѩ@R��a�����@O�����>R8��xI,K���tP=(ۤ$��)U6Y��y�`>!��!W�RU3'���~z��&0�������3����?�k���kx� mV���H!��kr*r8>�uո0��7a_��Q��3l�4'�j	����,�oM����aJ4'�������$u��2��_.���T��Lb]iT�5I��nl�*�G[$�R-��z���������� �14_�I��p%��s\����ď5��q����D<�,��o�/\iHz	o�,�����j/	���+F���BϾFT3�p�x��Х��v�~�{��I5�?��S֛{]?p�Z}���a'S�8@�����������<�2z�m9u	W�>��^�K�J���0wͰ���6�Ӳ��*����$ԋPkì�ӭ	ɥ�T��O�fi�Hn��P�����$5�daB�\�񯤿��@tG&O5y;�ی��#\�I=\C�N�DH��k^Tj�����%.j���/���=�o֜���59|�8���1Pe�l�u9;wdm�O�V��w�#l�����n�'rX�Ս@^����N��������#��$�hU����(�>�>E;�6=�}B�	*�����"�^� ���Z�:��O5����.�żӉ���&U�"��W����ޯ%G"&s~o�{kۗ��͗���삿����w�;��~}���^�!�3uG�x���GAf��[���QCe�U��0��(o��c6���-�B�Y9�ar��_�j��߀^;���k�C�~α�˝# 9���炽6�ɠg�ʃ^� B��['<ZmS�a4�Ҭ�{��Ht��q�>{���uye�u�VL
H�I1�M�we�3�I���+����ýݩ�fg$��s�ϯU��e*c`��_����	��Kt�YoTX2�a��P@���&]��^�t�[�/ϧ�aZ*6��o�w��K��m� rx!� ����y��`M�_�����]�[���.��{���#�5ԞXP-A�@>���]8��e��]��5�*��A>ܢPejT�w���L��%z�`:ݚ�J����/YN!Ñ��k����2cmgTQ��e[;?k�nz�K �E���T�l8Z-������BwP��';�Q>����Z�	���ʎv	x���02Fwz����������g! ���a������Y�v��i ��Ov�I(��5�3�RH�ˋ�ʠ:��u*O~89�/m�V�3�e1�B�r�L�qN@.�9AT	�`S���=O62~$�F���f�Y*uGs�C3$�Ap������f9�V�Q��Ы9 @"$c1��ֵ{���fԓ�h6������G/%�4���Z�B��7JS��J�Ѧ�\�����|�{�A�8��`s�$ �Fօ��>�mI��_���\Pr���.(� exΥ�������7�3!�r��H�${�*ɒ��ߌ��]����}l� W�gS��]SM�qV��}�S�{��f�$O�(*S��NC��:2��ޜ� ��۽C��df��89Z��g����3
(S�݊�֤g/=�j���>o����(-d����vZ�{�Ee^>ѹc��m11�e!�h�J.�o	G1��P�1�.��w�q&���{��1����J[��F�X�3d=�5��Y��U��a���{�zFDꨨ�.�I����軝7����w^l;�͡=��l[L�;*oc�,�q(��ϣ�j=��	�\U��x����D�J�]Ԯb��7��*ʹ��VD��P
�37f�SZnP�d�騼]��aOP�j�x�t��M&w$�f[٨E��,kC��|߳�؈��b!�Ez�^��x*#{J�OPb?T�xO�/���:�vჲF����&�aˇ��R� �oN���c ��$��ll�I���WZm
K4�G��m��EsJsQ�72����R����n3)epK:�(�����T�9~��Ā���2~Rɠ���^�BŖ�'��.�4/��MWz1�2� %(���x0�Q���K&����Fi*rt�h�%=q+���ϯ��<ʋ"��}p8+�{+꺄V<�}F&5���	�YyB%n��n�E#���)�D�Y�k3�����]^�Z�8���P�z��AE =Ҟ��yJ'�Ba=�A������݃iI��l6S`8�:���ĭ_��ɖ����G�w*�Hl����u�M$^���~�u�r�B-r��c���zA���� �k��c�~��;��s��NX��o�\-�� Hk�M�a31�,P���O�ii�"��=DC%gҩW��}*r�3%'���+m_�]O����/��ū9a9��ncl�oE ��Uea�����x�r�D�^�5p��@��_bՍ {��T����Uت�_��=g�ª�$L�#�B��M��� ��i1�7�Ь��)�m8�����1�ޟq>Η�ji$3NIq�sqdհrp�="�X��sq�	~�-M.�(:K7`,�x#QO*0��	Nlr�g�z�w۟z�15Q?,L]Ǭ�'�=�M	e�����������O���������N� �6u"�ת��#rl8�z�;�8�dP.Z�7��4�{�����,�N�΂��H� �	ȳ�T��LM�::�>�HͿ�%ME�����mo�"�MS���21+���],qQ��
����K���۪��{9s��-�K|Vo�$����R�GCv�U��x�>�ƄQ2�/R��|[c�U��l��� ��>�$�����|��h����@�9g:kx�4���RG��W�`j8����d�Ћ��g�d��\���{���/F�Z20�h�9&f�M����]����qlԞ7�&=��1;�@1���{�<ݗ�5}**�;�ȁ�n5 ��z��z}��Ba�A�X���b �[#�v;��}��]�q��/~�ۇv]'��i*��b����2��s�FM�Ъ,��-x_�o�D;0p�[C�h ��]���s6���~	� ��K���רF'fO��!�[g"o*�W��n���M���0�m	�̰/��"�����g��l�N����?Y�p3��&5ð�z��pB��Q�eN{��m+���'xorc����Tz����~�Mf9Z�������Fz���*:X��ۈd��݀�=z� �}��i��Y@)r�W1�v?W8�X��~]j�zf�K���A��}�x:>a�l�����1��
,��8ޯ~a�~�w~O&3���-���)�� �OS��'v����3ul��n�����^��)Z��1���H�WF��O�[_/���@lWU!}6'�;l}�[f�i���@7��6j� Xsrr���n
F#ʲF-n��FGq���D�m�31sp�H�d�~,36�����
�:�׭mz�N���X=����E�r�q���z��b�v���[����(n
������ؘ��K��Z"�.�c&�-�\�'٬���-��[����g�0؏'7d�����s��ܬYg����~�̈́�EO~+`�#�#ro�`�������c@;�sФ��X��Hzl���w~ΙI����T���Ws�ɑJ�*�/�w�"�I0�p���J�'%�=�c9sW���!�P�PC�!!�j�s���c�oi���v�#+�{��J�QH<�C�Qh�# �Z.�YYq������&)D���V��'��d���.�E��(��Xj���Pez���	�
�(����U+zd��g��%����x͋��S��Q��o��r�VJ�K�Q�H*T+�1��z*w��M�햌.�:O���+ȃG���̑��~]��uaX,u^�ێT��xƠ}Z�6���1�Wgv��q��1Z���{���-~�[��l�o�/�(��]-�و�@?���+�5�ߌ6G:sɃ˃S�8�p#�L⃼�(��şioK�b�e�[ �C�ivb��5~-�<M��_]�� A�B�ԥ@i�+��!��ȋ��I�U�-H�n�-r��ib�k�q���vP����������S�<�!�.�ŋo�D��i�OG�]�#pK�%��&V_��2�HK�r�a���r�v ~B�%���F�M�!��+��K��$���+G�PNwY)\��	ޡ�9���7���6�Fj0%%��uE9����[�Ax�����a�-�C�}E�sBC��D��	YߒZ����+�:�t�e8�\���q��.����`z$��c�ƨτ�Ǭּ@�[���ЍG��2V�w9'��Ȑ���9w���<�W��?%u"�C����p�!j`�}z9�����*L}��%���]<ѥM&6i�Ȝ�F�)`^�O��T� 2�;���r�;��a�43�������I^�@����`��G����˸	��u�5-x���w���!;�e�������M�R��o!�����M���C�)��\�2"��ꖱ9����n$�G/����sqaD�����|�=��f����Xw� �x�̀/>�sQ q��E�jh����Ma�	��b&�<�B�N��]Q�?̑m2��4�y��"�'�r	��e�#�wj�]��r��B(��;w����{��$���Wxum�3P%����{)�O����R)�cn��5�J)U h�<;� ɱG�l����`p��=���ֹx��7�eZ?�\N��Fkڬ3��c��
�g�-�!�zi��&%XZC,\�xh�B}��fo)6h)=_5C���Vva2��O�CH�( �eLJ1������}�?e�z�����SΡM�ď!]1m,�����;2�H��4dH����W��׶�R��j�d� J;�������)	���t�^tW~@X�I.��┇�v��/�7r�&.E3H��r����IPc�.�Y�<iM���_J�/�td�����V���s�t��ʶ�����.M��I�����!��殺�%�.�Z�Y² �K,'��1h��_&��ӽY�d妶����ISƫ�E7&�95��+y3&-	ܗ�P��b��ŨUY���\J��G᫝�~]̝=�ƋF��K�Y�B�-$�Hy�=t�*jY����� ��g3#?$=���蕴���{��,�HP��]��_�&��8����H8���ErA���:�CI-j�۱Y,Z��M�+�*��c���,Tzn��t�-˭�������i�8[�D��v�[�>L�.�B�!._0R���Aʊ��*7�b�R������:���,���3^Ia�,�����1�ɟ�IW5$}	b};��0�"rN��T�BZ"ע"�=�_�԰=�&���OCn��	��%ޟ}ί�C�F%z����<'��^���c��-��SGǐ�xg�H>)RL��$���|�|[����7���y��X������9�HX�"�%���.KWŌ �Pz�/���MѬN�8p@L%=��q� ^&�N��o6]^�2�@Y/̬@��}!XM%*7g�?��ǯ��.�<{��F��i��i|X�O:�^>�n�Οׂ�FOaf�76�#5��㰮J?%+!�,S��?� x�&�@�L�K��FN���{9��=vtê�h�IńUi�R��'�&p��զ�qYZxڦ�5�?�ٗ�!%6u�э���/ב@�(�W_�M5����i@p���1� �o��G:Oa?$��s:r����u�����urS /N��]�hJS<~�z�(��Z��Yt�dX��=�`����h�O�K|m��3�}ͥ�&�:�TZ�]�ZV��~F`u�^{t�e���isa��H���H=���U�.��F �f�����Z��O��eMlE�M1M�u|�4�`�"��D������h4���8�|�!��Hi^����/�����#��z�=��R��3<Gf���4E-���ց�"�rX���!��)�F��8�,�9��'*�g�1q�>�<�i�Id�CM"e�?$���{s=mL�\e��э0�e��G���.�̻XA4��I]�C��92�B*\�+M<큊q����\z�7���?�6F �E���@�A���2��%�ަ#P�*������� �ݚ�*�jp������k�[�6=�9�#!t�|������.�@��O�*>y���p��'��&�	�2�|+����	l1u��]����Kp��ma~Qv�d?��Q�&�n�RJ��<�9�<e.FLzO��식ď'���X��,UK����-,�/��B�Vj��M���p�t���yh���;��B����V�R��Baw3K^ڔӠ}x�t����5��K/vU�4�O�ޮ�̳Qf~��1���<S]�D_y�}�)�:�����S_&hG���2��t����`�e���1C$/������ݼO83r�,qs���W�tP��A$����$���s���<���y�l���0	/�Cc5�%�����)M�G�VG�"u0;��U���]��O��w���.%���	Կ"��#�Ȃ��)��zOٍ�&����FF�O�p1�S��xJ�Y�H%����v,�p}�a�.wW���qg6j�{$.`���g��D&�-!�LW��ګ��1�����Ỳ`�53�����Y�_�!�[iy.����y��_��fza�Z�����]�\_A!����DY��t�~��aǝe~r��\����7<�Yi1��tGz�w$(a���)�fMF��
kr?���=��"�ʅ�t�Ĝ������'�̜?�֓W'���=��lz]ib����"��~���>�����&��YRI������n�:[j�������6�h�`w�E�py l��hІ �ɐhs(�h�0�r���W��Rnx�ۥ��\TyD�1CB����blq3�
m�T�+,�y.��pz�� ��-Ku.T+�s?b䝸���rf�"GnN_)�@�h.�����&�SQ���MMc��(H߽Q2!�+H˨�$��<�@r
;Z\o�A�ʀ_�r���.;C�&_f�x{�m���a,M|;��IcWH�$�]�c��MW��hB������O6���T�5�r�ZZeyfN�@ R�Z�k�i)z��5���Oq�M�9�&�(qEXvƺ�RƵ7x�f�(�y���o�L`k��c�D�:�5d��iV�vx�xF0{�y�߽4x�r��
�_@�9@ ��-R��S� ���P�'�+i�c�����&w�a�X����w+���Y�.�ؤ�ZE�
B�*����y�q����ژ��p�c�k��	�x�t���eg$��� �#l���^LΣ�;�9�{(�l�?�����M^���MP(Y�58<�`��'cvZ�VS�`7��HE�}�1m�q�r�U=�������}`�1M���������Ru�
�(�\�O[�V��fy+#S�^bmi1#u�v�2�ڥ��s��_L��[<;�?R�N���gE�b��|���i�N.�S7>Yv�m���Q�\��SY)ڂ���b��B~D�ҏ��4Zе�χ?w@<3�LAM��'K�qufi�� S'Y�ڛ��&�O�J�á3����rl��9� 
7	eXGC��vF-6$����|8*2�ϗ�I�T���gf��˥y������3R.���hv����S�5D�_�h1�\N����Ĥ�֯�h�G�U�.qY����B�P��B�w�\an*gqh�5�*r�Z��oz	��7,F�AN�S/��A��(�"���\�-����@T�~�o��G�/��LPe�
8	�W	I��z��$E�;D(.��ŏl�+l~}�ys��>�j{�K.)��2���ԓ�%!(7�
A��W0YL8X$Q4Mը9�[R�ÛRt6&�U��˟0��T�i��mZ�4�È�%�gD|��_o&*y�34��d&�=��V�^�:"����%v� >��ʬ�j�Iykh�Ԩ%��`��me�b��p�Fi��)p�Sn�)����4��=�>?�nc�A{Nq�(���t�#�w1��; D���G���	
_.E�7�c����	*#��5��#���0���b�>q�lw���MgىS�V���<�[�#HDD��U�����}�!|v�lH�;*V�h�d�W�*��o�4�]P����Tկc68ol�$����xI�զm:�"X�H�l�\o3������IXǂ� ���*՟y2�??�V����f��z���@Y,-�!cQ��~%%P��=#���]���N�:�U��j Z6���IJ�6�uȪ��9q��1��=�/-�m�Զ��t�=� 5Z!G��@�fŁ)�|�E6�-�����Kp�	� �� Э���ۂ��'Ք.�Ŝ�2R|��-
n�#+��㦺��\��\�W;"w���*t�U��Z������N�h�o7U��[�f��~�G1���m��B���[y�{�Zֿ�v����d�y=1�Q�' �G��@&'˥u��Yir�Sr勼 |+�B0'�w������5Θ�GO���KYi���n����N�rA<��Y��?����!X��v`"�`<j]�N����wI,�b��t4�A��4�20'��q����"1�{6�U��Rp<"_�V��-,�V#���(�&S��i���8�|��
A.:ش��lZ)9�Z��P���8Hh���V}�,�"�D�!��u�����g��+@R���h�o'&���8�6���%�K�@���o�F�Г+����Sn.貒�,�`�@����Ʃ�I��Eiul`�ݰf�����1I�:\WW1��i���_KL	��oo�et��j�Ӛa)��	VG<�@.�G�����Ú���I���,���xV#��-)���A����W��Z�
�w2$98;�NƗ:��5~��� (D�B��f_Q�W ��ym���~��-h[A�c�s��ZkX�'�F	ȴt�:`i�)4��G�� ���#-ko"��gC@̶cw�������L�tF�B/v��<�?�Z=�#��0��0$�7U2�=B���跚q�N���	S�Ln	.L�rp���%T3�b @��k{Ff:Ǆ\��*���*~gLي�ˁ`�'�@�D��x�\ZB��'�B��t�B7`u�����y�	��(����{��h�we��B=H�b_�=9ߣF@��,�:;QQ�RW��-_�T%��`>��S���x�����d��n}A���-�[4S�)(�s,8K0���ӡ�P̧�Z"�E�JDS��e��]�����7�u�X��K$���3̲l� ��qX���fx�^�Z۩�ǡ�lϙ�LW���k�,r;��U��<�M�B�(�Ǳ��A�s髳�Zޱ��l���I�wM�x�V;c�ז�&_9��>���L���7�_��y����Y�����/����Ԇ�����x!s�ӅVJ�8����H�[_Ne����.%������z%>3!���޽��jH�XƢ7!9�e�J��&�y#p�Jϒ�ԖO$p��)i4��!] ~�0c� ��a�\Wpv}��ޣ+L�`�S�R-+����5,4X4=�=9K���*���'��>�W�������"�2���a"�\��*�_�{#��#�^��?Ne 8����Y���IK���w������P�)�̒3\��CN����~��^�~0�M#�xܨ٪�8��m��M�`��s,(�d��q^r"��,[$�c/e\y���y����-�#x�{wXS��N F��kG�
�rJ���� ������	3�*�M�h�|$�H�$`�X�6h?��B�4q���z�Ew�,>	�*���=&�:��"ŝ]�4KH�2؆��aPF ���?7�?i謏GuF9�X�W�Z���	���"��2QeB��D((�%ʮv������IJ
ɒ�>9:�w�睸��o�\�� c��K��(ݓx�V$a%�2����=�����z��A�ٵ��; �%j��|�-�ǭ��D�6���Sޥ]'k�q쫎��Uߪ��'���'�nT�ʐ��J�0�8Ҁ<�@FE�*;�F�i�����@����)�;G^%���-����X��N'$q�f�N�Jp���<���\�BT�=���/��g�XzQd�䬊�\�/vQ�j���8u͆b���@l�y� �w�5��n`?�&5�����副�g$;3Y]�1Mo_| I=�����$d�����A���}BG���\s,��|b�L>c�r������5Y8� fx��tW}Q���]��CODn:�-)��ד,T}N�qkUo?���`ҵ��>B�<�I��~�}��`���Գ����U��������$z��>5*���Sr�(8�"�B�v�/��Ӄ�% :'�
]z�������%!
v� xq1��9?C�Q�;�&2_&�_7� ����k h*���Vg
�標�'1���-w�R��a|�f\��~���&����uPh/z�걳��ܳe�T��a]RV6�����D��{&4Dhan�(����������h�t�1��(����XZ.�H�;�k$��{uc9�X肵��~�ϒ��K� #�u��%lI�L�*0��V�p�x�(�:�D��>�X���%���ly���RA�/�?�WM�.<�a.�w_Jj��b�N��=��P�,������u��&�YI@ʓ�v��$W���X���HCʎ3�0�|�4�Qݟ���J G��`�L9��O�F˂&���0Xd��3�ܬ,9 �T�֪��B;�t�g�3a e%�"�
 &��Cql��������5keR
΄����f�]��h�*i=��E\`�����ς�):�N��0ƒ%�_+o!i�\F@	����?\�_1��ȪG�n��%j���L1i�WSۜ�:>-�c���h�ϓBT��@�,�z�4�����?�/Y%0�'���RE�ׅ�����j�����Ă���8U �P��ps�c�I4����%_���>��Y�l8���j8u�u�N�����_�U�϶a�l���z�Ýgb��ԍ���a�-C�(G`�j�'h���C�qc��f�s;�8/@��Q�Vթ7�CoU"��A&�<��"\f�^��9���z\��j�et%����d�?&���3c�z�47�@V))�N�ط����vg	�[���E�)��_�ۈ���:X���醙����H�l����y�+���r5�.i�����}�^���Q�w�w��#�|!	�6�'4����cGe��ǰ ���nshߪ�	+ .Ճ����;t5r~��W?FS��)M%�"���� l���s��0��(��@�<p�>���D�&���
��<˰�Jm��)|���.��Fs�߼������כ�J�1N���fO��_Y"�_�v	�eu�t�Q�~�S�`��� �Qj�5�����_��.A�t*6�C@$��?��I����2��Q�spd�H�sǉ6�'nr�RN>�B�3��nz�~��~����9,�]Z&4�k�ܓ��kr�;��D7q�&&�"`w�6��z���j��Uxd������r:մL0������^�'fqV\�}#r�Z�^R����|I�;��X� 
� v����φlX�8�~����4���Zda�`%�bK��4���~�+��.�;��|ʐj) *]�!��N���Pu-�~�4���8��T��U�N�EN�;�4��J�k�b8J���;W�3 �^�d�;�z��;H%m��-����ϐ��J*u��ߏ��?����~�䁽&��X�+��IV�{�)W������C�"��\g�YR��6|��c�O�/?W^05���0��R��!cضM��V_��'�)dA݌�ov��2V61���?e�������K��̱��֟�	�����p��_M�p����q$�ݖ��m�{�'\#��F����t�.���^�f�K�ӑ�d4� #ZW7���i��h:���z�O�D�¦'�z"@��t�?����c��$���;1{6�DJ����E�燾��x���~����P��ӆA3�3?{���!��1V��{8<v
�p${<���ǫ��kcǵ8e�D��&eF}�W4�!��h�Nо{�V�3[�hz���	{�(��ord�k@$�S�����=����� ����z����xt롯j�J��XZ�7�]nDF*9x�V`ouSH>�Nmֹk0-Է���1ȟk�ڻt��&�����Z�>��e�%�me}�OS^����J̧�����F3r ���c|!4\E�O�d/I�� <0����{���I�Y��1�.yJ���I�*%JHF�,���P#�bu�;7�ᬎVI<�&y��d�K�~��ܵ�V]yv�@!��i��o�n8�tJ��}7R��,P#Q��HE��uB	n$��=cw$������4G)sz�[�v����3�� SH��j��
w�sL��jל��|Њ�a�)���T%_�P7���$�7�]}᝙.X6�뺭���!'�X�s�>�+#ɰ��Ȝ�%;��Sӏ��HcV/���tF�n�)�NV�_b���I1D	Է�Q#����(�X��۷(_H��yv1;���+�IA�%7JD �8��G��^I�	S2�:ق���zx�-�l�`��K�p�L�/($�K8�z02�r�϶���[�}h�E���Pӣٲ���[�.Y�$�ܠoSsQY_z��(��$ȎMX��YevdBI�/f2Uh��l7(����GP+4E�09;E��;�7A��tj�ek�[v>��!m%`]�[�ly&�
��R����/eE���Tn��ID$��[e�-�
{��b.N��6`Щ����]d�������|E5��|��
uS=X�M��E�F.{�n"!3��!��lFw� pU���ꤽZ��W��}�!��Z���J)I��ݰ�$���pC��er�d���������i�L�$�Wօm-����?�˷z�E����'�}��WO�HF ���uB��Z�Z�H��n%�\(TZ�Q�J����4KS�q�b'�A�2<T����Kf]��;ǋCg����OJ6�Ҙ�#����QH����緒����D�1N��=�e��t̉�i���Ġ�S�����۪������ṸU���;l������ٸY��C]��oM�(���}
���pq#:Yl8�׵Ǜ��j��w=񡫄1�$��q�OZ��C!
��<E���Ì��Fc��ղ�.f5- O��W;%��q>AS�>^4�e�)�YP���c��e��H�֝u����{}��[���H ��lv�im�E��9�X�yd,�s:WW��������~6g��^tq�ډڎ�`�1b���1"�F��1��eˉ����iF��r�|�&�v��ޒ9L��g�@_�/�=���.l�����o�E��j������Ѱ���9��9���~�u^d>�U��l��C���R��M��ƣ�y��|�K��\<_#�>��z]	Za��P��Z��E�/?��L�s�y�C�H�_HkV��	&H�_^w{,����Yݧۤ�\5K^��ޱ�S��rR��b��ԙ�GN���S�(���3U���~�b���O�[t{E��^����o�b��l)�hW�� ���*�8�4,��s��,+Z�-@k2��
y���»E2G���"�L�1�f�|2x��&����~a{{Y�뢙�o�1�	ȹ��٪`T��>-h�@/��"&�g�I&|���"�?S	�:G�9y�l��4�˛x�����t�Q	�W7���~H [з쮿B5��:8�9�P���}�'I��m�B�&�.+j����	�\�O�2�V <�5`�Jt@-������tޮ�r���1� HN�>A��A��3+�^k��:B�|���~X�g�c'm����	?�����	�=��Uj��ݛ����4��$T�aͶ���=�� ��Vy���)�z�W��]����ʁ�Cn�V���e+e{��l�d�{f�m� M^�'��d�t���{)�5�b�oƚ@�U�QKN'�s��|QP��qTcga���v"'m�$ ���'���8��m�i�.����و�q>{|,+��Q�rìu��i������3f��������+.���?� p���W��x!��0�\�@��ҷ�Z��/V��I� O�a�cYѕ�^��M�~�y�:/��_
~��3<�}Ͼ�w��*I�[ň����HPI�����݂.c��ds�$�a�� ��Iw�giC踈��I?�N-q�����n��U���'
F�D�i�1)*�π��Q�ѳ��Ρ��p�6�'�m�{����cJ�^2#�Fl�7N);��x��z��H= ���2Y��d]X�y-"��{�k��L��[�F��~�I�Zu"�����G��s�_��.���BK�­3`+�T�^�-z9
�Q炅1=��2!��C�� �0���/��XR2_� ��\#J/ _���f'}l.�W�S)����2)� 65j\�>���&��6il<`?�,&z��v�1��!��w���[2V i�T;rO᝼BB=r7�Q>@�Ӌy�"MW��i���V&�C��E5��;��%w�d�O�/�Y�����MV�Tv��`3,'\��c�I��=����ZVp$�0��ї�ʥ\"H���`�*�$(s�3�.�O�MΗ?4�R@k"�S���ڟ&C)�=�w��N����1���`>��d�B?�����Pco*5r���;���L)GԦ�	��3@D̃��ߊ��`j�%?���2�����A�<�T-d=}	���#TK<)��cC��{H?}��e�d��*�}��BFq����V��ӟڢ�Wоe6� �V|�R�=�0�������`�{���W�k[8Q��]��9�^[����r����'�F�Ltd �G�M���ZD�Ϳ ��4`�> ��M���#��?�}4��Rg'T ��=%?���@(����D
�nI���:M ���;�	�o�	�V�.'�磼���3q0v:#��vf��!��j}��?��&�����k&s���:
�2���*.��X_�ӏc�;g�kw~nF���ee�������N���cBx���-��_'��QS�X�٫�)2�m�N�8����ݳ�d:��|��2^#`C>�"c�Cӛժ�1-ŲJ/� qd�X��w'�K�ɽĢ�qSE����Ð!N�@�3����l9�p����"1:������ݪ���c :��Y�y���AɰMь��ٽ;�x�f�2�B�8�@/��* ��k�5/[Z _%�� �S��[:�.�(�!I��_�T���x���[��
��pY(#<+H����ls/���H%s�$�T�绽�U����r8��;@8;Z�^'Q�I��4��b�lr'�G y���H�p�q��б��\?؟8b8���ػ�����t��;�
�= }�H����5R%`���W*������2/���-�N�������]�O/�'�-�צxr�q�!��	�hs��{���b>�.(���GZu5����l�婀'��f�J�r�Ij�	(,�t�J��9�7&4�0M�}�SdBq.��SIy^ޘ#�����1������٘<�М'fr�~]S��R�n�-�$��,{����ʡ%2 6;�|*����'9���`!^0��tB��f�@�� �h�Z"?���'?��βW1�#��h�~e�ш�p쾆#�|�SH�|�	�2bڵ�w=�@�vM!<gݥ!�w�\ڕ:;8_��S��zܛ���dA?;�+Ch]ͷ_^~�C/��L٫���rp�n�<��� ��, ��_��[��:6�3#��ʜ�8����qqd�e?}�x� K�՝���}�u��Y8�-��ɢ�,�������(\B���ŵ��#��ٽ�D�M9A5]̸�V[5}B��F��+.1��tqG��l��w+6�ˊޢ8Og��^un��_K��<�P�l�A<nQn�F��[����d3��|�X3bf\-ZZ	�p���2��w�3�ߒ.��l��!Uv���e�'�'�6d�7�������*�6 �����0ᷛ���3�h3�ߣM.�K��b�����
Xr�;Z��~�OkB"��U�e>o&�f̫��t���5�^�O�^J�࿈:C4��8��i�6�A�R�5�dW�bF>9��%��hZ�24�;�s�Eo@��
�-zW���YI�pڟz!�1ݱ+0�y8;�ކ{�$��a�q��9�u8<��ԣ9��G�}�n�6���x�L�@~ऺV��^B=1^"ˏ�<���	��-��An��kf�����E��!1��=��:V�`Ur�@&~G��_�`����z�-h�CWj�^��lW�>3���`����#���z�ScW��{`0=�A��J��Ip�y~�2�i�gr�e^���V��VlWΰ����5
ܣ����2���E-ڙ�[�gΗ�ۍn�g�l�Zn�04�S��H�uw��V���ˋ)� ��Y@����I� �_1+�ӾB�v��N�)f�����n��@��#q��͹4�<��L���a��`�`��&2׾Q�"�R|,�@��[�B�0ҡC�+r$��;�O7�,2li�>�]̙���?�LW}��(/x�R��y�5N�h������Z5(>D�h��43�AH��Ɣ������[�0��;���=���_����>=�j��{t���� ��J�۠�׍�{l�}��� :� �y-2wX�aW������h�2��I�O��5�h��/�$)��(�
��qkzH�F+.�S�qY_��2��>�JloF��EMx��.CH�h�ϝn�:i��O��Y�)^h��W9������n�9>�_���ׁ�!"��N����{g=Y���l�϶��}u$1�jj��-�>�3���������:OK���+��F���L�㠈��m�a�_o�/�ٛ���^�dN�6M|�8�1�O�;lFyQ/��hg`l��� ��I��)���={;���#��q��@����C
��@�bx��qE�p�"��Xly\�̓T��I{�8��֋�,"9́%���;pq~�a����N`{�sk�*��\,p7y��1b�l����Xy��n�ݕ&����u�.���e{�?.}|�蛆�3U�,
�H�����+��ʩ�S�����M����S��lS�\�3FY���ܜ�d�a2 ��:���&
��9x��㺹�����,�)U\�(0®9;!��D�������Y@"���1-���
:��Z2l|�}c�x���a	T�#Ǭ:��0Z����h���Im��{H\Mߢm��H�82~x�����_Ё	~�����w��n��fu�֟J&p���<��,� 3�`�3�ד�<���*��{�l��h'�+J����T*y�	��y�L2�DwS>��C6��Cۓ.R����&�b��1��D���7�Ё�H��62N�׾�L1�Yp @��;S�pʼ����G���~��?��y	2k��6�X!�Rﴶ�qnc �ڊ��|rUY�6Lpb7�t�W\gg��w�cq�Sr\�w����J�π�ƛ�3谎��=�&�b��0�	j8���6j���ւ9RW����cބ?D��(�Ҍ%l��&6��Rp�ѤE��z;+�Ϛ{���j�G���?�`{���y�엇<f@�R�-���'�9ؾ���@��vV��F0 WѮ9q,�����F�v���ۦ')S��2a]�cN(Bk7���*��{�g lIe~I��p�q��!������q�"!H�_[���!R*�U��H�**�~����X�¦�o<i[/�
1�W��2�ق��Q�����o^�p�V��/��ޓ����6jEǌ�/�vq:�hZ�"��SguX�{o֨;�=��<��k�q烸�^\_ę�:%CSw�;��L���ڰ�����aΰ6�U[�)�J�4Ԕ:7-\1�ݡ�A��1�ї<����vҰ�W��.--�,e�d λ�ݱ�����!�,��-A������;�����,.]>b�菙��߂�����+:�l]y���m�b�l�A�����V�����?�ף�D�é`fg�~(Ce*xI�`>��5�R��rJ-��aA��+���v8����?��St�``\���mĨbu�(���Fq��/VFP�O��/�iv�⬎���Q=o��IR�2�ס[��@Q���1%�t������n�$�r�%�w	�9F�d[:�{p��jƘ�7�*2��̴���	ZFs�i���뎦�B.ڜW�nņ#1ϝG�&o۪���U�F�Ys&w5����s��\u�.��j�W������o�|��aJQ�l:#��g���}66���z`Ť*r5�u>��;���"i4Q�v��,|e���%*u>��u�=�*,��_�V� ^.E�4:W�x����(�H�/D��/*��7 V��]�+f���J���hc^�Ё�D�=>;�>��~.���pAA�̿��b��o���xa^�"�%7]����&.�z��R���$����:e�.u�eJ�%�Y�X`�*�%Iz*R������6,��gW 
���[��'���!N۹���Jo�ףC�����X4�_���8�ٜE��l�S�Y�.�!.P�Q:hAW������hA���k�Z�_ ~b��/�D�ؚ8`���W��s~��d-�<Ԝ 9�s��;,�����~o˰sk��ݷ&=��_��:�\�h����n:�ў�zuI�Dp�%s���j�9b �������T����TTe��n��*y�&�d���h��8[�f�>��I��c}�#������M�5Wxv?�F<��a�l�>Y�_���uf�����L%e�`��4=��crg`����Ps����^�����J�ճ�`���uS#7��DK�8оu/��0rH�R�8���l��E���f+ۄ���{�3����IbA0�Z�P,� �<J�0)Y%�$D�/F�,YR�?������p���k*{c\�k/6|��~8��Ӡ8��W�f�&�~y�2�^�xknژ��%?�C����>�9s�`,yU�F���̜j!b���]�� d����s'�1r��H��|�֠��y�,ɭ����\�4�4glM���1�_���6�E��aK��E!��V�����3�]?�xx��e]��n揀?�q�;]x>J�s����Xw�`�cH2��,,�Q�_t�=�����L�ׁ�ƭ��b8<{"_��`7�%9ot��H���������J����*.ɽ�,@d��WJ�w59FB�"׌�NL��dH9��#(('o&��$x<t�E������<�P�Fz��1ږ�S9VNݏ�)2+Ꞇ���+�g��ox�Z`����ʋ�>cۅ�?�s	���V�+���� s�U�7�Th�(�0���ǁ��_
֖��4;���.�)� �AvG���lD�&�`B��v5uA�c�ם�10�N ���;� UI�T�nN�P2��m�oX
7��"R��z{�B'���^�lʿg"]�"��xh���JW|բu���\��?��W���u`����lgĽ�<���l�M� 8���(�%!un�S��o�����Z`E�*S=�S�b���6�d\1W'�p=I�׋�zэ1z���[� �H3�L|!�O��p%1%�n�zQ;i�-�J�c�!wC�v|�h}D�"=a�"Y���R)&WB���H��&?�m�c ���FD�-թ��ܧ��J��59�_u�~+Vb�6�GDF�o_��
�n����ͧl�=�m^�����m;�����r饕m�j�{��a�4E�*I`�i�Yv�O�!C����e�Mr������l��M�r��8��՛��gP�������/< ��|��SUՐs�L=�
�4���z��P��a��}>}�Ɠ�k��w���?�<�$g��o�}�]V��yG�gRxWS�x7������ľ!/�@�/MQ<v6T���bY�.��<0_ol�ܝ����nBq��/�@�M´��C�V�4��k�zL_��O��m��DZR�Gu��{A�!% w�27�c���F�x��c+�v~V   h|UXm(�*_��V�n���>�[��x��5�>�d�ʦأ�{����G�f�K�?OpMF�����砱x�x:�Tp��0�m��3��g�.�q a�X�i^�E�Ӑ�t���\��]�,�[X]B���=$��0�[9%�����H���.�w:���$��*�)��g!�/��ߥ8�Ily���uOa��v�]rZg�&��)�EÚ8P�>䫧Y�+rush\5t���w����pS�?�`��ϸ ��c�CxZm�I���l��uN࿂�PD&���(,�g�K@=�,�7YtK�b���SMPMO���|��U�8<���L:�v�����lq��{ �9dV�����9�S�kY0@Y3���99���l:J�f��f%��b&㮌KY��#z�gP�]QF��n]]��}H��x/�v���֣g�k}��[���+Վ�Xm����5)�*�M�g,��� ��m�<�����#�x�O��G����gTb�q\�`��N5U�_\���
脥cB����ڵ��z���<g���9r3��yn�ٖ;�`���4��<����|�/�V�y̻AY��=�}g�����TJ�kS������w�����k�֐�M����>jT�������2��) ���+ 2����V w�������!�1Sֳ[伍�d��Mm��V=�oH�fi�9��N�q��5r	��K.x��Ȑz�+��O!Е�a:�+� �Y�m��y+��5U��:���^�Ojk�KK���T_����oP�WI�H� �b^Z�nz[�[�._ȅ/O��RC�7�$�K?h��|l[��}�@��[*��t��Q!*F�!�0~�K6�_'��j@��D��I.͛�J9�H,H���ꂞ���=Mf�½C�cN�-&�FY�RLS�Y�- �`-:,��6Yd�����g��~>��I�$��X���G�0|�p�`�4�-�����Rw�f�0�� ��*�������KŚu�qu�%�I��
�D=7u��=h�/�3K�NRT������(��|_l]>�-�s��3|��v:��~p
DFE�5X�Wλ������o����pc���@Ç�V��:������j�Т�ӉOyG��$�ȼ.�[�, �~~!��y�D��6օ@`Aa�s���c�������u=���Ԫ�����t�Sl$L��j� ���.a�n���^�����j�EY��_pދq�.�=��s�%��,6��`��*�c��$��_?�hw1��'��Ҹ͝'�{�ĿY����ć�F2���ΐ��0ʎ�O��p�|�ucI�����Rěy�]�	���&�:�Č�-�WY��^.���_!])�W�Ȑ1��s���6c�:�sJS@�3��0+VUD�bs��/V{W�?hz�
�;kJ����FQf���:�V�£�6�`P�̉saƮ�4t�*��qc$���Q�o]��@>T�c�:o��mK�g��O��(�Oqƃ����x
c���k�č(����Ͷ��6�K�a���:��[��K�Ri�PC�ڸF*�J����]?5��!?�&γ�-'b�QbI�왓�I}����8��>8uc9�%��~9EZ\9�8���t�iбq(��G���@��{x�{I�$!2.v:�%��I��b�8KX2�T���";R�d��p�P+����OX��T'Nf�����uPȇ���,��$y�TX�qt��aP�,"�H�d��Ӟ���	c�xz�3Ei�8�s�76B�:�$@Ju��x���S�n��Kv����`.����M�MU����Hɬ���c�����#�ӼG�ńYR��)����/�E�e�4�ϑxvb��Vg�}ݻ�Za������X�݁cWV	W�Y���>e�_�~�4j����b`�|!���cC)���Ө�h��.�߉f7�1���M<=v\��-#l,��ɗJz�t?���a�;��{�⣆�X�.�B�<:O���	�S9髵}�9�� ��hΟ? ��@9g�j�����ض���&!B�#=Ccd��1���U?�9���6:b��3V�M�ۈT
2��x���;/�$kR����_��A���⣖�qOr8����4���a)߷����&�ˇ<�7�*K���1���{��ƧZNصx}���C�Z)SA2ę��D0��T��x>�j5.�{FzŊ���s���1�f�Y��+�ZbO�q���i���8�h0ʚj��y�ۏ�=�U*�����<;��v	��^:
�ɰ@��yv�D�Ӛ�xN��zabR�R���g�>s�DfՏ�A�ΊE�}ʻ���	L'�%a���e�����C�j���p�5��Kάcc)�Z��N���
��0�<��������[O���Hs����r�#m��J�3��	w�	_z�����W؍�!үc����N	�n�ƪD���+,�9����
hpo�U
�q+g������Fh~�ǎf�����8aN ﵊V��y�l�^]ŶJh����<�؀,\![7���
�o����Y]�uU�ӄ���md�#�
Z���b��@x�3�N��n80�Y��	�
ً�e\�)�����%�T�M�"8���WZ�X��aa��&��6C� �O3 rU�l�7�xn sC�v�<�¿�t����\+�7{��o�g�|��W�����c�ɳ�0��$R�O9L��jW1�υ��
G��P促�+~pr�H$�A��# $�9���I��V�n�����0�r�����-� �\��"V���J^�]��>i�M3D,`e�ƥ1�Y�,�r��o7
L�/�3%L��f�����>��%Æ+v֪	kC�Fa�Q���>HȨ���k�*㌘�T����`����|�n	�BY�eI�[�:,�
�!����@�8�n'6Щs8B��9C�ȑ�Ǚ�'�yYF�>���R��<���I������%Pi���k]�t5�'씺%����Ŏ]=M�/��HDAE
C}B���2�;?T��|]����5yj�;A����c~%8�C%������AV�vx�D���c�3���21L���_@�+!�;j�ix�r<���[��8� u��F����2R�[&�o�ʩ;x�L��mU���V��mn+�AS��{�{�i�W�%����~hK��Ȱ �\-EFiR���\��ܮp�Qj�R����| O^���>G��#��exYBã!z��ĳR0mMBM���G@��F)�h��_���c�S�������H���~�r��0G�����Q�+`��h%k�2�#kSP�vxeeT��ٻ�_Rm�$�!��R����JʳGM��-���}���-_��&
%^����;�x�4_�tZ�A��'�|pP�a�����į�9�D�L˸���?"q�ɷ�+LM�<��k��S�	���k�?"9&���B��g�Gb�Bn�r�L��`lI\z��q���8�+��P�9�aѩ��/��ń�Dej��=��LM��t\	;�������ù��On�!����o��Y2D����T��Y�܅`�������r.�t`NU|?s��V ��y��5�$��UD�f폋$-�o����}=����R��§����,=�3a������N�|�qv���������Rp�=��m���F���rl���߂*��c Sxe,rG(,֤�0z�븿��Rԣ��΀TJ�YlU�V���M������V4��Lp1ߘGI�����ٚ�s��ql�n@��O�噐f�ƣ��D7_2���E�m0�̲R���d���r�e����V�s�w���ŕ��X�������I�� d��Ư*�m��u����zap�v��u�FX�����'V�H���k�������]QuA�Gl��d��a0�l��~0L�$�"Q�jc&�T��g֨��s���{�(��D��~���Z�ƴ��/��?׹�WfN2=���?�k�)ki���W?)T�Z��c��1;��qAƕ�{F|��N�:��TK�
�U���4�y9 M�E�A3��2�`�5��&|�IԻ������z��3��)1�h��t掫�g2l��|��ߗ���T� ��&�S��I�I�'
IOt;��(��T� ��]%Dl����s�#ߖ#�
O��5XA���A��"���Dy��{'�j��c	�.h��W$�d�U���B�!8���l�|#ߪt,�wU~"m�*ʒ��DŤ��S���|L�à���M� f����+�NB>�޻p�5H_��X�����n|�H@Ĝ�#_iE��yn�v���/f�dk�\`� ���u��U}�ٚ��Hp ������'��T��������=TK�p�A-����%��Z/#�iW?`ʵ����u{W�G1_�Ȏ�oC�M��HS2�0��i�Ʈ�Q��.�_�2��S3��L�0��ԏ\���c����b��$���N������FrC>���N����ۻT^�E;"\���7Kr��aü&�Ҡ��SAJ����,׼&)��ԟ�s�����ڍ��ĳV�$�G�%��3v�\��s7� �u�T��������^����0�|[P4����q���"]�Jኩ���n��M��NV�tp�9��,�m1
�e�{�i�F�l�c{q�sW���1/a^y���3$P�����ѓ��b>��Պ�@�������1�׫�|�Ƙ9����0d�oWc�0�qU0ZʑY�i&!l�%�|�X2%o��E��t�\�_���{DaE�L:�ϰ��&�־4ӒqJ��D�@��wN�ɧ
V!��7��^�\o����lGԧr�/���/�b��8ȶ���؅������~� ��j�����I�����r~0~<�s�Y�����:�=�ޭg= �L��	qwҮ%@�����Ck�� J��8�Ӏ2��g7�{dAR�S���(�g���UL�Q$��2 '���oa~ptg����Z랇M�v���r���o���1j�>�C. ��8ޓd�@�vE���?Ĉb2Y��3:����ln�����CU�5��nsrtn������*��_�TE���cW�5���r����M����0ns5KF���إ���qݽ)<�Į[�T\��HnO�iJ|*�g��H�V^�"G�m��nad�j��|��aO'�E/ӥE6@��ɛU�T&��d��s7uv���3�v,��DN�7�C{�M��l�/f�o�����5�eT&�I4o���8%����ڷ�/��$��:����k#�
��T3�?��-�w��ٞB���Ԣ�h?�;˒��\U�VP��T�I�B<�o}E��g�G+�, ��=�%8-Ħ5�q���
�)���+
,c?�;��Q	4�;�aR����%pk�"�����H��AP�dA�^�̝m;���z��(e!�v�I����ET�U��u-w�*B�E����-P(�F��<��V·���)[�p* �M���e�#a-��Ӌ�n��@"�c�s?]�v9t^:��=�4��*>�?���_X.�H����Ϗ&�BvA��\��9�9d3z
�|c��&u�'J�j'�^�@�2z�8��𷚮$��1?�l3�"�Go7_�/��2:>�ѯ!�T�Kg]�ﷻh �����tGN�{m��?uq��IS3|6,*I��YW��?n���� ����]����m��I�^��O�kn�l��@V1fq�1CL�o�GN5# k޲�ڲ�>��Ԏo�z�W����U�Q��4��X~B�����?�I�'�e���[8�+W�Y�hF�@����<�d;�u��yV;�t����	Rr��;�U���ޯ��\,�=☔��c&�v7�� �n��g�BJ7���q�O�Ƅ�GG#!�����%`>��`���ي��S����oc;��a
�c������_�Ca+5n��'�>쀆Y��[h�o�C�]�v���j��'�@F:B��@�n�|�D�����!���OE�>�Rz0r���(I%���(�//��O��kd7 ��܇�i�z/�)�K��|�J�p��f�hE6+�z?�����v�]���2LP��F�B2��O�a���8�\o%�w��E��^���o%
�{����M^��&%02�}����m�x�T��Pb���*f�陴A�ۄQ��{~sG��K��4+g�~Y&�l5����bp���@)�� �%ChOx���.v~��p�'4��r�8�_Y�)��ׯQ� c7����r����{Q��}�f��q�f�N�Hv����8q�F�_�aT���-7���6�rO톡h��d5.إ�}�C]V䬤M���1].�i�!��!:-���V )���B�I<B����ϔiW�r<xw'�}*z�F�[؟�}A� f��ZbPm�p	^Z���+*��m���S��5S�8�e�̔����j�̇�V�m�dz }F�O���0����rB���P�������0���sd����QT�s����]f��Kst^:s�S�n����.�ɋ�<�x̼:��P�>���UV2�K)rDh��~G��;�ܡ���#��0���y���Z�nu�+ҚG�|=��Q7DɔN0������c1�g����a߬~'[+��y��Զ�hR_&P����y�(YI�K���];�y4.$Je���Y���9B�":�Mvs���m��o�p����hcn�JW៲�Mo;�(�a�^�
���ƣS�YIɸA���N�Մn�a���i�)��'ҿ�����m[�yɰV��p4Lg���D^$n�r>-�ԟ�t}���1=������#�$&�����EEM�Nuz�'c3��t��5TP��r�E�%������?N�[���#���Y��E�u�[ws�9�4�8W�B�HRo3�'枫|'����$脆���4�2NY.+����;E�!���	~�Ŕ��p�jBq"��^r3l�#S�����>H<j�f����5���C/1;�1}Q��h�gI�ƛP�Ԋ=W�,��Xʹ����9mG!,�l���U�εnJ#�Ԣ$�Ъ�mJ��![$rW8����k�[\A%��e�2���d���X�w�#��6���ʋzQlx~ރ����m�}y�ý0�`�/�d�)�w�˲���"j,�*Ѻ���@,Hw��`{�#ܪ�Q0��k�9>]��vmb�����u��8����Q�d4�;Q=�}mh�L*�)3�Ҷ���Y`�هF�hv��[���>��,،���$r���y\��l9&V�S/�"�@;�9'�jF1��TX�Yu���fe7�П
j�SY&�)k�M�������r��;]`DhM��G�p.�����n�Y���O`˃�/��P�)��ܰ�~'�0�"�"ob�2��~Hϖw���C�rUw���`�R�Ю��Rhk��&S8���ym�����u�ܲ�Ɋ�&��oq�^�FJ�L-`�9跼7W|��^(��D�K�p��^��NxH�S���|���!�5�_4W��q�W�e��\�E�a,�ޚr������)�6ex���Nn�$���LoZ;���~�3-���ׯ�I&�D�<O��	���9A���Z��e<���&㲪9y������9JtP<Pj��^������S!�ȟEvG{��0��%�Oj�O.��cÌ�܏`���c8g���/)�o����-#�ռ��I����}~�����Nt��!�\3_�c3�{�nr���-����:�P��C������q-�ޕ��+U�ɠ�$d�W�!�6l
d�I��.�1��|G5����E�-eƳ'*<�\L�����y�o��YO����n0��������N�6�^��>��oǨ�$��`�F��m[<Kǐ0�C5�Y��qP,h���׸E �9&5[⃽�-��z �nƫ!5��I�󿚋bW��c�%���$e�a|����[{� ]�9�
ٮ�����4��Gׁ�x��+,c[}RZG����s+���7%9DPW
vwdm�rt_8u+~���Q_�o���@{}����[��Z^Kz3rM���n�&%�PZ�?]g���a8��&.����w$22�π��� ���>A����y�"�%=����b�����%������|~�ES�t�'��w�[��:��H���W�U.��k*�tϱ;���s��Hǎ����5�yC�(D�W1]�Ծ����y��W�&����'�p�\�V��5W��⥞��I��S2��w��V�����)H�n�
��n�U����D�%�B�İ��Ӥ�DH}G3��ϋ
+��B���)Tcqyɨ�ޡ�;.�=���@��:�a箌 B��hz��~��PRf�M�j�g�HXf��!R�l����d��ۉ�(K��Ω�p��%a0�����\x�e� ԍ�D�!��G ��y%����wp�!#1��,�PrЏݤ��)gI5S���?/1�C��1Na=gE��O5
u��<?I�KM~�� ��(ޫ��7���A��9���[��y��Bj9@ݝHʁ�ݘ(��6�`�W$5r��ڗL,�������"��^!�ld��_-;�)u���R�N}B�t��8���lfh
��,+Z�r�C����w+t;�ZM���}�2����E��Q��:H.��Eo?j���˛�?�6ʻV�vmg����=�r�f���k�-��s��QU�F���/�I�4�M�@g�\`�
'�9��^����d���`�ڶ�4��x\��o�Yf�GR?���L�6W��Q辨X��W6�Ym�	����O�)�a�G��R����X���h4��(b�2i�&ȑ:� �%�8b[}-2n_d�, U�'�!��7�?�h��)�ux1q�L�{?�Cij�QÍ�b�� (�{�����M�����ft��ɍ@�4eX��� ��4�	Li�k(��L�	����As�=IK_�ˍ��@]w���;J$A1k�Jn}AG�g����#q�=I[�{t*â�dvJ���"U��&S����Ҡ���獄7|6�Q�EU�
���#�U�Si}�0�jͳ��-ob�Dw|�߮�w:�2�qJD��ק�:��Ěd����k�L�䓱��z�"�	`�V;+MO����I�p��Z��3E���k��B�RL�݉�z�4r�?u
^����0��G���&蝁��LX1��qY��M�o1� ��v�T�S�����}��Eҧ�B������/�O����Y�a=ӀSl(Gj�c�2u�҈W�Eݖ��*��v"ˉ�C�ȇ�=L���ް��s�ztt�>��U� n�f����ܵ��w�����#�+$��ͩ} ����J�z�ݷ6}^��g�����|�z�����������F���[������i���D�]Mn����C�2"^�Z���E3X?G����r�r��V�-C�,��M:�j��Cۨ�������D:a�w�&����(�����{Ѫg4�۷o�Z�%C"��ѓ�[������O�Y8/3a �Ed�����T%�����¥غ:��.�O��w0�7��$���S҂�,��*��-޷Vs��/uJ���`�4`��(��@�5s�n'�.�ٜ����ιG�����9�Z��n�����=�����Wȫ9yq�<�~bI�05�>���0|�E�he�a����\|���mH\E�����\��2k�':����"o�U��]�<�����3�da�� �B������l��o�#�:Q��ݍ�-C���M:)��F����NH���t7��	Y�`�IC���l����
F^ ���VE$��}���~����KKoG����8m�����^�X*���~9��l��i�%OT{ E�������l;EiHƸ���%��S�D��}���ζ�� �0�
���W�(��N�BV����a��"3j��s%���{=���j��93�_����@߸I�%�yaM�����T�|�2Ly�i�)7��/��5II� �6YO�h�#/���	��>!2ͶӲG���ne	|?�1͎��U4��NXK����5���3h�G�:��u+$�6��Bs�u� Jn��"Ϫ:@�t>g����ܼb��x�_ấe��/��N-@���RM�ސ<���ϋ(m
1ys�a�%B>KtT4p=wv/8���)˭n/^�l�%��e��X��]vkf�i�zs=����h7m�xJqZ��w��B�b����j�^^=>C��sS�W�%�٬����6ߗ�Z)Եŏ(�/9����̔���|�:���u���΅��GA?��tAw�,�~�5��� ��Q)���58��[֬�<hJ�$�9w �gcH[�ܸ�:�U����Ĺ����[�jDRP�O j�ObZ� �X-��x�\g��s6V�����k��!�v�Ꮊ!�桠�r���-���B��@��(16��eLu@4�h�����^Y�j�&[�TbR�0�<��
�B]�{w��f�+k`�wr�sb���}�b7�ҥN(	ouyl��~8b�m���t�n��O!]au�z��j*^�f��TT��zrH�64
i&�����P�r�SfӂO6�\B�����}>!nYf��
��+���΍I�9��B��;J�Rh��6�i�s�/p+��U^�Sd���kt����曈;�0�J �1$cα��o�G�V����*������
�MA��xD�|0��(K��4���2���V�â�|�?x�rz�:}����+·,)}��]V��#-a��!�@[��ѿ1��o��K #I��d���-+�t�[��}���IR%u,����O!���(�>�e����>o[J2oI�U�U��H�uI�{d�֦��_�<JC�MYw�#ALh�\?�E;(N�k���j�\�h^�QY�����0�:��A?�����d8?s���=5K<}dlG�9�1Cj�㈋����͒8��q�3���QT9`��n 2���2�:�����O�9�W��k�1� .Qv��IW����gX��n��^��m�h4���,s7��w����~�=�
,���4T��N"x����]��F��:!��W�'a6�ler�צ���{�5��-)��8��U��c��v��x��E}m�b4"(���p�(KfiBWdH`�A@���W0��G�Mׅ��]n3�E�����R:��0���a<�Wr�p7�'��\��Q���Gs*,L�r[f�#��9��NGnΠ� ���y�6[�6�[����&� �*C�۹4B#7�?�D�[å��,��<�m/�&	�JWu�n��uD	�R��@�(�ö�6�Q�p������%�)"��<��-Ӱd�.�����R5��&3c$�>�.�I���"֭�VPD(v�Ȗd�L���7(,�	�k�}�Gخ]̪"(�9$r���Ϡ�
`�D�R� �]Uq�X�0Hg�}wr|��/���|���-gM�y�4���P?.�af��^������""�<=g���}�:L��׃�,5��
|�tК��Ͷ�KWE��ep��ז!y��S0%�f��H���_�4;�,<�?@<nf���;;i�YH;zT+��^ht��zG�o@t� s�b��!ˣmJg�[ /����fx;��F8�0����]�:<���a{��N�:���׬�_|?�@3���.f����5�ZRF-�md��7����W{����*48H<�2�c����N�G�
�j�D�-C򔛼_ُJ'�6��J���>1����&�?�G�E���_��*'5�,���aO�dm\�`��g���T�B�?њ�;��
ď��FA�#.lDa�����0�pR�ʗn��_�x�Or�,�j0q��B>��6zye"ϗ=����~�?�f��;@E�����	��R,H�HT�P�:̅��1>S`���m��(��I�(�^<kEXZ�B�]���g��(�5�vvy��BOVe�n�Q��Ut�e��oYؓ�Ygƥ��+�"B5TR��^4P3����p��%^��~�5̎+�~���P����x�������a)@P�kNQ�\<�;�������w�%�M�RT?ᣧ߁���J8cV<�x�yZ�Hg���~)�7�+��A7������%A����s�p91�a�D��53:�/��s0�&�ￒ�SUγ�(_�B{����N���Z�یL@	 Dv����ݫ�u��a����6��!��+v�Z�Yֵ$4Q��B�!��:ð�J�܉9��Z^�d9��2�p,y|jD�3&�F��n�,�
�Dș����h��3�\[�LAX�>�RИ���q�%[p9=9��Qp�A��ׯ�8���W=MD2%Lɐ�ń�/~�@��I�b�A����n5��x*4W�j��3�yO#�OB���1������_
�Ih-��0��V)-v�e�iy����+4c����5����A��H/Q�9���,Uxjj�tz2rc6��I���e}I�A{@]�|C"4�0��$�Y��5�icjZ�y��Kj�k�/J�hہ�d�*`�M�}?_ �8�$��X�$��?� ��`��jz܋�`#v0,�H�R���j��=�86n�G֕|�U�#*�`��=ZA�y-6]y�a��\4^���.^]T޸�9��*8ښ ��}l2�撞t�[�1�ogׇͣ���r�+[�J�o�dA���:���q���$�)�(�����R�Ӏ����z.��%��D�����^E���x�ʩ˞���F�14c�D4�+;�:�9;�x!qUɈ�wz3��I���|���A)���8P��L��`��At�����b��(�)�j�Z6$s��nh�~��㺉�đ)�,�ɽy�n�����KQ�(�e�J�i�ޔ7v�L�B��^���k���% ~Ɂ���)L���y�1@ʴ�}M]fF�#|�mG�^d�ьj�x&�l�3��$�1�MM��¡à�)�a��r�C~ ��1w�!fЍꖸ�.�c3r�#p���P�������g�W����q�Ɋu.�3vl�\���\�y�M2���(_9><*� /�h�f�B�cl@}��{���R��ib�f≹̩#���D1����'/� IIߟ�Y/t���=7�Q�<����y�ז�`l�^Z�^��F'Og�"�.R�J��D���Y�9rUP���=�
3G5fl,�z�
���A끌��A�|Ö2\\���N�l�C��F��5Jr�i\��׭�]T�6&�(�x��q�c&4A\D)�G,ۨ����f�n��Nt��^�"��Y��jk[�E鳝fi��C�ؾ���bjp1N�ܒU��b�jP I��k�_�O�Ң4 R���2��:q��*��UO�>�7�E��ɀ�A���j��W��m1�_}�W���>I<n�{�2~mm��^@@�S1I�2+�ϙj��d�Mtj�0o�|9�<	�L${oc��(^��eW`�K��ӃZOQe��V]��UV�R��<$�@����ĢY�X�Q�@�Z�{ni��2Uu�, N��9�U��;�?�@� ��Pm��,�E�;�V�g�������Y,���)R�����ߙi��XU�4�F-S��\
�a*Y�����gR�̺���������~��j��m� �O/��M�����D�eS��V9����5�ѣ�3=aD��lN\��|�b?qG�W���ti/���*(A�0ǔǤ-c�b�n��g�:� �W��3s��_�W����ëm=�iXN��ĜPU��4���hܥy��� LF�U�̿z���D7tT	{n�B�s� �&��͘d����=pU�(0�}Jɷ���͒Ͽ_�49lO�4𤮌tx�L��5U���?�r\YD�ҥ���c������w� �ƶ�[��_wѴ~�؂����Ro!�
?���[#u�Ѵ��}�¬jc[�qB����t��o��BƓ$����2�k]o�3�b�� �@�~v��c
�Q�wQ��7	Β����][���iU��Wc�5����cu�*\�,k��V3��+8z��=UR�į!�P�$@o�������N�h�@�����_��
������W-��B��J����w��	)z�N���y
҄
(Q��R�6F003/��MC���J<�t�:� ����J�����|��q�����0*=r���k����´�8o��a��L4�+r��|R����9�T�LQ��6��r�_�E<��������wO�(a��M��9vo9��v�Ի���X�B�f�����}ů(X���=��;|���Y��t��%�^�_�,��n�q������o�ݩu����%��m�!�?D^/��Hv���;��B�*�+��˝�n[`��DgL�艮ʪ�|Qa!�Z�gY��
>�$ʹ���`�J#W�}�X-��Lrމp|��x�c�=�*�\%?h~*�U�+�ϜjY�PK��pծ�^�[��%)_j4 OzvT��u�<��Z�F^q���^�28Ǌ1�N�+�8@�x�g�c˗#��:��V�mjn3��B�Y��Iz?CBR$4_!�.�ꞃ :ƀ�r��}ʟ�[���1�V.s�4c���w�G�ި$�z8@�]C�#��^�����F���B�ɫ�f�W@dͅ<_&~�w��G�<Jf�C*@�~	E9bj��t!J�3/</�cږMr(�p�E{Yk�vP�Իk�M��r���/[�Uv.7p��1e�c�Er�I�~��%�(.��*���l>�0�H +o&'�p���"�18õ_m��Ή� �$kf�d�������Ɔ��qo��i�N�[zω�w�����1 �Nm@�z�.����Ig��q*�A���0NWcYM�m���Ҥ�}�
�Rޫa>�(r(�lU���E�jNNA� �y� ��V�NV1fs� ���sS\�~b;�7�'�n�t�䎑xB{n��՞}e��P<��<S>��^�)=w�O�*�h���#&�2��$�x�����p8j�J�g-Ǘ�lp�k8Ȗ�<�UW��Lr޽��w��	�e��X�+�%ܑ��Rua Y]7
z#5���)Ve�q�'	뤾h���_qD������?<FM��pX>�U�T�X�a����.h�*��U�=}���0SOR��nJ/����gvxF�r�����k�i�/�J��u���.?2�ݹ��T�. e`%�7~Wł8�Ԗ�-	�[��b5��y��B���6���6}w��oA�P�)!�p�⋫�{�D����t'�]�  ��K�-���{?��Ojҡ�h>�n��f}fYx��ْR"^L,r|���p���g�>_�:���
T^ƢQ@�(G��������U�k��_�I�2���=K����^�Á9��/�_���p�3S���i=����y������x �f��şK��e��k�Z>"�ʚ����\Ac� �S�۳]�z�S�H' *���A�,*�l����Ǭr�\]C��T��|MS0�A��Y�aM���U��J���GYC��O>S�,"�/�N/���T}�F���s*�و7cVd��u�l�����UaoM�4S�-Ab�"Y��1m��B�Ӊ3�	~|`e2x����j���/4����]]�y���K��Ar��(����X�\8�o���~��|<�޽w��86�Z���_v&~֬�dUz���fM�|����%�Շ��7ZB����a�k���2NB֥U�d���v!�;9�%�f�%����"�"�v]�/�[)3n1���?�ޛG�=��)(�4��h�Ӡ��[��r�2�V�����!5{��y���d)|�j��B�Ł���΄}쀥X��
��|ڲ��>��t5�C̏_�9�I;���4���h��d�y)6~=��#�|.���-�r�< S�F"��{~p>
l�_�+[K[AóN[	f�5�ҍ��^5���x��W����ZK®T�:.lO��U�b���[YTb��`+6�뇨`�t�<=n,`Pl��gಡ����G�F��* @�ʫK�3�n"�ͤ��� \o��w���'p;�H�c.�S���sIlX^���y��0�/Z�-�X���߾�+�ғ�N�-�����:�Z,T�&� ��\�G:lw�+��\���
"�;��ؓ�f�9}Ǖ�s��t2`�*�[m�/�s�)�g�L\r���h$�U`���<�����3#�uς��2&�*������Di����
yO�V��#���Z��H������]���Y3�ZWU,�����5������q��bq�T�Uz�UPR�KX���$����~�A�<�g�ޘ�WS��\�^�׭E����  3�͂.^��~F~v	z�����_B�:�A|�k�#y�f6��il��}0Z(���tǹ�Q)�qM�9�iG�,�'*�E�Ft��壶�eL���_��c2����gJ�o��i̊�\���@1�H}\s�����k]*�.�7�m�r��I?�%ƍp�t�R��P�^I��l�X���'�/j����iK�w�5n�Y����i�Ԑ�h�rY��0�c�!0,�
��aw,V�s�r6q����yqI��8�!���\h��A�+�+��R"��i�w���':�e�udٛ
h�����e7ߟ>���L���q���k���d @h	9�ɉ[�e$H�cA��5�7�o� � ��w� �pǆE���	���؃��-��$5��r�[��or�2���(	�no�۝ȩ��^T�"[�n�_*$Wn.�1����)]hc ������.`k4�SԫZ��o#�X�a�CUFW��m尌��+�Յ�V�NԞ?��[��E����jq��=a�R�l���o����
}������<�#?��_�bmw�q
��9�<v���Ãz�ù!�!n��ؐ>*�\�9�>WR�kC��F�i2]�/�t	���yi��ꈏDT�/ׇ0�k�̞
6�<O��|����E�@Y��p�B�kYw��MX�)F,o��,���i���y&��o�����?�R��,=)6)�4�,{�;ʁ�G�e�H��	H���
�N�\c�bv��V=ZkJ�:�oc���[N�����b9�=��(
3��׎/v�����;����-�a���Nv�o����V;�kJ�v����#+�}V�r��4Dk�QG��^��$j
T':��v&)��*�K�Z?�K6l!b״;gT���p������ӗ�K~���B�z�X:��]ͬ��t�KV�5��,����� L{�o�G�����վ��Kd`V9ɯ�6GN)]%I��V��-F�Dت �hj.��UV�L��w���I0��d��i�}W4��"�L�4Pl�Vd���"�b�:p��UjJW@���u�Z�r��	;�A�Q�YY.�1�G�.��(.�5�[�Ij���9���=�@��%dG�e�P�]�(��֝	�������Y��`d �Zq�w�Ѓ��wN�8��r]�>�H�؆�� ��Q��lՓY����Pf�7�/>����B$¬m<"krg�N,��Ѭ�^17l�di����J��0Mf��׾:��	5���F|�}���fE��V���jo#QBMR���L��r���K���n?���u�
�M�1"ck�����nڿ�E�G�̗;�)xކ^�p�h"�n��}[z�V� �;����3pr���}?�S�sa
^�c�9�_�+ 3�m�,j�u<8����l��j�NQ��.vA��+IğJp4s�����4E��.w��ah%��b�ڻ� L�>Y�0�vW�km�,]A�G�()�u���<mn`ہ�~��#�ƣهW���|�!��JHX���x��P�������K.9=}4!1�B@�܋�GJ��^8sU����W���b��UM�ߟJ��{�}M�^Αدo� ����Ylx:(��W��&���Zi,�&��6~���(e�ߋ-G�oCϐ;u�铂�d��?�v<p%?ʐ@2Ux��9� �tϘ�v�P�Ǭ�'����d~y�������vUL�ȕw�ӹ��U̹q�0���l��M��w�w��{�h��ch��K�<�t�}A�r?�@�
� ��h���';K��|��sFרt��� ���v<Ň���\�o�����ۋ%��iY$&S��\�M�x���ޟ�YP�!�e&�X�\�Q+_:�/p��m�������FP5p����6�$�Փ�eS�`Y��u�텙�SѓU.ʏ+|�x�5R;�J���i8Ae}�F���fƜ�E��T_����;ࢧq6;h1c[�+��ɐ���Lt��|��~�TE�9�>uP��&8S	a��Ve�vEʼ�x:്
pw��qz�Ճn|b�vc��x���c�9�K)k�Ҥ"A(q��|:��3b�xA;_3Y��J�8�6���I�-��v��-�4�ح\�I!la�W�	�}���И p'�H��U�cf>����H��S��oMx�'-���~ �X���fg��4�8(�������x��r���[z�Njr=���F����P�+�B�� �� q����i5�v�Ngm����\�u����
$
~gmk��?�P�]q1�D+��0ܘ{lus:��<\���KJ�i�+�g��%=oF�u���В��$�����7!���""�j#��u��Kw��֍�!M�	F/| ��0���7�O}8m�8���
�&i̒h;T�v)|�t�M����ق�;�5Q��|Ѻ|u;���(*��AW%�����3`�ۜ3�o�t�r ���*7��;:|D=J�"|p�����Z��w�k�a��"o�!�d��CvT!3c{�<(N�wRU�䜈.GK�J�JbC9��=�'�̺�gb��������3@֚=}���l�F�VV q��1�3\��(:��j(�3�	!6y�3�vA(����\B�'�+LF{vӛ��/������Ha_D�	�Q.�r�,\z��B�;�����yUX4ES���-٫hT���?��~@2%Z��C�^f>�X��#�8�-�.�;������?�����Q
Ī���v�$�O���p�֏geg3��O�sGv��́_��^�X����`Yc�R��M�'ix���%�"��'&G!�³J46�ٸ�Z�a���{4a �n�K!^���6GuDG��� -Ϯ��.0�`;!an��Φ��3jɮ(I��������m�^�v�Rl� ������- 7����T����\5b�	�2�
P������+�3��T�U�/ʖD@���N��qv�2���� O7n�E�u� ��P����S���/�(4��b�x>�	�����-��v�z�@�wj�$��0���G�S��Gy����G�����++�+^B.x�����3OH�������&?uRv���th�/�L���nA%;�su��A���������pP�)N����)�j�p��xih�\6��4$g
��k�Ф7V��˙El�ha��9�Qo�o��	����c�X-\�L�U3X�*���4��$Q	�SlV��%���Y 7��������� ��ݝa�'#-�c�.���mm!N����m�S������~�j���HZ���	$�s-���z�����2��ʞ��)��h��4Mc�#�˖�)����-�H�3�a���;���ʒ0 �����YK#n�8R��<>�qt��g��v*��K������ݙX�̗��� �=��x����k0jO�~��S��Fp���ň �\J�
����'�/��ܔ&tM8G��zH���[/���<X��6gu�K���U���g]UP�L"x��$[�z��j��y�S���V�ۂ�W)�Y�?ِG�]��[8^>6�]jބ>��cMX����r�Cd�
X`Um�yo�]�:$�/��ډ�ʁM�#^�'���g�E�f�Yt�d�OY��VW[�3�J�J�papR�ɟ�U�D�뙍��cRT���(��P��Uײ�@��8�h���qs)�\�>A�@/{}1'v��Q�Rb1���{n����m�������>=x���g����-�����ٸ/u�����0V��W���:W��n�n��uƾ@���NmF���!��,,�]LZ�6�!p�?@n<#}��9"#1��5b�T�l=F> ���;Ͱ�M N��Ϻ�#F�u�_��p�e��A%*L���O�ԫi��32tý N$s�ө��4z3$|��-�?��.}y�)
��x-Ǯ+��P���~6�s/�03rQ?c��gC�Y@+\aH�n;���q�;Ȟ]T���{J΁h�<6�xۑ��%�����[q��
.��Һ��L��k�6��6���`&����~�-%.ߵ.���/	?2�b��^09Q0mu�(3�E@�����Q[��cl�͌�_���J�9�[$t�7�A��6�,ak,���ډ.��#��;��D��Y��%F�_$/���,X\h��w��e�]|p��<G����u�5��}��ϐ��~:����☺˻�$eI�9��-���N����}ş[̞�
[���;����[�|Ct5��4Tv�r\[��o�_H�l�Ev/��?��D 5�W�ت��X<,� �V9�j�th�ST=9��ԛ9��He� N��*��9� Y+���c�xs9.� C(*�~�E
����ĕН|@��M���8~�CT����H�`Ք�}tǱ��!�S��y�o�f��|OJ��bz)af6�Tё������l��1m�C�0�de)Ԡ訸�>��V+04��S5�`�����v�UM�CSm�ړ¿����VNZ�A�jA�M���/����r`��%��=�w˘+w-踶�������˂T���TSO���[L�L����^�׾m=�#J�^�n��Ċ�O\�����D�ELA!� �Z��~�v8�D��\�����r};->��7�b`9]��hȐ�����>b�a6�3&״5]��]�t2��������_#7��o�5Z��?�d���1�k@%�	姇�B^D��bcb�������`g�>��{�7�T�3�_�Q�y�� є�*rS�{aH�(�*�� ��>
�v�I��~�/f�l�`o=��p��,��m�5�2|D�ň�-��z@���i�@iTw/袨*E�Иm�%�$�HG�3��5���I��
�K�>e���v0�M�>�=v1j��e-�U�*�B��nzH~ȝ����b�]��?�i�c�nj�ւO��f��~@�Kl��/6��qd%��m�7�Q�]i�S���x!e�N��a�	=)�.�Y�;�SUc��9����T�*�N���9$)VD0S-��7�A��Gn���Ow�Ѝt���rgI������@�zzE�M-����, !�k��ͨ�!mT�nk���8�O��O:��4�2�3�q5h3��o�wH�a���#����r���珴l�}���+��Å�+q:4 &iPD�Ub��p� L�~��5��(^�s�sC�t�pp��
�9�Ȋ�"C҆h��Wp,C�
��R[m�C�7F�Wd����U�-~�T�O1�6��-	��j��z�RX<�3�M�N
&�6��ڄ�1�B�n6<�
�͏�wpB=���j�S�H��s�T�)�1!M������`n�5~������?,��?1�*
E~���/{p)l�Zy-���ؘA�>����̀���/������'�_���R�z�rCãOqë"�o��s�֩_ID�N5�h{��"+g%UJ��iQ��>?iZL�(����z4�l�pƌ:s���d�0�?!��`��GC�*e�fc԰]���1g=�u�"3����h"3����]���k�5��:	��p�@#��+��N�w�5]��(�פ�X;*��گ����3�e�>ނ+m�S��)�����o�=�S'*G�y����ڬQU�r�Hp���>RR�J���@i�j�H
X~�q?D�[@�iZ��_�����Lܔ�v@�)��|Vi����W�����iU_z�� �P�5��t��*�BTJuXn�f�@>��Y��P��3�˯�q�}�T"?(6؟���	��skrU�>g�98K��BO��} ��ba$����\�}{�q㩉VM���]4Ҹ8��-k�m��ԉfj�X&WHb1�*��ms��ͬ�V?���u6ISC�Tz���5Ň�1������؂/j�>��z/���\�j�W5o���s6�6�b��;Wm������%�ތ2����}�8��V)^������?Dm�EY��;%"HV��&�Ѻ^eg��((Y3�ƾM��;��8����{v/Y��rh�
mKS_��{lϲynE��l��ٷE5*b��=��7��v{cSf-|���)��p11S�m�y���>$��o�/jjs�)&N�� �Qf(0'a�a^m,j�^�KH���>DK�`-A&���V���P@s�~?
)`���~s�����ת�D`��Y@[�y}Ԡ�@��骪/e�� ��b�(���i�lH)���G����Կ�%�`��=�z��V������Zc�]Z���-�6�.S¿�՗wn��+��a\F-t5�]�~<�3n��{�ڍOA͡%Nk(���Qu�9����TU��7T�S�e֬`���
���iᬩ`�M�?F�.9��W���t
]��>8 G'P�j����.Vra��������ԑ������oq�G��;}� |*B�~U^���	Ł���}�JP<��<i�Z����X���)B������)�V6����Y;����>|0��J�n�v'-��c��HW�������&OX��7�Ot�b��	;�0
zKQ���!�7}Q)�/�/����nWs$���C��������A=�^��BH�ڿ��ӧ��j��JH�[ªr���Km�D�⥂L����j��tc#C���C[w�d���t�\�]�=/^���0]��>KbN:-�7����MKgޏ4�N��)� ͹@��
S��������3tm��QHB.��5��H�x���708��o�bJ�x	d��QѴ��;����C�Y���`P�|�l)�%�1��W�������`�w�׍�8�Ց�����٤�c���9����1�Ө�������)Et	����� jM�WF�G��d�0�Gģ�g���O@`ߘm���Ղe:�EL��-���T�J�2cnu*O\�=A�;(Jd��j�f��Ȥ>7�w�sh�K|gȢO�{��Pz�￴^/o�t��~� ���,ҥw]m��Yh��g���̰�1f�1�x�[_+���Ҷ�H�"�oy�Ɲ�.�1�^!W���
օ җ�"�E��T�>)��.�n%;�*��4kք%�k$��U�4Ku�|Z�J�7�j&��C�*�"+-`�XP��v2���Ǖ�)sr���������zI�/��J#��Y�����#|���J��[��W�ɕ)&sS��")sB�?�&�7ȹ�������0��L��������0
j�>��U���;v!�ܯF�/A�{X��4�Mo�RkP%c��yi��?�
 �4uH�xs��(P�j$=i$�4�:2�W'nq}�wn���ƠoJ�H�Q���:#k�}$C�3�Y��MK+y��c0]��3+i#ģ��;���N��def>a��3����u~�;���{&�z*xX)	A��z��eп�-?�LO��w�K)B���ᴼx2r��]
�Qh�U�g�R��m#r3�`�SI�G$�(���e�,el�����\��Qmi:^_�}��)I9$+U�����-��-@��/���,���p���3����5���D]�4n��Ŏ�1Y�?�X�3���Oo�9�3U��%&���ma'�^�T���Ǘli�Z�ܿi��t6f��	J�_���ɿ��[3��XF��-v&��&�k3}��������iWș"LG�Dv�
f��b@�-���i�tr�)b������s�5�%�e{1�B�̕p��������Ƿ�'0�ƪ�Ê����*����ާ�8��y�5����&�9���ny�wQĤ�UR��ط��N���n
8�I5���6���a���s��z�-�'F
��t)|@Jߗ�-o�D�r��X�$�L������h�O>�݄a�����l�A��{����y~ppe"��Jq���a�ju>���1�;9���ݳ)�ȯ��U�Y2�2���q�d�y��00�Vnŗ�(� �#��*a��8dAUU���f2�ܴB��_uꨄkW�}��[�_U��1q��#�]�଑�R���u|s�O�q����x}���)�'�+*@��/�vl����%���s��Ɛ;��a��a-�O�6X*�ý��E d���F�2ް��Ie@������|�B�H�j���=L0��K��a�Fj�=��h���G�:6 ���=�RB�Ҕ�sG2�B��p�ƶvN����=ۥ#�(i���o}�m��+ʲ��Xk��CZR��k�5i��U��9˩+��^��L� �x�.�
ܔ��Rw@➕��'�_ĲRE��%v6�Q���Վ+_�*4��%+i��A+�՗^݄�E��xI�ޥ��)�U����ǒ
�*؋�m���hR���2�B�Fx�W.=N��H���x�b�[���DjTbh���8W�%g�kB	��Q � ���5�FY�m�ML1#ط{�+�%��\�K�-�'�=����!c`L�i�?����!A7�To4/�ZA��u7?�~��<�����)��^pdwz�
+H���O�y�Hʛ\Gp"5wy�"tV���6�B�}i&��Q�]Rv�:C���Xa�1�q����k8ra���.^%N����3W�wO�����	&�^pѼ���K�[�+��U��R���Ñv�����Fh'�
bsamYW6.�$��4z6-Uv�Q��nƻ�,\�Yu;�#��[*5�G�����4vI��bׁ���	j�S��z�x��JD(W�HT�*�I��L�[Du�bA�J�|��V����%�e�E �2�o�zY�b���!���ì��\���Gg�[�}k`����&�(9e��	�ɠ������Aq�'�"S��klIDbš�L:ɶ�9
}[ 3 ��"�_��$[�/rl�_�1��7Ln�=n�Z�����ڢcǗ�g1�ɷX��u��`>�F��@\	�.���f�dET�կ�"[2İA	�Ud���S0�m��
���{�ZL2�b���>�zެ��_��F���XP	�K�O�W��Ϟ�P����=��>b|��Ɉ�t}�9߷��.4�ʞ7-�+=hlk]�W�{�z5��ӱ���b��������&m\"H�A��/ҧ���%�xG��M3Π�)��Ilc5��2�깥R��r���6���^���W$�D��nN�5�E���wX-�Hx��{1�a�bj�������W��f:@GW�?��������3����SO09�`pQ/L�?�	�F��M� �*)[jh��B�����S�g��w�;����9r[�C�bָd�B�-N�[T+c��c��,c)�OܳXhv�V�E8��[@��:����>�K�ekݐk|,~�I뮓-����o9P��a~�+�Q}�d`���~�<*�C�~*h�M�(��*�e�W�x��i.8uT;��]-���^����*���G+��;S�T�/���eD]C�O���^�&�Ea���U��7�`l�\2]��l���Iwe����iw�(��!dE1�3��󬲉=��@٦eѳf��RȌy'��C�������L�=-��-,��9�؞s�{���YXw4,�ߏډ�ѮG"0W�g��_��r����db
8�?���8C[3��ĸ����a���*��(��=���%��Wz:�#L]C���9JïD�EV&��~Ìl���)�N;�nc�<��At�@�d_h���.�9!t�}�|1^�����rW��`��j��_�G�"���zg��n�����գb�D����{D&T_N�E�<ћ�*/:X2=8�zO�S�e�^����#��q��X&^,YWs�,'���(	wc�[8���e8�a��'�����2r���-0G���+X��kӭ��2^H.�M�{�g7�4fv���{�7ZSaŲ|�xs�J���h�m�����`o��A��)
&�D����LP �.Ѣ�Ծ�	׌�h)y�9{�t{��v��;���V��<@��.0��S��u�CBr�����!w��a#}��'B+�~g�NP���w���?"�Aס�DI+S���� B�&6��p7�.���A3v�8C4��:�7�Y$2�`��T�r�^(��\��-fF@�q�(_�
�"�L��yC��?�;w�+�T7)�B�'e��a
�K��,r��u�pS����7��F����yk#B����LU{�򈞪t��٘����/����Ф�m6e8��Q�
A3�T�X}�!~c���x���/ʲ!H�p��~/ҍǢ�_��K�sx���;Yvz��N��p�^���`՝S��_��?Q�wjrN;&�_�`��Kdf������K�wxq�g�@\�?�%{OՇ�1:z}��2G��v�|m�:�E6����H��6J�=�9�	`^n
�7̛x���LoN�mA�HA�[�򜒆��rٺ0.F�_�;�Ō%-�|���@�Y�l��|�����@mХu�6%�{�n�:c������b�C�9F�G��)����)ğ�e��/�L��k���.odtb����V��פBf~𫏔��c���������I[���>����k����o���#�/�$gVܼ���S�`SBbn�֯�˫���,w�A���^�b�]"��j3�u:#h��l�������7�8����7�e�U9�H
趮,N~N�5���L�ap�+�vH��sG������S��DG�l.�k�o���,�DʸL���6`rZyBy�P���բ{ā����/�}�t)��L��_�
��u�ZB�U�d���a*=���ע�R�G��*'��۴I8�KTiR�3���h.��#�sED��^�%p	$��*Y���k���v��ɥt��a�Kc�.J����IL���O�$�n�|�� ����b)Z��fA$G~� ������}�/7TK���XWB�<�qNL{AU��=T��
��a�55���Ӝ�0�"��ű&̾{v[/S�2��@�E�˜�F߃6MVMf������z��p��b�[{t��>��q9���'����䷲��ɞ(Ml���_Rd"�6�R��^�+e�	��5�U�����/��C�S�vL?����G��A�h��W��]��pm��3���\�/��X�!����v�8N��M���1��AZ����
c���8��k!�|��k8�%�FF#��p�~��`=#5d���ul2j��M����A���<�B�J�ܞ��A�y�ٸ�3���hU髑�me����L*��ײHw�;.,/ud�����w�e2f-j�n�yK���@}�d���>��_�E�|���1�����yI�=4�J��	hs�k�+v���I����C`ʓ�l0�C�?�5��4�Fʂ� .�^G��u/��S/���6�*�*Z��z�O��"��~�\�K\f����4�@H�T��n��驳�9�}!Ӊ,s�rڶQ��O�e�
��Y���x|��|LWQ�e�pF;S*�z���+.|� {b�~�"�'��w�-,�C�ë�P*����2��Q�u�������AM�%B)�ɜ��fR�'P$5��%%�š��.Qa�jʟ��/fl�΂�w�� 6)��i��G�sL7a�45�� D�}(�'�]�m��D�$ا{���~�G����6jai��xS>x\�k��!
�U�w�b�@�n�~|�i#�`��{?�4=���������	�n�b�t�`֤�kЬ��3?{1I����i�UmU����;��ZK����$v\��IY��,�%��.}W�C��tH���j����><T}�V�ݮ�$���<�d��������ѽ����i�h4'��� ���8�s�+��u�ۥ9��)2%�B8�f6��)�d�2���?���Dw\��F;��]�y�}�s���
س #$�{g+����r��q�����^m���N���+_�|�@蘹�'�`�y6����8��W�7H�3�s-����f8�I��7��8�u��@�W�����w"w�{1cq�1t�lU�k&�	�N�Z?G�.�[=������-z����Ҙ�\�Ze�&����%�O˽|��3v&w�Ɯ�S���a^�ͥ�d�ar��U��̜t�����6�)��J��ri^A�c��>��j�&��rs�tI��ix��G���U ����y:��6 5��E�bs�����I�ǅ-�4��xS��D�6�Qb����*�Z��1y��=;c�	5s[������t����;�N����NRF�M�)���8����-� &�6`�m�&:�ł��K�L�9՛5�v
3l$qLYQ+jJ3�7a	ds�ӱMH$rL�jE�Z ���5��9�L\~\f��ڼ!��y���:��ܕ��k#5�
p�\(��j��,ݍ��C�ܳ`(eC�a�lh����T5����}��|e� ^���E^u��6lM�@�������4lk�UG&�4=����;6�3��`������)�wP4�bՏ�S0�Z���ן	�dB�w�o��	��x�\�q(��D.��XٚW������_���=[KñR(� ���]��J��������G��a�'�7��������L=�>yb�V�S���8���䌲W���J�W�P=���*�B�0��=��F���d5k3�m��O��̒��h�i�d4 ���?�c1ۿ��_4*=��2�w��/�I�0�٢;bZ�j�ȭX��U���$�^
$:K�PjE��"��!�P��L}�L!mޠ|]��9oB
#��RBmөJr��̐�	d�P�"px�V)�~	e!����aN�K��P�C�%b�l&F"<�HE�8�Z[���kW)+��V	f�q���u�Ԣ	W>D(~.����d6Vp��߻��>�> �L���
')�`C4�:�ϫ/��h$#���&�X��@���(���[V�Dh 14�]��c��=p������٩�b��Yd�⏤�!�I�=n8�p�C�/�б	:�n�U���;v%9+1K���O?˴���l�w���-�V�/��>�(�8�k�t'�����L�eP��3�����<�1�ӡ��6�Y�0�����g���ӕ�L���!��2ycy�y����AR촔��b�,a�]�	�j�"�kE{��xK�[�&����~*2� �1ٟ"�4[m�H8	qS�fy��#�eY2�1\�f(�$�ե��q�|-�+��q�WoSm��P��/3<i����o�|U�7�i�fĦbH�B�#���  Q���\.�"2��Nӗ�pc���獧�b&��܃�;Z'�S6r��-��X+B^Q7.����]9gq
q�.�Z9B�UCP۞�;?����ڂ�`1�wz�Lҏz���>�<B�"�1#n��R��ӏ֓���N�@a�`�~�C'TL�M���B�>YĽR� �1��W����~�����S��dF�ez0r�ۭ�����$u\k�;�ƈI�����L_�G�,+ۜB��!�q��W-%�yi�Pg5�� k�D�dr\Q�;[�Z��8����߳�$64OȽK���0eJ���p$8�R2������,�oaT��	�)��N �?�����v���Y�ߗp�++�y�˷�8��X�6P��PMQ_��G�g0*�K �c,fP�!_�h�Q�gm3��a�-n�Bv�Zwv���m�c�;�A\�f{���a�R�]�����!�0n������w�����<�A����s�aV*��YC
��X���mq����j#�<�`�s��[�����
T��/(�t�dIIZJ����0��kcMV��gIK�����,V���_$�ŘϨ�8���?���RN3D�{�Ԧ��WWDL/Ƕ���s�]��W2�Ù�T��D|�|�fIh�c��rf��C1ږ���}~IXs���'cvm�Y���.�� �X֔��v�:�~�z�I۫�<ָ�-�.�O	��V��"����Ք�{V��#H6�1���M���B;�p}����,#�R��a�ڡ��E��[1�83*���]�f���.5c	R��|űԡ���/8�x�i����g���D��:(�X�uU�ʀ9�Yz���LN[�qh�䌇:����PH����J�['ꮉF�tS���G[z���c�?�޸��F2���?Q,�� ��_Dr�H��i�<ksͺ v�\k�&���eF�s��n��
��t
��誕z�Ka�mh-mɥ�R\:��o�� �$�O9��!{� �i���cB�lf�/�K�.^�2 ��*y�G����TU�2�%хpг�Y\��m���O!u�:~%.f�d��ye>�"��Jt������.���F�?���"u�Q�M��ћׇf�9h������%����w�Ѹ��W�}	b
U�\��2�_l{�g��QqL\�*К�ڃr�Sl�	��D{�dN�ڼ��J�آWR�QG@�3�}f�o����qO�p4n>y]<��M��˼<�&!�_g���(��R_�%���ǹ;�Rj1�Rdӡ)-e%�7>|��,��;/�j���m��!�r'�ܝ;4ܦ�S��"Sֱʮ1��
W�l�:����l�QC�0���%Pa�j�����}�?oS�@����������Ñ���$d���D�b�Fꓚa^ ;�2( ��G���j�؋�O��`�U�QX�(W�*��e����|��,C���*��X'�w�+5Lm#>9��p7�k���⫄\	���e�0�sYgZ�������
1���C�.(��h7��R��@!����#�~�0.������.���d1ꦏ)���O͖�����n����Mq�s��91�}����E��I8����������"0�|ry�s.�zގ�мёe���a��r��z���͑n|����% +���x�>X1�Z3�X�_��g����8�p�8���p/n�ŋ�sꢹ;Mb���n��oϚ$���R����jYB�*&�r�����,�؁d�
��
�������
��6�jna�����d��q'Pf����=���d؉���-�b�	��O�^�6C��L�rt���B�K��Ოzdv9x;6N��(���Ŷ��92��||�u�*�!��sk�|�J9��d�pn�-�܆M��="4�  o�U�'�<�[#pNL^W(I���3��n;��O��Q�\�Kך�v]��m�K�#A�\y�C*8o���2o�wr!�~xT]_y,7�cm�t��v�>?�^��O�,�]�׽P���)��^�g9�#��x��C�+׀F6����O����p�y� �UfW#��_I��ܰ��Q�ټe&�qǧl��BQ��=�x�F7��}|X%�&�o`�����`.Nor�<.@F`66�v�<�L�d�R�2s��S-�&N��u̴oʜ�����G�y��W��2��V��5Yg���մ��	���A�hfK!%%:US�
��@Wc�����zd�/Qea��+Pb��X_*4�s�I�.����w]����e���m���_�JR��D%�e��ť	z�](w��m�5���^uN��<;��P�vw�A�����&��(��M�R�\��fM�����ըPV�i�Ԇ֤��� ��.�#+;6(;#Y4e�p�b֡Q�m�1���4~��"i(������X���P��Ի#�2���M����Shn��"���&
\WOÐ����ǎj=@���Kd�����%Slzh٩�4�.[x���zv�o��1o�&B���Q���+��I�����Kp��-1˼��@_�ax��7ؘ��/}aQ��R��I�pW�MH�2��G���Rg�tE�JGԓ����@�f����������z;i�G%~[)�p���?iY��WA���yE�
��%��T̘Ⱔ��)C'�BP��[�Q/�o9��-A�.zG�UQ����b�g�)��ic�O���R_4G�/�7�{�#��8kf�7�9�k��-j|����g���[��Ȁӵ���elI��G�&�(��fi'$e+ݘF��[Υ��`�>���f�]���ɑ�����Rx��[�-=� >~��+�F��X�����(
�KkJR�	�Mk��hX�^���qj�"��(��Z����"&�X@ƌV�I��/���ծڕ��l5�0	7��?R�˄�$�[7o��!�A�͠Sh,ﶰ�I���&��F�ޖ����V��5p4��0:��]�UܿJ R�vrs]��h3��+0��@���&�ۻ;��z~�o��L�$�f�^|Р��`.Rs�e.��_bd�^�f��#�PN��?g�ö�_}QM��7N���:4s+];S����gd���椺�����Ch�C�Չ_J=1jz-xe5�6��<�&�c��L0	ah�/���'>���`+������Ԃ���>3�r�7�� ��WD��.�k?�	����m��W�C�2uG�H�)��I�J.2u�����r۪
k�J�/iM����g/p\�K���������b_<��m�H=��������2Qmׅ d�>��?��t����\:YkJnѕ+PN���S霅k?�aə��4"���Yo1�Hb��h��V�V���B7l�5��7�𙽠iFqΖ��� ��@�U��p@^��?�����*��AמP�-'��:yc��^<��/��fe��>���D���Uʴ�F�͑޺{I}1Rf�X�Ħ� zՖ�N����j�l�ʹ�����|�d9����"��0��&�\�	�'��"��
���Qd~ޡgx��,�nث5l��`ܠ��u�0 =�^�jGB���ލ�c3�jK{+������ ��?V�UDȾ��Ƌ�(�l]?������l�hVU6h4/1+2ލ�x��K���Nй���5y'%��;��71��C����1�1�_]M��2��=�T@RC�_V��<a�c��);�+o��i���ܞ�!��%�0IocI>��y~�H�_K��VB����@�e�N���T�����Z^��Z��C݅�]i�.�|��vf1Nށ��=Ӈ�G��"݇���S#P�Y)gۃ������K��TG��wsS
�Y7#U��(�W��F����>�6?!u�7�U)���Jrfc�N��^b;�9	�_�]N)�$�u���~��Ę|�H+H�5?���,Q�jrYD�{�k��s�����ms�F15g�N��RmBfpKŏ�`��]7�F�d�)���Ą�p����C���KVn&"@#4D�F�η�e]g�|������DeP�2N���^�A�j�NE�P����=����*J�ʒ!��sI"'����fn���w�}^*���k� �m�E�� �uMÕ`ħ������sC?�\�+E�b�6j�MJ��y��	�5j�|�hn(H��k��+V[eQu�J0�'�E��'�wSs�z��UX�i�n�<���{�V5sA�9h yn�GAc���'��u%���,��N�{�TJ�Ƌ/[�5FE�x����*<�3�w���:`o��B���Bu���W��٩<���߈�B�qㄠi��զ�cR�QѪ?����u��ɯ���Ar�=�v=�76	. �/|�ZP��Ա ��š�	�3F�ն~554��D���n���E����v�+���U�w�!����p�����K)�ο�F��:-i��ɸ�ow~��~�Cv�̙��C'��^�l�^d0���%�sE
>_#�\F2��=4���i��
����+Oh�Sa�q͞���r�54��%%���1�(��4Ό�1�7}|ЏE��=)��Q�j]P&o�ƛ��%��DUK��%?O�py��5�������p�D���p17 W�3����ɋ�5�i��I�u���Jδ3t�[-�Ï�#.G���ni*�T�#H�9Q�f�j�6"������-F�{��t���ձ��۳̿�U�Cޛ>�q9����?��g�0�p��iT�Q�ꎰ��J�&�:�&�<f�(i�	�^�~K2m��W���ڞޝ�%���EE6Dw��+�8�z��}�R�.9��q���g>`��h(
�m%�������?G��;�eJ`8�w?Z����S>�E�7g����Y/�"Xk�1U�E�J�����F�Z�%�Tk��e�u���X[��̜mM����y"Ƽ�A6�f�¬T� '�@�(�ٔ��s-���ш��#��+�X1�e�<K#�4ҥ���n��)�ά\{C=)�;Q�h������,��?N<�X�4�Z��+�T�u8����!//[ǃ9��)}|��<��Nm}�Q�n�a����B�qB&7�d���m9M&YF��7Y���� HA������ݓȫf:'���ɭ^\��h;q�Yy�s1kU�ER����Fs��ȅL�U�*�'Mg�%����TF�Fs�Eo}	,��~97m��Ԟ�VB��\Y�j���1�ic�լ���Rst��ucP��)��q79[k���:���:VP��1�q[���0ء\p�Qf[��U���DF"P�R��>n<jN��Q<��R���4����@6�/�w���P@<z��%�|���%�}5�
{�/�{�d�l>L��C���wCI���_Z7��PB�	;O�N0����T߅�!��sS��ݓ�
!�࢙�5�%�wy]vd��'��s�u��x����֧��|}��0+�Q���q�fa�>�z�I��u�$Gˇ�~bN�����#�@9?b;��@��]&�j����uR�	7��hlX��M�U��^������lu�#wţ�F�WyDLW�N_���!��@�2{=n ��x��M��	�<٦�D���'�(�Q8��[\���Pz%�ѕ��܋��Zܕ���ne�6�ũ�|᭝��g�f��~C���i�(6Y��⒍I�4��4���8oc��R}�����3��a�m=b����k�W �����qb�oƱo０�����|$@�4BC's���a[}*!=�>4Š�1^*�q��h�*�lu�B�4ڦ2�����Y��qF�qN�B`s=L����LD*����k5���ɶ���b�-��.M�/c�e�2Z�(훬��[�67��a��Mk��3��w�����-���"��u �MlQ����/�Ӊ��×���#�u^�u<\�!iK�7�F��{Pf�%ȱX��yg�+�\.)M��/5�:��a�1|�d��?���#�2���=/��jU�2�C%�G�.�v�%�`��rـ�QC�e�ط�{#�}�0���z�����ĸC�@�~1#�SI6h��;3S��DS�v�� �ۻ��ϯ�D�:�$��hs�ۃ��Ϻ�����V���siT�X]�-��c�:�y���s��s4�m{��V����gIn,���q&��2N�-��jH�daܨGf#~>Ս�A.{о����� K7��0ܯt���
�]k;?�!��s��<��[���*8�U@�g0u�&�B*~�k]�w�ʿJVJN���!Z��^2��Z��b>��-����`Kw�E�s�Y<�n���.NS:�S�������Rѥk�����Z�Nf�W��k Wv��'167МBJ�ʳK;\�_�&_��rע�"�&�׏ht�������^�'��`&���M4���,�b�V>�����3F� ��$�����cm�����\N��#����^˚�'g�n�CE��G��a���oXM�|����cv�������!6�%��t�<�QV�բ&%k��3̪� ����P�g�ƎrT>ɫګ�d�cg���4��y��.�h_����Յ�n{�i{I��Q�"��Eh�o��9�"���We�LV�J�.���K(�D�����o��IF��٢ڠ>%�eBq�:H��I��@AQ�c�x�@{������3�^X�.��k�s��2� <�p�ڧ�<c�0a+��ۙ��@&��eL%�î}Cp%��7���r����yQ�cra���c�{�8־edfĮ$W�̾(l��}o֑3X}�ھ�d)�t��,�LE��E���{��9��iVUf��݉�|1���#u�$��=�?Jҁ�	��;��<�
8�3bJJ���x5��B?��lQ͒��,J�|b��3Vp -?[���qх���#�A��!���w�Q��4O��q�t�T(��^U�M�[���L�r�lXr�0�&1Awp�nYj���a�����l'�m�YU\y�bd��AMJ�湂�ޙ]h���z9;t�U�����_��̇o��cc7�X��r v�L�L�<9�=��}�����$��M�dN�� ��%U��j�K��w䂸í D�ߐ8GJ𸗰In8^-P3C����_B�2�S�n�5,�~�����H�X��o���Ӳ=��b�Zq8m��"ʹ.wW�M��>��*���~N6bkH7L����-�Rs��� G� 3���b�~#��T�?(8<���5#�{$�	�4�x��խ�o��62���9o6%zw���󠝜�P�u�ъ��\���FSP"3��J��n�g���/-ա��4���*�ؾ�8�&�p��rU�ޙ���Bv�%�\���6?(����^a�[D9�.ԁ��K���ٍ�d[p�.��_�d�E�ݴor�HD"W�8#5L'�h0�z�|�|B$�} �5֠�8�*�.TB��.À��u�Kֵ 5c*��� �B���Nva�M�`r�����ɠ}uq���o�T)x��Hw@�{���N� �;�
K�K��9�}�������;�P��7���)��l�;P�	�t�r�Қ��s����[�z�Ru����UZ���Exδ�����g�&k�B���LEV�v�Ij	������WM�^���u�<@6�į���غ��Ĥ]X�w�>2t{vpg%%A���?���W(5��C�6!��M�^z�w���T��4��a-��h������=�8!�E������Fv��h�{.DQN���M ��}��<a���,s�`�%�p�_J�	z����D6�!�߫E���*����ANzYIM���uja��P1����ӕ�k!fy��C��]-��э�˚@�)(��Z��9'�L��k�ޯ��p�̀�_ҟ�8v���w�͜���&Y�>���{����5����EG��4/}���Ο}Íak���'�|� �2�dR8:�ޱ}�6Ꜥ(9�>#��Rյ.�Y���{�Ȓ��$����~����(�ؠ�E��U�om�q �1K1xO�nά���C�0��n������i���i���43�_>���x{�`�>s�_�.�,b�>D�8F�:��}D��0��k�0j�&�ÂIJh*5㪝wTF�O����� �u3�!�]�qҫ���Q�.�uˑ��ݙ�.=�w���j/�p=��f����:�Ξ0��bWtϏ�0/���j���������:Ǣ����uc�^�
���54��z�7}x�.���M=Py�!G�/�$�>|���k9���7s�����+S�|u�9!pI��I��[=$x
<Fj[`�"���u��<�߲���.fR�}�AD�Z���6�_S�O�t�ݔ�RU��ֲ��>��c��E���z�^sb��W��N�^`l���Ah(D���P>��ΐ�Q�[�7c6Pg����֏q�G+����<T<A��Ԅ?U��՝K�dY{r�[Q?��G�����a`h	����-��1��@I7�]*��z��\z5;��u 7�0�
Ah��R>�� >�yx���R��-�b3�3v!�W�ݹ�dz6���Y�90�kaHz�Ff��f�
{��D��!
�4I��'�l�7h���֎�X�6�����i��ӯ+G�%\�SElU��#����S{tG����C,0aZa��xd���5��{y�=��R`�x�>�P���x�ou>�9������|��pq�+VH����Zk��I"�=����6��`WU0d���=W>P|�wa��t�B�F��ٔ�� ��S@����3#}2��� 19b��(C&ENu���(H�-�`-��%4��
%���-�C�k
8U�c*b� �+⳴�����ަ^���}ѽ����ʚ�!O9�ɗM� �;#/��_tz�V�����(G$���䷤igr�㘙u�S<!�dh�4����b�u���4�.~߰R#F�Oޱbo{-�#n�Kj����JD�-����6�Y$����1,��A�f1I��ڀ[�4��XS&��Յh���b���9w][�$�]od��0��)C���,���w��ybU�&�^����C�N/��޸f � ��ߙv�?�}?�̣�v㧜E=n���HܯY�vHe�5g�n5pc��펩�쥘�L����Ͻ~	ˣ�O��G,���@�{�h_b�
�b��
1��c�B�d ���#��G���%�B�;ہ �AO�*ʔ������c�=4&G��b	9�r�\>V��ZQ�\��P)r̼5�v��W�n�B�#E7[�^o��?n��K��Z.?ك*���-bU��������݀q��A#��f_M=��4���ʹ�6�����a��BɄ���m]��������A����k�`Q�
�qw�B�E��a�d$��D:�PM"����Q�~��Tfq�P�%\#맹�jH���^A�\;\�ϟ��K{����p<�>d73�����0�
��C6G�|���g���0�Z�Mg����꯫�2������v��?a*#(=�N��������P��|���G �`�:�x�V�u��� J����h�����K��(���f���s0E�X=�╏_� ���D�+�[G45�BtK���%���H�4�&J�'��qWi�b��!rZ�Rrbk��.6�����῝�^�,pnsu�;Mƹ��
��%�R���a��B|�ۜ�7c�ܰM�ޏ�]v=^=����^"��c�)T���4V\=������6�&sq;�-�(�����锾S�)%�6j�lܸ�͢��^��Q휄��Q��w���`'Pi6W���9i@�ݩ���r7�0N���MHt_f�b�p�+K���ka��3%�.����H �NeH��]��8ϋf$�#0��R�ڦ�D��6�<F>w�'c?�8�bS�Je���i��ð�9���V�a&�D�{O���}9Gi�x��!ݎ�n�ܩ!�3��M�@m����GU�~��p@��l�&����&|��n���t��zS���Og�2h������+o"��rZ��:��,�<�$��9��+k�m��;Y�쌷sw���[��C~�X��6:.�9d�K�5C�jO��D^9��Ϫ7ӕ���K���ѵ˿B[<��'��MQI�ye\���S�JI���	���/�]��^{l� �v�_�{v��w(I��_0���1�e��Y�Z�~jF[J�)#���.�({��ޡ@�wp��G>Xߓ{|nV9U�°�@C���}�G�2ݲ0M�<�)ė�s��c�0W����WN��z1�C,K3φ�P�	i��WVJ^�}�K:�` �,��*s��+�η��2^���z�a��ڃO�נd��MB��x�4��5��y6ԑF|uZ�1�*�����v �yW��(�!D������4So�^�O>�Ŀm�o�"��*)��i�1�o��������N�RVJ��s���К?t������x���%'�������eD����Ԛؿ�~s������.K �4�s��=s�d��#��C�K���gv�	ȅuw%ۗ`���ӡ	.Edt��5�x|�W���,Umc�g;K@y1E��'�����8����������w���_?6�����0�;c��X�L���`�V�V�N�N�����|QM/O��� t����ƹ� k��7�q�_��'�S���<����K�.�6J}v��B�B�̪.�<��M��mq��0��xwj�@�;+eP���0I�/������I~��4��'�PXa:����7b�TM ;�`�Ifj�w�Ǡ� ��Ƅ$�0Y('�)ҍk.�@��K�D�5��wq3��zv�-%C�x�UX�ZLjm������IS�����v��b�d\��U�p�A@�U h��̀�W��-��Ǣ�$����N���c:^�M(��@8;ĥ%���;�޷�^,΀�7��j:�D�!x4�=a�0,��mjY�k��IIs��Q��2Xm�^���؎���:=ơ_��g�h_v%c�:��@ Eō�F�!)��4�Pl�.�8�TTܵ"�k���2R�ާCD�^�i曈���u3�k@��U&p{s���z�^ ����7$x�X�%%�-�����B�#:t��}Ǘ-����������"��Q��x<�>��F��[���BY��D��(`͢�WAK\�<�]��XT=�~�Ϩ�̑���s<-H"Ԣ��ъU�ڋ
Z}�=h��AcBU�E��J_�;�9�wu�uw!�߫�M��B�2��L���4�
��N�^3������eٰo ��0_&_麎�>�(Ut��R�	D3{ |�2���D"/Ro�����X3��g�O�Mv+��|�=��ѻ�b��ɡ���?B�J�q�Խ��͹H���k�(Y�`���} f��i���$3�k���Sf�X�ƣ��O�xLJV���h߂���� �^O��@��|�Iw}��Q�'��5��@3:���P����ǁo*�i��Fk
���x�&���m�jܬGH>mMY�CR��L�87�d+1�g��������@����	N��|����N$[3��ׅ��U���[�~x���~��@�������p�&��{Z
���l%�<VD_�y!�b�g���>ٰ��3 -�"A�0�qy�"�4z��b�ީeckmm��c2-����!�>C0����8}�
����%[q���>�QJ��O�Ҳ��%��]eA�(�5)����Rh���� �ߦ��?�?=��7i>EF�Ky���B�Q��C0�V��<���y�C�?d5�^\�-�sbخ����,B�J���&$��fs_�.�r�a�b�<#�CL���Y��;q�E�a�!��y �̮���>�d�Q�J[�|�c�R}(F�M>���3E��>���.Y�.�֨M�lv��&��_4�#��E��� ���F�ɣ@`-���h�6�,����G�L+~�H�7�Y�ppN�7�n���-x]&D��N�����?��;t����ZEX�*��\k��J�궞s��n���z�g�غ���	�~�ǭ�{*&?Oj����D4�mDH,�G$�N�0�c�
uQ���ݖ��B����3zr���o���Z�i�9Nt#��; 4|ƘmY�T="�e�9�ӱ��٢t��+��[p9E��k���2(�yF��e\�lIb�,&v�ư~$�&~���O���B;6�S�%��˩ux�&�L9��ʸv�.%g���wO'@�|�C��E'?����!����W���?��4�bk��E���Ҝt*����@Y���	�ì#��ͽ�>+ y�������6�<��i&#�߭�E�� f�r<Jc4�4��H�;�Q�%,����UR���q��H"D�U2J(�jlA��2q��)-dg��k�%�N!3�۾�����+ (VrdA/��拱�M���B#��u�l*� S;��Á<����.5���Z��P-����7T��¶eJ�;�Q�_V����"�a�t�h�9k-�:��}G������FdL3*����Rp��>t2W
��(�H�m{��:bF�ϒ�|$��r���(ƴg��D���km�:Uww���:@����hwDE*�rEy��&A��ĳ{3�0�=T����ϒl��g��t�H��6�H�Èv�fs�Jj'{�g��K`�p7����>�I���TN���BY�F������ڍ���#�o�RژS~vn-�����7������1 b���=�;�B����Zkg��\�O�؋tU 
m�Wr�[�g����qnl�L����Ȍ�$N���Dcs����/c�wӿ�=r�������9���tx]^�Oi*D���B�c���ȸ����BF
����v�&ف�s�����Ih��9�W7�n��������پ�X�r�wk"\x�>W5
�����"u�@�����M`���Q�Y�ll��aj�C�$:L�S|X���f�"
���_~j��W�_Iļ���M{Q�_e<�\?�|*�j+#�����������P��.0���+�z-�}^�y��UG�L�z�r�i��&]C9"���.�:�
n� B�@�������h�\���	��B�|�~(��>(�C��1x�a��^+�v~-I�^T����k�yj��a?z�K|ځX6��^����S�c�r{#�s�4*L/wd#:sG<��uY�'���0`��}�%���:	���J!2���7��W�w$g��ʋ!wc��Իp���v2\ ��$��p':�0b��s�/8K�V�! ,����Fcƃڭ?�1�Jr�9ƕ��:r���2�yB
�(��h�j'���𪯨!K.�ɻ�x�j��	�>��u�^���_sq�(���j@�6%����y�I�����l��W�kr��+������
d�q�(ht/�}��{U)?yY�=9�Q��NP-�A��<�J	���	���ɲ�1��z:��ҘO��tp�`$4����78Q]�ƭK}��	?�M�����c�>
AbB<c�l]R����9o3�;�S��e+!�@����5l�9*�^�aQwZ-��-��]:t��}���ne��S���7wm�.:�;4�O���XT���$i�;st�&�a������j0dfZJܹ�+��5�����ChwW���1�����s��&<0�8�vW�55�F����ۊ��\&���O-	�Xft��TIB��`d�sY�l��({J��P�_3�/���H�[r
�����.Y����.�%X� ��؛O����OFZ���\Ɗ[�*�L+x���jbܧ�<�r�;'����#��5 L���;�����=g���pB���ơz��ŨrOD5~��L��l�V����$�>��k�~��+�t�9��7����hDVT�_b�*��en-�<Ik���A�&��{j�J��2�j�|4���?s����/�?g6�~:��������Ԏz��I�~fj�����%@���n��h�5qW���+�c�������K�~s�����������Y�ϙҚj�n ��9�d����e��Ѿz���:��g�b�h�@>��v�\TҔ�b��k��_�ٻ|K|�ײ?�V��?�$�A�Q�@N�b����\�-�l(��j��L���^'p�XN�O���Pp[�Cp����<�@)�*�9�<�9x�,�k6���%%WM �L�@#Kд1ڲ<��>HJ�̒��TGFA���5����#��o�/G�	smW�]�{xL�[f��O�z9��#����IjE���z��@�%�}���̿�J��Ꚋ_|��R��]O2�bM�<_("��n����A2l���=��<&��"�G���Rݛ2t�7m_��
B��]��\j.����.=M���0�h��.��C�P-���>��8��-"�>1��x�xG�L�I=�m�k����z*�Ή��7�St�Ov��5 ��Qn`� �$V�h�{��������S �{��Yć`��������%Ĭ�0��k){�#1���
�{^�q�啉���I�HO�������C؜~�>s��P�#ަx�4��9����������$-(�,֠���5�A;z�nˍ/��^\#K�&32嶃r[�2�2t��}�X��TN�{�}��r*r=�� FT+%���s�3 �֠9���ݓ~��?�pK7��i�u��j�Vcr�/�|CM��A���ۋ���'���9.PL���b�L$�$��V��@�����2�8�LL��Q��O�UW1! T��'�!K ��Tri��X����ڏ|J����6�|.\fF�����8�tb��W���ʙh�� ቼÛ�G��;Rb��=�����F����Q��ۜ;��d��L�����K~�K�i;j�����X_{v+�����������r�]���ީT��a\h���N�����j	k�q�\	!�]*�� ��m�Dhe|)(����Mn�vj��TjT��z:~��K��k����z�Z����.qY��q�5�J�iJ>��t��F
���T� �@a�-v\c]��:��X����&��M�8�J�*���eY�Y���T�u�T�T�����0����k��dk����Q�RZ����˧�|��D�J<E��9�l���R���uў9e��'@���S�J�vŪ5+���w�z��<��O��;E+�v��zz�`&n��ox_�u�)�A����A��>��^���CRC��Od�U��'�l�I���9y�������gx���{�'n����)�M8��C�{ue��g �hR�C�N�T����.��!A�+���r�k�q-G]/�9��{Q��um�ڟ�!��㛲�w$�8m&�֧̎�����h5}�=�d!��H�>��/�Up66]��9��K��O`�( X��F�V�c�X��9+&�Qv��Ǘ��f�,��8�����_=S7kjC�Y���n��S��B���)x��dD�w���%Eu���b����d{=����>t���v(')�#ZT�\j�tOMbŀ"� \w�<�k;��֑V�'�,f�yY���7p�綕��L�%G��'��3_H�"ȧ�cH��QG%����$�'��j�#�U��o�v�w`/g�|8b�@��-��{�k�n:�������-.�&�Y"vz������������ys9���qq�/=�����-�p�Ƭ��N����!f Bi|O���X�|��N����p�
}�����0�1���HY0 �?]���)P�A4V���ժK�"K(>�5h�]�N�R�K��9k���=�W�ur2a�F���Miʗ���a��ʲ��T,K3)�ݰ�T���$k�ت�u��$����`�lf��ҊSY�2��u���bp�\��������9,^@E)�)+�hN�|��H�v �)QR���J��z4VA%b��ܚCcf�����*&�ۿt�x�mM�u�#��@�x�h��Ŭ}��װ�gx�D����qUB�	#On�p���;J9�ܼ�C�1ɓ$�pe�U�6��*��j�r��&'�&�S�q�H��F�*��u��p�v[�a��n�l!_���F��_�tL�tT�إ�륌���I8>�iv_g1�a|����"3f�#��(�q:�=p�&� �1W�xI���4��!�}i=(:�Q"�	9���Xǃ�Z4�3X�5��*������mqأ�*r�nbYW��R�~dv3F �/�cg���`솝~()���yoM��� "��)4��J�}�'��.C��c�L�x���%���g��뫖�R{x8 G~�"i��@N�ʍa���P䦙�a�=�咳?���;p}�6�w���Ti��x,-�W�����x,Z��v��e�laC��h�뭇�b�H�+1��L{I��V�
k-5���{9���a���@�=E#<�3e��k�;��T��ƴ�t[� b��N�3	���"5x��uݿIA�e�4Υzj�~c%n�����зXO0�Gf15<���j���!���℩��;.l4,�$~�¶[<�j�BF��L��� �i�e��CWgnj���@@���${��@$�K� o3�W�V�s��9�̯�>�Ъ8�-͞���e?�A���ج(*��@�o�N�w{�U��Z���D>Vt��2n�[�/�]���Ѽ��|蹕��~<�Wg������QTwإ��(�V�
�1J�+�f�= ,�@��NeGˆ��(���rn�:�c�Nr�Y�2�~P��Q̷����#���W.��AW+m�s����"^������jb�|"c��u�7�뙊�O7*0��\�:�gãa�7����VE=�{*�d�ϱ�F��~�2�N`i�����-�=�/�J��C㜤�U���[�'�5\�:Ȃa�L-yz�	Zp��&�m=dS�S����r+l������q,�<���0B�>����: �e[!Ƹ�,c��aA��m
.fz���E>��3yV��3��������v�o|2������H0vt뭘��4��l[���sR���@�
>�<O���Ʋ��T��ԭj�C��,�=��x�<:GB��鴝�y�2Mo�Ǉ/�`�cY*r��Vn�`����ٰ��Է�)�fNO[�ڨ��Y�Q���ˢ���m�Y�;	\�|ՠ���n��vJ����U�r���\zq%6�i2Q�$���N 7v��<`�Oǜ��_/U{�YX)��Ŧ�?�c�6ͅ��d]R�,^���b��>�T������b�VN����M2?�np"|�5��uTN���U�ߕ��K!9��haY�#p�+�"��"�pn�y�z�(rF���*��=��,� �0�RV��V��Z���4�����Xg�R&y�1N�awN��^�<,)�)l]s[�壭42X5��g�cE-[��;Vշ�I�j��~CP�E ��:��w�Op�4��0A�_M[@��.�����E&*��[���:�:�v��#tӃW���΁��whC��]�mkD��fIW�{ټ�ŉ9F�{�����!zh���:����[���_�����K߄ɛ���9w�����)�f� ���}F�a]��$��`�ĩ��k�nn^�X�Ed�"�/?�I�n�g�ω�u�B��fw��^�����LuK�1`Z!F�O���]�v�Z X�6�8�ϻߌ9�A1�����+��,EEqD��~�ޤT�Wo��"R��u$I�Ʃ��TiY�Y[;4���9�qGK_�d]�p�8�V�R!)��p�6(���Ɣ.��9e��_�)��8e���1Ю�q�a.���%�p�Qa��Y�r��Y�e	��5D~�P�F[2^'������ç�<�"�����'>$��j�p��S0�����+R@T�渿��sZ���b�Wn~P��͵�'�ۋ�aX2x�%�>^�I�0y��GC@�^|�|�"J�e�!�H�:6�h�1�cڿ��U'����\���5G�MШ����5��)xA�'�,f5�vB4Y�G�pL�g�P�F�ilj��ѠN��0�0Ob��Į���w���z��>�AD��8�qV��Phϱ|O��0���g���ʫ�VLJ}*z]�*Wh���2<�$T���@0J����`x�fD�H�]UX]�8}Vgިt67I�$>P;��M*�H"b��b���#�(��}K�����H��X���r��p�$r��O�B�,KF٭H�d�����^����g��@��r��T�N�.���R�D��rDSD���:�o��l�ص+�

�2d$�?)sƔ�N�N[�ܲ��&K�9�Ƞ��S�|����k�%�WY�O�k|��[?;��9r:��ﺍ%�C�DQ�Y�|:�U0�Í[`��^ ��͋u#���3\�o��AI���1�R�ۼJ	��F�e��$� j���5�Ah�Mc��Jԟ?���O�A.�bV�ZA��e=�x�lf�=�����&��j�J3:��
Rж�d������v!K�X6����O�:�i�>� !z/��{0�_l�g_�u��q!��	u�o��=�7�U�ɧ_�ȫ:h��pk	�X^MSj�� ϖ��ѝɿ��9�u;��Z'K�X���9��#l�a�M�:*�����3����������h�>qI1\�?)�Ţ�zʹD�*d=U�F���b��j��ƛA�r�Ձ>\V�t�A�3szz7w@�q�}Y5�3ه�f��<Uu��׀���D��c����¥d��S��e�Po��O�+Z�(��D�9~��P��������i0�m�X�2� %깚7l��.rJl�.u ��N9�d�A��uj�� {g&_�gF�����PxțpR!ܾ6%q�0hY��Nʝ8��Q��.���Dv�טf���L����lsJ���6i��۾�$�S�t%��j^,�]#S��Gx�'�Dtk����%��Sz ������'�!'?y ����H܊�}�8K��G��یLѮt~� A`��P��k�Iԧ�
W"*�3R�bڥ3�����E,�jPl�P�	��=��ST��a�&<�=��L/CSV�z�{�m�����&��h���
Ͷ�f^��9H��#
b3��K��j,{��P�Λ l#Ss�7���9�XX�6ôS
@�"t�6?� B��d�O�QRg���pd��	�!�WY�_|�oe6q^�|���2���/y�k$�fq˓i�o�N�/:���Ib��vQÿ�=.��-���4Z�E(�Yp/�o�(�ǋ ��g�8��~���'i�/%��i�Q�{�����31�#�-A�BgC{h"��0'�+8�$���1�4�$�/}�=�x����-ާrI��s����>v���[�("x�H��F}���Q�r �M����s1���`����0���H�����0r��w������;�$g�Rb�D���P�L#���@"�6����x�ɝPI�+o��T���� ����n*/U2��c�%%�cމ~���S�Lt�lf'��cX��q�=ԢN�J۠>MGݸopd�7-���R��C昛�ӳue-�@Z�Rg��+������/���ҷ$20E���d���[�Rt;1cը�M�A���qV��!'D����)ʛ�Pc�c�yob{�=cN/(�-�>	Q�]}�뫫R�ʈN����Ɯ*��{�
O�i1L�?<_�YR�8s� Kd3V�7'�s���� ��?d�> [UY��۝����3�|蟗GD�c��0�=PHo���`~8?�腾$�4�~4�@���=�{_-H��3���!��@M�X7{�0���*��� ��E��AD,�E����$=�AG"�8s9�Ht;u�M5�1�[�PێЦ��S2��E՚����Gv�V�}ʛ>������b�����fz���Ñ,tf�yyтs�>j����<���A0@'�Ԗ�v3K���od�8��*H�󫈂�9�@�$H���bN�8V�|?-��O��Hz�V ��#�5�B��8��nr�9ER)U�hI��[�S����S|6O��($2q}X�X-�1�&&��F��;�-��#6 �@2�����,U�!!׷�c�i�j���U���o���c$[���߽���7��� ��6�H��Lbl�����*�ً��ݜ��̉����⼛�o�`o��4��Y�0��p��!��d�(j�vS�F�J��eJ�H@�|�2��4�'���0�Ӷ�~�^��aaLlmL ���%���vr�8L*���<S李P.0���!�2��Iwoy�Q>�Umn��o�/9����1�y�%M�6A���+�4К.+��"���p2uv�����G�K�Q�:nC����Z`��v���qh�d;�z���gA���S�`s���W=ѠD�X�6����d����g�l����v�3�Qѯu���瓉�t�8�wg͋`͊M7��2 i�8�&EF���GH�����Nϣ��6ǷT}�����^(�s�E�y��=Oc���LmE=���S��HݲN?j$�u��_��a(��JɎ1�Us=�BF1���:+����zR�%C��+X��w���;q��W��,���;��@-m%�z�;�>Ʒ�����Н�.]��tD�Ýi6d�
�i�����X�3q�D�P64�W>��}5m1�7�w���<���U�3^�u�tR�6�O�z�g1Qe�S�%wc1�]m�Z{oNU*as]�ʋq}¾�]Da��}�C��q�ÿ����Q�3�¸�H�緋Pb�<�O�S9��*b�xz�;��M�)���M�]�\�"��o��#�	�2�h��ދ��[�3l�&�j�`�J������+U��$��4�;Ӆ�ˌ	�;����-[�GȜ@�t�]�ț��둊�S��dk�/����J�45��G(��8��6[��E*s���| 4�-�Z�V��Ԓ?��.Vd��f3���FMo4?6O�⡳_ŽV�z��_�1?ȸ§^WӤ���G��`8{퇈�r%�%��Mq��_�k�p�2��g'F�a1��S���5krD�t���G$)�i�2fٶ��Mh%B�a�O��L�s��O$;�~�ZΪ�I�D�۵��n�|�f�@���`��ibz�����~�{=g�Ȫ��'t{޴[����(�@&i �7��9љ	�Ə8$��+�>oœC|��"[�6��g���0�/�X�^���ot�����I���^9�S*.��hn4$�`��˱[�&]��1����n�vm��*��^�t`{1 M9`�Q��	��׍ȊN>���zpY;�W�6F'�'��\P���n��E�9W� 8{B�M��4��[��\\d���Ӭht�^���!��r���0��Ϛ:
V�R�է��C�m��f�����4ċP�Φ& �}\�~rg���x4���öȳU���̨�ж'���O����#8_��?��2����rxFxe���Ɍb)�"c�4�%)�ɼVa�ާ+'�="����EV�����/ݷ�34��q�����&�g�ť���`������q�l]0�ʠ��W)�{�a�]7qd(���C�
^
�
�|�����&���@技�M�=���K�"Hs�r������a� �Q\>��7�+U,+���f�1�����^A���R�����i9���+5���e�9S��͠<�8	�Ƚ�/�ʸL5�w�U��p�-_��0��]24ha���L����'J�۷%��R��H�8�<	n<X�Ww`��J��	�vQ;��3ڃ@j��!³M�t����T�����ƴ��R�c�^������f�6������@��m�|GL��S��r��h��tg�+��*��WF��g����g翨��c�p�c���;vAg����Q��w�I	F��iӾ�e$�f��b����,g0ΰe�I�C&��w*KG���`�/���H�������R�υ��\�@G�(j����>�{�f�w�'Ң�fiB�5��}���ߢ�6�`�.��oh��]�	�f:?1��#�_%f��2��{�j��|}5Iz�;�~��4f�+9Q~�.�N��<nȊ��;��N���bW�Iu4��%}���rLl�쪨��͐p���T��L~9�-8������Fj4\"���u&����3  ��j�K�F:�����ܯ�~[�(���y��HF')�P��aJ@S��+����\=��vZ��c7�g��s�;���j ��=��{Tc��(���
W����=��5�*�J3���E��T~>�K}�^I�׋i��o�X�������,��ܫ��S��:h�.0T�XO����M���NS*��y����Ut�!���/(�4|ʶ˲ v K�a�iE|�v�Ҙ��`���L��#9Hq�s�0��|G�������@�벉��D�����:���g�[`p�n�9bҳ�:�Od���)�YR��0 �� v�ed�J���߶c�n�3�,�&b�PyI����``O0(w�7���εd�K��{��d:t�<-z
�1�篑Q�}��bMH���s��Ī��{i�l�"鈹�!�:<	��%����P��o�6:duJ{j��A	^GM�I�W�of0{�7<I��o�5�4a}�5�V:�]�t �D�e?��69��9������A��j}�9�R^	�Վ�|�/����܂��Q���M`��<�2���/6b}6D� ��$�U��ﺶ5,ꇧ��|�t��}����F�\a���uj��4�T�v��UX�(�,�b%�z	��R����c@����}H�ڒ-M�|u�������_M�a����1࿊d��b�>RG}NCE���H!���U��h�_�㰉s�L:�<4�U�L�PX��r���-��X��;�%�I�v�hED����$��b��gm��%){kBI5���+��5�,����	�R�(�s����4�ym�[]�������PX"~%�R��>�S�c}�_[X�F�~q��"f���q�[�.��5Q�.��{�^玮Cږ�x^�I�u���j���I�,^���z��7^%/�$B���<�2Kt�K�6���pBdȀ���V9g�.w����'^�"��t��C���~v��jW�:�F��hЦ�9$���	�����ۯ�?�V^>V��bh�H�ɩ\XEc	���5!鿆��g{�?����㴺�l�WkeI��c�n[����T��&TBw�@�H� ���zV%�� b��$�<�(��L�	+�8�o����@�H�ŏ�`�;.'�5)�.?;���k��; �o�[���3اK�*�Ϳ;%��M���Mw�B�r��<�V%��VƖQ-����	�H�R��mB�� L���r�����ٿt�)7 �����	T�z���v�wңA���z� L�O�L�|���͵��C�<��#4��ǂM E��;ٯ}�nU�L'���[�{�C���@�{N�	�{/	�*���b�J�Y���ϺU���C���p!O�O�L�>]ڗ_�C���d�l	g[0����L_u��PS
�#�Bp �'�)�	�	V Ӷ��>Ҵ��it��L:cMh*�\%)�k`���SS���z%\��"�n��D{E뭸1���N��u�R�g:EҠ�ا�%��AG��R*���`�����><�%[-�oV~|�xH�La;&���y���X�˗u�
Q�\}\(�/RR����1�j�B^�vm�;Suh��jr�n��%^Q�7��	��i��~�����q�/��1�V��b�q�]���A®c��7U.L)+����7���P���DTX�s˝d|��I-�0����b��/|ux/VJ"��Z@�Fz\�Ao���䚳�ҳ�����@uV��ا��� �j��7]�2o ��G�hK�`r\a��q�V05Қ�����*{PEO�Cd�})�y��%�=h�8M7jr��Ѫ]z
m1�M����VX��ި���
_CT�|E�c�|�x�6:W���K�&�M�b�8���B)�?�z[s�IО���G��hc�e�,gm�7�c��s���� +���Hb/��������	�c5B!z�&�P�P����qf.��E��S�z�:teT+%�U�k��;Oњ}�NtA���C�lW����*AU�w �y'4#�:�U6�E%
P.G����<|��
�pq�І��i���͹���Ľ� �bl$��sڼAB�e1o�E�fJh���E��oS�W�:
��� �F�[W��F�S����Dş1(,�ȴ��f7/!�n��ɿ����xe�J�Mh�w��J��
/wuI�x���R�U��u�����ԣ�K[����c7�}�JضAO�/��5���sfi�S��v퀟Z�M��X�I�I��e�۪��]
(���� *X�r�0�.=�K�Z�t���-ݏ8kK�n��"�m&��/�����,bS�u����������͐W�*ߓõ�"��# �q��4m�o2�$�"5qd�[�^�(}����������VT��1*®�k�C�yM]��]G�E�p�4U�qD��,P�y�>�u�PJ�������ˍ�	������pL�7wÀi��d?;�yR�,(q;��	\4��
Evt�na �·N+�G�N����
7�/3s��KK�,`y y��1�^�%���7��'3^]s/A��>4auV@�����Q���9������& ��Q�b|fWsl9��Bg�ԥ���5���lx���*K�E���(:=RN?�sHl�h�%`*/oF�fǠj	�L���K������z4�Ӄ�;�K 5�m��S�N�U�M}$��\`�m�����+dƺ�'k�4�q*�9v�5��6��d�M��T��ZU�w��q�� �g�I�r7���!
K���;��c�� V56�/��t��k�]qόqq[F���>bTs��"]�~{5�)S��B-J���ǽA�@!+,�(�Q:(�w#��I�[>�?��h/�͏UH����O&����W1�3��8� !J��09&�C�(�[Q���82�<�n}���S��0P7^+8�J�Z�qO�dj�����'��x�yީ4D���:����4���>��0�����C��9j�ӑc����Z�RB6<��4W4�A,�����w��Tg,&�']>�!D�ɦa����E��ε�Sl퀝�?�P�!��rXW��6�Q/�(�d;6z�`�h^?��f<��7���<����kN>/���Ǒ�|��y˜�I���iU�Mu�Y��i�ۂ����������
�:�����uI�%�cc�[=�
��;K���H8ۖB��x6��v�I�__�|%�AɉqO�w��h7ƶgO_�F^���T=��\�X���n����b9['�%}�>p��H�Ե�s4%vU[��%̎�8蛾����k��h���&[���q!\��wB����镳��ɇ�<���*3mwj��6,������zd�P<��Ē�S�����u��H��6X�Z��3�1��)�s:��d�
��ƭ��&x�����z?yh$4r�um`�8��N�׼3��d*��,��&���H��kl�� �%��5c��(���fXd�Y�~P-�j�7v^�[�C��I� 4�۞����Y�C�H/�G���f=x�3���8�������8_�X��W�5��R��n3�
h�+M?;�R��vˣ�KBE+�8x�H��|z�Bza�q��ȗ<>$m�T_mxq�O��ˁ	\�Z��p (q���C�Q�~4�~�#�9����C��*���ݭ���b��d�wb3������Cv^��T���F��ʴ݂V�.?�ד?�>r��$�O��W}c$���$l�4:mn�R�Wv�]<�ϣ��w����G�rf�ͤ֏d�%��7�͋dkM��#z�`�\TW�а9*��z5�D�(B��f����%����z=�P9�S��Qi����V�$+�z.=]z~C����˿�W�ت����L��;�$5���q��?O7���^�ݞ�7|8��4z��JP�ˤ�����
P�;���^v�m�� �}����>��+!,Qs�^+W�����|����7��Cl����ği�-oCd���y�sF	n�KPGl=�ѱ_W�Ṻa�������!��vlH���RQ�����~��Gms ���4��׼���F�9�;��ע)l���n�$<jz!�2~m
���kf`����P^<�2�9}ֿ(�������O��_F�W��_���˜~ĨE�G[%�ԷS�T�m� ����#� U;}+���1�!�����*��*>����Dg>J@�BaY�ɬ#}�����z��9�E+;�s�rS�u>x�o��v�I�n9����^�LKD���<0���S��P���]/sor��)�ZcpU.GJO����U<"��W[����;�N�9տ����S�ߊų389�"({"p{c��@�$$a~��ХD���6[�&�I9��']e��OQ�FXچ��/�y��>�A���Ɍi���Q��Τ��̻yg%��v������\��M���	�����/�{��!�l���7�X)�<�o�b�<Y��8a2��^��Wg7��[�U�������;�X����̪hI�{�5���1q�p���=;�q�{uMʺwj��i���sπ��&�=7�졌J�*�A"H��J�_/�A;�U.J�W6�3<[�N���T�B�a����.]R�2:�D"�p'�V�U�~$����ɦ':���P&�g�̎�e��	�^9������ �-�(��}cZ`��{9Ùd~�-Jņy����]�M�������X�8͸����a��)����$�_�ټ����H-<$�S�2�1B���o��h����p��@K�
G��>�F&�x8�+���G�I8v��Z<m~�<�#
r��C!�����V�&A����2�`�+B�W�Ar۾���e2��R#}Cҩ7���(ԑ2Yݨzؠ��᭰����[T(ފK����J{S���$�P�=�ڝ@�*��:?LYV�bW�
e��?wL(*2���̗�D�C:>3-��m&�������4��`6���+,6;B
����jHǑI�<R<Րrbm�}�m���\E�9بr��TT��Z7ձ���W	Rd0@��j�����g�����!h��ѝ���Q�1ճ�̙xo��Z��5����H/��������������N�X���Fa���*�9 �`�!պ[%�)ƽ��"��"��õ�B�x��/��{О�o(g��Q�H�.h@�r�3�W��GR{��.|.=�س��=���M�C|HWR8Y�< ��-�(#]�UO74���wI�i��LZ���r:	�2*�A�8;������ՖO̊ȉ�H$���������kv�g��IQ�_o��X�G\5�p��^t��?6<����<�2�9��L�(P�P�S��>�Kr�$�A��O���o݌R��?����J���c�Ųe7����;_���`�k�?B�D!䄓S���}K��R$��	dW��WpR��{�H�ԅ�o����K�i�;|��}t�B�M�,ә�5�6�0$Y;��_�K�}�����]�����ǔ���W��*1�*`�}����Ҿ�OI��NN?��]3Y���!�K���*��K�Ev`g%*��Ͻؓ���\�d�l[B4��F'��Eq[@���|�4����Ĭ������P�H��+�|.�~,�t��� �)���'�����V�����?>��EO?wjE��� <c���6�$�OT�S!+~�XثTظB�D�L3�_2ٛ��ڤmFu�Bin˾����A����(
�D!�kB�z��5�򨠁�	��2,"+d ��rQd?�����������%/o爼L�*���n�x���\$�_mO9��p��3�qe�NQ�����K�jM�7�.k�tbm�H��o� ��s�x�ߕ���_Cl�y}���i��R�	���To�,�W�����5�&RI�jV�����R�:�yHA�`e Bv�O'>�(� �P�n�F�ݰy�6%�VB�.�b��9�����eKX��K�����%g��t����v����;oVe����^b3�
nHA	-�]�Nc.�U���)�O��k�:#�������1���h��rp�!�~�(��j��uA\�w�?Yg���֮EF��j;��X�-��T���1ޟG7d���6K���u�k�؞9�DBCM]��Y���ʿ��mm_���n��#)՛�y2����f��q+�UQ�_��9��g��9��9n�5@#=k\�n�>1��}��Vv�`6ӓ�%ZC4oz�빕���r���?��
FħT��t<](����Y��P���9�^Ԗ�Z`�H'�kT�nɳO��@$��*y�²�T& ���<~)�P:�H$��K:^b_P�l��wt�g:M��ao��R)�a��8����,�A�w��e-�[QK�� I�*I&oS>+�~�Ԇa��Q������S�Sd{6�R��r;��^A�(őq� ]yҟE�l��
38XE�s�N�O��(�~R1In�O�u�-O��EI���)4Z�ǫz��B�;0Y�ƾ,Q�'K"<fO2��d�bG:@ X~l��**��!��/�/���������ѤB���ͨL����ʷIi��0wyE����ɤ�D;	
�Ad?4H���s�	u�yĚ���8z��r�q3U�I��us��/I�ل�F�Ц��6:�@���8�2�T/-��O&W�}<��k�g���nR c�mh+_~�]��uӠ@�5M%)O�	�T�#���|���M�)���6���A^���`�Dʗc�����������zD܄��>K>�N�a�&*M��-��W
��|��cҢ�+Y�X�8Zn#K��|���P�8;j�������T%j�yӝ�m�i���]�<$�LLɹ����n�ťlqM=��=�3�h���]�b�0��Vd�D��"�}N��nt�[�u���E��M�̼Hʹ��|n�5o]�/�������l�%��ڊ)��0^qu��~�x�/;��;�����
~(ӓU�6�p۵���d�+��r��KLa�$��d���AAz�Ļ�	M�R�pT�Cİ���J�]"EBL`o�T�t3!nh�o-XN��A�O��L�c@�5),��N�6U���S�}m�ɇ�Y��>Ʋ��̔�_�X�����B��]MR��F�w����Bq7�Ğ:��Q�7���@/�3�K��d���;���
<SMs�r�P�Y�Z����"2�� �EbۥD(���GKdk��X��h��	�KC���[�0� ��Q�5���*�[��p�S�ʋVyu��r�e�?o.����C���/d���������Q��l�{����{���,cY��OM�`��e�a(�֎����Mj�3[R%qAǤc8�cs�M��m��/Jm�#�Q8�-�]^�-����3�"��>�:�Ċ#o�>�7ʛ���zP_"�eB�E��J��2�Z�I��s��9�H�n�Ȏ�������z�@T�6?n��(\F/TS�k��%�W���aE3�s����(�-,�������EWx,}g��#��/"`��B~����Q��mZ� �����qmz�"1��8]v�(������I���y��	@��/�w�tkS�)Eu��Ξf4���*��9=�%[$���O�������1��@��#�\���l_��.�,��.LKs%��s�̦%�#רFk%��8�笗��!G�t�8��*�س09���xWǗ�1��$m�q�9`s�����^�2�0u��	:���~5�U1��MX.*�o<鲿E��G;?���nh�k��i�bL�b���o
H���9�}"Tŝ�g�	r\epw
�1��Ma�Բ�ќ�ӣ���C��
�IQ�W<�T%���S��:�*�vh5V�S/1�R���N~��PA�m�J��ߖtv�tP���=;E߆���MK��*�,V�����<m������V�����? ��8W!�,1�?ý[�����a�W9��i�NE"��i���6��H�wl�)�_�?3���~n�?3c��6�d�
9/2��auIH�^��xⓍ������4ӾlI���7�3g���Q���jja�"�#q��T�b���v�>a����Tt)5M�w4ٙ}�jlm>�+�Ӏ5���8�Z���RP?!��Z6���@�\�<,���N�y!������f	�C���j�D~�ޘPpnӯOsX��U������I���*����@�dhs/*.�r����Pa���e�Ga�Ӿ�M `hD�/n}��M��8s�o�Z��M��M��W�R-N\�����f�9�>d�'������+oK�k�Zht=�����>������A�wC�I�/��UU7++��d��������%���� u��P�����@d���?�HZ�s�{��l^}���~D?H�Z�T8f+�$��zF�3O�T9m�H4��Y��Q�t�m�����L���ㆆ�H㰲�H��C<ѩ?=SP�L��� @��
2��N��9�[�Q^nc���)��~�������(���Qr-j���r�����>v�?�>#(���ԍ8����lP�+|TR��&vY�q��_�-�nٻ�u���w��c���X���\J�������l��١���N#hmQ�9�B f��.1Ej.�إ�
��R��Q�H����@[�4��3J{�~ۥ�8���b^��*�9/���Ąh�i��N<:e����Sbx�7�b�+Y՝00���d9�8#	_��^���S��z���.�'NA:��I��B�b�<&���F��a6��~��w�����@�t	��N�Ic��P�y�o/��?r���G9�=~	)�6���9�4����z�N�%B��'<���ɦP�&E�$��4p��p�VO�NUf�U$�N�ʴ����-*���9=z�W&Z
��̇G⣼���v�	�a�g}�Zn��r�~��+��m�$8�=���|�� ��i�r���" ��|�vc&��gJ�B�o�8XYķF���i��qR�����"�w�@��=����"�<��J���+���L4s��w���f�@�{^'���c�h�@.K.��)sy���C�[����*X���NL�s�Hf�kl����i(��9��h�.��R�IF��Cz�
-��0���2�EBդY��q�U=˒���]C�H��\��(
-)���n���K�8���u��C��ny�n�Ć��wą0�|4q!�$�E6]���454|��00�=[��D���J��4��U= �"��O�e�3�k��}��:M�LI�� �i�����x��y�7���C�4N�cjXYOI`�m1�S:�8���*�c���Dl�������<�F����P6]����q�Y�T��U
��u�W:sl�5�p��V���ő󬎠�.��\M�����-�@<f�k!���Gˊ���>�ŸQ[�ǫ]��ҹ�V��u��@��?�#R�t`�S[Qi�@K�m$T �!�n%���o�k�$ߒ�!BKTl]pȉь�i	.���6�'�x�F�D;u�W�b��,��Ϥyb@w�EK	�f���Gotx�HTe�)���.T�;Htj*�oa���7:k���@�|Hs�zW���2��1$�h�����ȥ5��0�2Ւ8�2\���,t�_��,㍌��0*�.8}���Q�ͺ����%-�G^>)���JW";a��^�)-=10b��[X*ο����L
F/�C���؝+�[$�g��U�'���'(fm߯��$GŤ��oO� �lxmy[������qn�t�UT.J�~�@����C0^0gvb��;�����q���7[��}|�h�}z��!�m(��A��H�F\�A��vY�d~����uy��1���ۥ
���e�Y>R��㖽o^�76�0�N��e��YP����W����b�KD�����&�[����������ᜫ�O��^D�X^���xn&�Y�-�5ޠ� ���?�,���Qj��^h����#���1(�W��C�5;������.\n�'�E��:�-i2VF��݁�w/��N6�וm��I�W�)w��2`�o���[n}��߯#l����P[��w��?��"IC:�9�o3�����_�7%��� �(������X"΃9�:��|EF�0�G�M<_�, ��mH皤��?�ޗ�\)��{�vW_���-�fߊ	Z]���Sp��Q��>����s�(�t�6���p츏a�i�3T�YjAg�l������U8`�I���z����ޮ~c��#�3o�;��1��_	�����,um"y�f+U�;����Q�N��&{g�쟡�/>e�M	AH�9KEZo����.b�u��l|[7�o�?�`�.����@��(�
>����t��X�o��%jWuW������U%��2x=UFp��}�/����cX�4������Q��	b�Fw�[��r$��G(�{t���4D� �M#0�l��)'SM"�q�mVuAol�T�qEJ�B:�o�ޭF{b�!%|47Cs�Mȅ7A�IZ�ކ�/�܌�����$�)�_��2pu�a��`�S�b��K#ГF�A����,�|��?b��\_������ō����ԥ�i�¿��=�c�;jr��������kse�u���}���Z�c��+nH�c��˘���0B�/[��u��Kt�`�E<o�$7�(D�u�.���|Z}����)+{0�&��GF*�z����n�R27A��1�kAqm�^��ٿ����$+)_h[#�)s�G�bl�0�p�U]��|��.\Ihb�`���U��,�4=���E�<_�\1�a<�ذ�������Y��"���F��1�q��SJj�r�Ɨh=���ߩe�K.I��r��a ���w�M�yQUe�#.#`�I���E����(%q��F/>��Ʒh�o#�?F�{�D�}�YAQp9�!�c��3�,07�k�^
��1��v>d-aLť���&�c�~��K��έc�F5/OZ�`�z���h�V���P�/@b�K���5q���I���,v� h�ÛI>�\pV���9�i�e��1��K8�P�|����x�M���/v���\�����k����F���z��U�!�8K)�Ox'�s�8u�G��}o�D���?Ddp�.������j��K����6���wh>9�Yh�yb��wAg�="�Nh�Ϋ�S�$��j;g�[EC����/���,����;�<j�U{��Y��
b���5�p�YA�AP,��$����B��2���L��s��4��!/Q{��?���j1nE�Wnyf��5����mV0����L�%�z��Ė'�|�i���5��&j{�	�� q���r�=m�ڥIWe��j����u��R�w^2�$�i��������q�#�FǫF��o���|y]�i��C�����Q���hV@b��	~`�~�W�>��t[9g|��Nq�u���D�Y�܈ ُ���T�"����x�Ir,�'x�b���\���a�|P�ck�, �{I��`�;�:�G��`&�l��L�޲1U�J����m���8m��#Y��X
�ݙ�
=(Ֆ�Ʋ��q@�}% )�X����0⽁XɓGc4:�ӭ.�$�:�K3�^V����y6��*�qM��-]&X����X��\��w�cDD�ϑ�3i3}��m��b���-�N�,�& zGKA���l��ϸg��ehz{y',�L�Ae�1N�*:*_�MF�v�$tj��c ~j�f즁�����%��=+)��V�>w�~&�;�X�%�G=2�Zrf�T�0�zF��;�V0�� Q���UC�LA��:;��)��(Ʒ�8�0m��z|�d�����S�;gsx�j6!2c�����\ꮼ��e�:���*Cw1�\�}6�QY�D�`Z��u�� ��,HE�����r�?#��R���h���E;�,�uҤ�=�H�F��Wtͤ�Ѩ1� 2�z)�<Dz�����4��͢o�Ӫ1���#U��f?w���zGQ�8v��������O)���޶�������Q��;�@�XP~�O�?�4H��Zf� �AD�U�IoyJ�R2�֢��_8�� �!���:�1h�_R7۹~��& ���������NK����+�7�����i��ם��V��~�V�DѯŇ�@�>�l��}��=�����w0;�(g�%����f��,X.$�^X��N&� i�ӳ���]������P�h]����o�'�z����6��5����R���C5h����_�0�!4��$/2�h�(I�Pl�Ej%#��ɽb��C;Θˡ+=��e���/d��fh���q��E�G5��
~��^z���=4�NwY�o��h�۩�S�L��4Q�g3�"�t����6)沐4�Y�`f�;�-q{UX�WCI.M�n2;�8�΃g�7rmD@MֱG^K����U�o�ï��[��b$5[y��ˁ�Sj�IH8�\x�RJ��fxxM��t�J�i�#kq�V�.cN�Z)��J�9��֏�W����KŻ
巁�Bf/��vQ�1���5L-�p�7_P.�~_������\#��z�B��.��b9�Dt���R��4����Z|%���B:�ԋ7k�P=������$�+E9�Vo��j�����Wh 2*��R+m�8���L��a%%$}$�W�����)�����,o�����!��FSb���6�d�M�&(˭;t��wa2,� ��M_8����	Dp��0���7A�m��Ok��7fP[�BUx\fe~Y�����Q7�Y��ݹ��ө�SD�g��ѥ�F�-U�e�9ޠI`H�Zp=µ6�#��g���{TK>s�l��֖�!�t��;�v������w�N4�؝kpX����꟮y�׈�����j����7�g�Aʡ(��l�!! ��E ��NUk
���j����M�P�]��3 �~W��U���O3"%�`@�v]�d�������'�^�G��[��u��T���s�B��xˍ67���������
��иy��{��8!=�����ޘ�*���2��7�犯=�P��5��[�����\���['G����ϥ�����smٝ4��Vx���/��sP$Xޫ1��+I �"�t�������5"�"+)z ��23�Q����4�>�W��[(�(�BPִ��{��N�H|�.�6��T�pN�2g�2M�!G�M�ӓ]5Jn������luc� :��¹rf3���[��N�6<3���7��~���߈��2�c6�M�l��ei�gB��5��2�2��3���[*iD����(B��w��T�^a����k���+�H���6g�B�C �h��=|G�򼕊_���T��Y ��(����X�l���l��T��7ꮁ���u9��T\��:�Y�BO�[ό!�����׭��3T����34��@Э�NM0vܑV���t�t��I}&n��'����I��1G�݀1�{z1Tz�����w���5�F5��``��Q�Lggi+���Ou�_W�P�:x��
d]-�!���0��O�oET&UO�P�پ�,n��>����e�C��70&e��%���J��8�g%n掃w��O�����kH�$�	���L���[9<c���*T j*C������Wn|�c虦�#�#��g���c� Z"��kB���5��������	�dI�#Z�jϴ~�q⦜���0����3B�d�oQ�-y��%��#�z��C.�0%G�$��;��c�IS�<�4�rD��W	)��Ѓ�&� sƾL[�i��!$�"�ل�T˃��r�7gV�[�h3k���ɻ��q�C�O5!�*��w+L���N��xk6dU�-0/^�����搌I s�W&��|W����rJw6�
+�9��o� �g�pK����k�'��JW�Ԑ���r�w��}͓ �6g��X��-!�����CWv�W�����P��^Ď��C{$Z��K���o���L����H���b7ڴ�M8@N�uJט�(�$�X�MJv\��
`��J�D/���fe��"�{G��7C�v��&I��ڡm`��>*C�x�FF�|�ȔRF�<��Օ�'�����Z�A�}��z�J�u�+m���^/�u�y�B
��(p�V3��D�Y~����������ɍZ�Z��H��v4P�rnP�� ��8L�3[dg���
�.a�x��	���R��
���XFI���3v�Yk9aG�˩f�����=r�,nDK3����+bb��bh/1��9Y�i@�!PT���#�2�h�:.�	�5H Z�O��$�S�}v�r���u��ӧ�#p.!�q�`r<m
Q�nn�'ɼ~��T��CZ=t��)X�d�Dc'��C�,?�L��vH��}<�9Y'�I�YUt�bS�j�:a�[���h2�(> ���F?����@�E���a2}[����ܘU�-��[�f��%��M'����%+ȳ�U@es	;<f��� L���&���J�G�H`3>G�oq��\� �W&:\L�2|����s����+��k�gE\
 `فJ�#3�bqe�����0�D >cf�S�n��%������@�%^y�6�����=�� ������VF�7�js4��e$d�b
���6��-��8\r�!g0m���i��f���˶�e�4y�g�-����e��j�R���9�'��S��Gu��Q�.�E��|�焰����i��)��j��-������l%6�h�k�V�1��J��\�wίm�D�/��F���&G�����×�#�L>�Q��m���śoX����an�ά�~�����`WWǼ��}��hN�������Z��s��Ke�ʊ�b�B�o�Τ�:�::%)�)��q�;�l�5�}���A#� ��O�9}�Q*cLai��L@_�Kab92�֬g%q6WJb[H�Ϭ��8z�E���߁�ɡy�}�W�H�8|�/W��oD�i�B�~��'4�Hّ+t��bs�Py|`	N�0m�kX��^g��sR=׊�h���x0a*�d��9�����d���.W_y#�M#~a��)��X��6����ɹ����P㔍� L>�t�v
 0Z����_�5zgx������ HG�_k2��D�Q�h�T�il�Pk)�p���`��o/�Լj�V�D�#�:qI(�$�WSXB[u݀�����T�Z����D�iB"�f�ɵ��X���=����q�p2w��s����y�pEO�,e�L����v���L%�ܭJv�{Za�9��75���6��Sbx����mI�Ѫ`X�J��8�B��O�"Z����B�&�a�<sЃ�c 	m�����o�}Įv��� �>	�~>���#��v�WT�gW���íR�CB�L�8�>��m�=�,r�<�:�WC���M�]�#+�,��^(���a�,�U¥i�u��A���AQ<7���J��Q�k�Fֵ#֚V����v �V�&Y�6�b*�n��%��`�P����c�e}�.��IS��ƾP__|���L��q�<���b��P�~��(�]��dW&3�M|�\���vG[I�Ѣat��%�T��M�j��0y���c��"V׈�e])�>$`��0c>U=t��ת�Lj�B���at ��n�����),ilP`H;	�;�zphpv�a)C<|��F)�r�(^�q�#d�, :�u3N�����������\�i�}�h�K,)��j�[��꾹�0�첈\�cs���9�=�g�.\I��S�}�e,vC��l��ݲ�!���	���Ϻ�>#�WX�
zm���a��&�pc $,^1H���2i���_� o�dd��7Ğf��w�ӏ��v����r�5�D�b�r�cL��:��T˥c�*-0�?[x��x�>V��끙iS¥Mk���kߎ����)�blJ3��TG���*��ʄ^�!U$C���3a��"|��N���,6N��%�rϜY�T����b�������RF�t�D`�wsp |��f*U��͎�����7����7W��>�	F���R��E��~�X��/w�c��u:�w�����I���Y��Y�t�Z��q�S�<G�sN��S�<23�s�`�H�ȧ0�2��
Ym�t��"�#��B�m��Yf��]�a�ԋ]��-��\)!�� {�~�n��l8j�{n�?+�`V^gc��}Ҧ�9��	*��"�s�%��2��3��zZ��@�淄mg�x+�dXtQ0v �<o2�TQ�Hab��F���p����n�RA�ڕ�l&\g��%��Ȱ���+�$�� �+��ړ]��mu
/E������^��] �)N8��)�+�qf���ALَVjی6bG�V;n��}�1ZK]���l�3�2؛�їJj�ݤ-�S�*�#���ǝ�3�D��,��)Q[Kb J�W�[�V����_��Zw�>���U6 F�����޵ԩ��k��:�Pq��W��L�]�D�nJS�K��y��!��㙘�,8�UD�9��5�O��Ae7�(,�}��5<8+�����٥�1Y��/ Q!Z:�_O��+��\�Nn%m�~8���ᒅ�Į݄�o�q$1C/�.ݓ��'{C��՜(��-!����;��އ�wI������A]R>B�7{�!3w����G�+�
�*�@@�U��d:x�tUL>R�i"D�b�D�'I�0���z^.�HJ�l��5�X��QP��ԙ	�X�#d��H�e���,7����DZ�)ph��}�MS��3K�����hi�Ay���h(�wc|O>�����	|
��i~w?(I�4�b]e�W�V ����؀@���wtA9�Qq� ���1���C�_�4T����_Pj��V"���'��q�F�ܓU�O��K�TJ��Py`C{LX�+�z_����hN踇
��x��s2���<ř����bF&!��$������b&P��\g%��BS#�����̼�e�J'ň.��btQ��j���#	ۮ�$3�'«$+$���F1��EmQj�q�w�h�QD���		3g��Ӄ���$xGa1Xh�IW�#�jH*��$3�G�)�C�)��Pݥ*DӤ�*�:�:�t�i�8ق��*
��
�a��!�IySRQ&���]�h}����e�غ��*�N�g\ܟu�f�z(|RD�\PИ{M���4�L����<����e@dl|�H�n�]�-'�l��{]�?��R,� m@�rϕ�闪�'X�t����{��=ģ=��	W��y%�j�M^�WQfG��d�:�h�.�E����_�Y˓�����!Ɓ!g�S�GReve�XC�O�"O�ִ�aSv)�w�ܧo��ϵVR	f5��OgIch��/�_;mb�,�:v,�#9w�]��/$�|K>=̍�eC�ds���;�M-9N��E;~��+#4`c*"��
`�;U�{V��;,Fs,J*y��r�ȡ�D��-��C5*�s������y7aXpk#m��1��j���œ�.8
/�:."b��q�ُct�V&
��jY�=�
/�C	��Q�?�DM�&��U���8�/�����<�����HƸ�y~,j(��'k���iɑ+��.c$��q���H�� ��gs�K'��;�r#�mБ`�P�7�U�'�س��	��'j��%ƫ��f<�Gd��go�4���)s;vdii%'���ʍʿR:��g�@#�
���!n>�p�h���`�ڐ՟�j�R��܌�R��ٱ=���(zn>%�Lw�p�3~�4�/�Ez嶖}0dYF|�҂�"/�*���ur��ƾ�6�3�\��c�:���2���5�}����i�J#lxG�;��ت�8�fo��C١鈕Y{���@ >��@<�ĈA^"H�I��L|!*��s�Z�9�z���LDl�j�G�ӕ�B�#Ú�����$4�|���13X}&�F��j�jw��g4�} �tZ�����$-7	����7V�,�~�G7�4 wɓ��.�2�'O�ҩd�V(*D��*?�	VE�N��]R��p��:M��Ώf -ƚ��4�D�qC�0+��=Q��ʕAjN���@j�	@����Y��t�dg���#�;_�H�F���I
yZ��HFN��.����$�Il�q���bISm�3恗�d�KJ����sήN|��y���+̗ǒ��/b+_����u��^p���p��V�1eS�ܸq�dk6�$!�҅O9u�#�un����]��1��'���޾E
�O��޴��?�Q��.�5��qsJ�������?��~����Y��i7�aͷ��<i���E��v��=��|Ŭt�U�,��̔��k���Y`��M ��#��:�v�,�#�M�]I�6T�3m�b�RV���²{N~�-���v�^]���b�'Z��ƴP�o9�Y9��b|�X�㠬&FS4�G�>9����9c��#��EYJ�N�L *�k��jqɳ2�m��� �`^'�1���d.�J*<W����'���Mr| �ѱ �bLt��-�G�&� M�mJ/��/!��2�4[F+!� #g��rW^�!�Li9G"��[y�9ˁå�	�fN#ԉ��P���(0S��g��}�<�5�/˸�8���r��"6qW����q���9�K����"�V� td����l���W��[��ml���®팲���T��΍��-�G�e;Jf�|�B�c`����sT�Y�����)�3���8m��Pj-�E)�q�]%�u��o�x [*?�2P^��D]oF�9^jno��'��]㣿)����\Ԝpw�$���Zw@�j��P�6�r��|u�3P�=r��m��(���N���qNIF�ɗ"5�`���|\t[�e(xZ�:'l�f��SFt�u���L��?(I)t��
����n���uT��a���!���+��L��_�u?��$��Q��!m[��\z����)z��D��u�Ck��J��ZT۳��o������(.Qz��C���ȿ���������TFm%�~|�H�R,�D
䜛Y�v��Ms,��»��M6�ȿ&hN�0�>%�X��X�����U��@���gH�X�v%�������\�C���6R��:BM>��p�y˙��sfApYB����#� x�;`X葉i�� ��"G
b�D�^q1�W��`�z&/.�l�'й�T�1{�e��U�^��4���U|���푡g����:�G��ɔ�,�����?��#C��[T.�K?[���m�-��`Ǝ��LC$!p+Q'e�x��{j���O�r�>��%Z�л�Ͽ�'{���56�4����{�K�z��l� d_�i2\	������E�$C������xV�L����+��pd��V��^��W�g=�'���1��\��8�-�����Q;�1�hT. Cqƞ�NC�P�"*K}@�z^ɑ��B��L3��w�����X>��C.��4�N���-�����>�<�h��|�?M��F�U�=}f-[{�9@�_�v�����ÎIf�]�;�UE�1�-��T����� ���Ak���ń�cǌ�W�%��o
����P�����P����4K�*�DI�n���@���#D��=p��O,t��Bh�7˄�mc1�Cڅv����,H��*��&���2WV]����}�"Z�O�`���o����&�z�k�ڠ��ji{G)t�B|<��fѓ�X�t,v�T5��2���U���k��ց��F�I����s�R��=͂Dۭ�|�@�t��[_��8��<���R���
	̋>�ៃ���
V�i��.�z:��KeB -1A��]S� ׬*k�̝xˋ5��G�7.,�����!��&�31�F��9����"���	>�)�N�%������iC�,Y�oz�  �l�RCǝDs'�ҕ�Ƌ�F�Uk	��N6���펖uE�y8);Cؒ(�j�r���GFo*�|<�^1Ub�9�%��WZ�$��R�O�TB)�s�r�ܑo�9�H�3�(���h�9#\��~h�X���6��8�
�J"hK�Ca
���P��������[�)*;��;�������+�}�DB���j�D�$��]� /2k��$Je�����$�W4�#�R�~u��{i
���,�˙�!�E��L�`����[gN�w�)�&{BF�$(�)8"�nOr6�`�x�Q4,Ʃhkr�ʒVШ�~e�$HƲ��m����vB ���x��q*n�*��Wg#��L D��c}O��z4�ȕF�<�e���`�1�vƤD)�kߣް���@j��ܚd'���@c��`4���]	��ǃ:�eDA�%�)���k�p��v�Α���� ���:��^n@��G��5�+��܇�s��?�p:��IsH);߈Jv���8�ާ����_�e*/dg���8�d�Z8'k�0¡�����K����G�2��ƷE`3ǘI���p�%�Ίe�0��DQt-�?�ϼ�j˥sZV��n�Q��da#"��|�Ӌ"�/�w��r�hJ���2:�q\�#��|R5�B�;�E���L������0�����ф����PY�ۦ^S�F���p�-<Zr�w�fH)V�y���M�L��b5b��6���Y1�NC�����'2Е6^h-C����N��!�"��FBD~[~�@�s��s�X�@�8�C��+ѻ���(Q�']�Ŀ�n4��(Nh�<I�M����Y�T�xR�n���s���&��.`���>0᏷����RėT	L�AΓ���;�!�Y`9��<Sf@bkR�] y��`A�)�c�S�Y�|�����J*�#w�x�vc�"l=#���@�"�TkA,,�������k2�k%2bY��~l�{�^r���
�����[�^�������lo6t��(�w��e�o+Ĩ2�^��������ֱ��|B>��O�]�5^��-^��&�'�耗d����8��5$��zP��`T��l��KY��7F�PWf��#��ԅ#8�T���`�ޚ_��_渷��$�(�'m�?Ze2�6c'�I��s�C�����քM�0т��Ƃ9�j}�6խ��.��˨��:F䅿��1	u���i��½�?� �DX�/������-J�P��^q �l=�0 �(7�W�����zV����Ί`,�U����$�`�n�S���	R�zc,�[�}&YQ��\��s��z����M!ų&Ǎ"}R�U�]�D���v��f��4S����I�����c��ݑ��p=�n��r����bLfҌ^d��?�f�YVs[^�eN|�UR��ȗ��Pc�}o��1NX~�c`�Z~U�ww;�#6�6"t�5.������� n,Y�6������'���<<��|�y�°ɭ,v�8̘���Ђ�(� �\��]V�'4���c0l#�H��B)�L�N�u;��ڔ�VuO��������m���#R��/�x��srk��y��*��v�������xe�#W_����>.��;�\��lf�*%4
t��X*"K|-�y��
^����@��و<:�������s#%_!	>9e�lN����~�����.Pb��`v��<r�(�#bGw48�X��yR���<l�޼$��7���yy�j�n�ੲ��O7�
�p�����{�߄���	P���4@��1~�E(=+�
y������}�o��F��	|��D��j��U~�IC`H����I<�ˤv��d�5�=�V���������ӊiYyE�j�=�gQ~��AP>f&�M)D~�6s-t���[�g�tn��@z�-.�O�پ�tt��]��4
���K����r�����l�'8�E�a���0w�KZ��n	�ꐌ��\�����/Y���w^�T'o��C�*�YϵէM5]Q�# F�)����"`�2S. �H�c�GQ�Ku�ʮ����pH��L��R�	G�!��Ǝ�\�*Y? �'��N_PM=��5M�2k�9�ﴌh����*�����n(
\�n�Æ>~�;�}�Y`߅t�y�8�e�P�����k�!�T�f��]2	\�W���b%��y�]�)P$�L�)�*ѾA���"����u ��M���J�NҎ-���}��n�`�?���k-��L"gbi���_�\k6�+�E�:*�{� t�	kZ�\�c=Pܿh�ёCo\��ȰEүJ�z�=��g���WՃ�jnh`��`�\g��O�Ţ��a5�S��a�Я?+�=wks���=��e=��H^��H���K� �f�!<͸�|'1J=�ڀ��V,zt	��jr/d�nP�t�)^��-����G2�c��l�hs��@���̲ڋ5�z��k��>�8܊y�/�l&eq����y�^|�w=e?3��F�k#���J����W�b�ȉ]]x��v�#~V�huW������z��MLY9ӗ�-rp��y����h��#,Q��P�aɆm���9��$x���&.�L��|$55N�L�� [�M�P$�X�g�c`�kQ��������YtW10�mK��|�oa�F��?Xc�f�����]Sױ�c�\I;����qa�M3�����`˗��Fͩ݀sR��ٓi�ir�`�UoU��h%L�$6�ɘ�i��	}c��:9���7�mˆ3�;�,��В�{��Td���+��rE�9M;���«����.T��
U� ���i����&�����w�yÿ��tؤd�9uc	gو8q.)Hߑ�Q
>�p����y�6�r�,�'bٛ\Lte	g�& ����.��~]*a*��3��40�����c��r�&#���6>�\�}�Pْ�+2���?9����RJ���u���+�ijKk�ѱ�b�fP��GՈ���h��v��13$���x���ޢ�)����G�&�F5o������*p�ں�tyf���$��y�D��QW.�U�yK%�\��=���?Xͫi9�za�K��b�3�|�=����=/�\�q��x:{%C��������*��.����r/榚�Z��/�sFU0eڮ���׼ �� ���H���t��"t<�}���%���&/:�k�R'F!/V��#��A�n��5�[�&1�e%.z�3�d��;�$1<k�7�b��g��� �v*���j}M�.e�^�%�Q���Y�`zHz	��B�M����l!2�ʷ��ɀA&ׯJ�>�����7u��?�(�n�ݑ�V��|�ݕ��#��˅�Y�T���HU�Z�T���/4����Gϛ�¬�(�4�S��\����!��/���tظ4{���%��g��G����1�,f�gB)��l����C�?J'��P�X9��Y�Ւ�������k��s$�L ���v8���Z�m��� ��%9��@M؏|��h7r|غm�tK'��6{ɉ�����(�x�l��y�/�]P�F͔MJ��re�R%(vs�L��I�="�(��,�E41�3:,��@���|XH0��v�����!�*ڸ
,�l��.+�s��H��q[ f��o���U�1��L^_�M�B��3�3Pg/T���M���O��W,��]ӧ��MM$Z�9�����&^��h/��C�UR��E��z�^B�_~�a'h2m�7'̙Ɍ���V噉G����*.��'
ͤ"��}��D�R7��p�a�j��=�/y�y*�Ui�)Wt���G��i��6�!���eUDb�@�^<2�'�&�"�r eG�C�b�u�����0���r#��,��D�Ez�B�Sˑ��k
�^�}�[�4U�+�SN�Ϙ9��S�,�-�Z����|�ᤪs��X'��kߤPr���x��bP���
�O0�_n��#4��o�Ϣ��d��q���0��:
�&�&@�L������8���\��t:���|͓�o�
WJq�4�Y=0X��(��Z�V4m��|��/~&b.�q�x�b]X���O����l&�˯{��j�`Q��Aɡ�Q�=W��� ��"�z��H���Rn���_TO���"�W�"�j���u~ey�ɪ�&e#�#h